* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VSS IB VINN VDD VINP OUT
X0 VSS.t49 a_8360_n43060.t15 OUT.t37 VSS.t48 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X1 a_16582_n43566.t1 a_n1924_n43526.t4 a_8360_n43060.t2 VSS.t6 nfet_06v0 ad=0.78p pd=3.52u as=2.19p ps=7.46u w=3u l=0.6u
X2 w_1750_n43456.t42 VINP.t0 a_8360_n43060.t4 w_1750_n43456.t41 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X3 w_1750_n43456.t45 VINN.t0 a_2044_n43060.t21 w_1750_n43456.t44 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X4 VSS.t47 a_8360_n43060.t16 OUT.t36 VSS.t46 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X5 a_8360_n43060.t5 VINP.t1 w_1750_n43456.t40 w_1750_n43456.t39 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X6 OUT.t6 IB.t4 VDD.t55 VDD.t54 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X7 a_2044_n43060.t1 a_2044_n43060.t0 VSS.t8 VSS.t7 nfet_06v0 ad=2.19p pd=7.46u as=2.19p ps=7.46u w=3u l=0.6u
X8 a_8360_n43060.t3 a_n1924_n43526.t5 a_16582_n43566.t0 VSS.t9 nfet_06v0 ad=2.19p pd=7.46u as=0.78p ps=3.52u w=3u l=0.6u
X9 VDD.t53 IB.t2 IB.t3 VDD.t52 pfet_06v0 ad=0.728p pd=3.32u as=2.156p ps=7.14u w=2.8u l=0.56u
X10 OUT.t40 a_16582_n43566.t2 cap_mim_2f0_m4m5_noshield c_width=50u c_length=10u
X11 w_1750_n43456.t47 VINN.t1 a_2044_n43060.t20 w_1750_n43456.t46 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X12 OUT.t35 a_8360_n43060.t17 VSS.t45 VSS.t44 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X13 VSS.t43 a_8360_n43060.t18 OUT.t34 VSS.t42 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X14 OUT.t33 a_8360_n43060.t19 VSS.t41 VSS.t40 nfet_06v0 ad=0.78p pd=3.52u as=2.19p ps=7.46u w=3u l=0.6u
X15 a_8360_n43060.t6 VINP.t2 w_1750_n43456.t38 w_1750_n43456.t37 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X16 VSS.t39 a_8360_n43060.t20 OUT.t32 VSS.t38 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X17 OUT.t31 a_8360_n43060.t21 VSS.t37 VSS.t36 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X18 a_8360_n43060.t7 VINP.t3 w_1750_n43456.t36 w_1750_n43456.t35 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X19 OUT.t30 a_8360_n43060.t22 VSS.t35 VSS.t34 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X20 a_2044_n43060.t19 VINN.t2 w_1750_n43456.t49 w_1750_n43456.t48 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X21 OUT.t8 IB.t5 VDD.t51 VDD.t50 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X22 VSS.t33 a_8360_n43060.t23 OUT.t29 VSS.t32 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X23 OUT.t28 a_8360_n43060.t24 VSS.t31 VSS.t30 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X24 VSS.t29 a_8360_n43060.t25 OUT.t27 VSS.t28 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X25 VDD.t45 IB.t6 w_1750_n43456.t0 VDD.t44 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X26 a_2044_n43060.t18 VINN.t3 w_1750_n43456.t51 w_1750_n43456.t50 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X27 VDD.t49 IB.t7 OUT.t38 VDD.t48 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X28 w_1750_n43456.t34 VINP.t4 a_8360_n43060.t8 w_1750_n43456.t33 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X29 w_1750_n43456.t53 VINN.t4 a_2044_n43060.t17 w_1750_n43456.t52 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X30 VDD.t47 IB.t8 OUT.t9 VDD.t46 pfet_06v0 ad=0.728p pd=3.32u as=2.156p ps=7.14u w=2.8u l=0.56u
X31 VSS.t27 a_8360_n43060.t26 OUT.t26 VSS.t26 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X32 w_1750_n43456.t55 VINN.t5 a_2044_n43060.t16 w_1750_n43456.t54 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X33 OUT.t14 IB.t9 VDD.t43 VDD.t42 pfet_06v0 ad=2.156p pd=7.14u as=0.728p ps=3.32u w=2.8u l=0.56u
X34 a_n1924_n46660 a_n1924_n43526.t2 a_n1924_n43526.t3 VSS.t4 nfet_06v0 ad=2.19p pd=7.46u as=2.19p ps=7.46u w=3u l=0.6u
X35 OUT.t25 a_8360_n43060.t27 VSS.t25 VSS.t24 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X36 VSS.t23 a_8360_n43060.t28 OUT.t24 VSS.t22 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X37 VSS.t5 a_n1924_n46660 a_n1924_n46660 VSS.t4 nfet_06v0 ad=2.19p pd=7.46u as=2.19p ps=7.46u w=3u l=0.6u
X38 a_8360_n43060.t9 VINP.t5 w_1750_n43456.t32 w_1750_n43456.t31 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X39 a_2044_n43060.t15 VINN.t6 w_1750_n43456.t57 w_1750_n43456.t56 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X40 OUT.t10 IB.t10 VDD.t41 VDD.t40 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X41 OUT.t23 a_8360_n43060.t29 VSS.t21 VSS.t20 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X42 a_8360_n43060.t10 VINP.t6 w_1750_n43456.t30 w_1750_n43456.t29 pfet_06v0 ad=2.156p pd=7.14u as=0.728p ps=3.32u w=2.8u l=0.56u
X43 w_1750_n43456.t1 IB.t11 VDD.t39 VDD.t38 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X44 VDD.t37 IB.t12 OUT.t17 VDD.t36 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X45 w_1750_n43456.t28 VINP.t7 a_8360_n43060.t11 w_1750_n43456.t27 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X46 OUT.t22 a_8360_n43060.t30 VSS.t19 VSS.t18 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X47 VSS.t17 a_8360_n43060.t31 OUT.t21 VSS.t16 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X48 VSS.t2 a_2044_n43060.t22 a_8360_n43060.t1 VSS.t1 nfet_06v0 ad=2.19p pd=7.46u as=2.19p ps=7.46u w=3u l=0.6u
X49 a_n1924_n43526.t1 IB.t13 VDD.t31 VDD.t30 pfet_06v0 ad=2.156p pd=7.14u as=0.728p ps=3.32u w=2.8u l=0.56u
X50 w_1750_n43456.t26 VINP.t8 a_8360_n43060.t5 w_1750_n43456.t25 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X51 VDD.t35 IB.t14 OUT.t1 VDD.t34 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X52 VDD.t33 IB.t15 OUT.t7 VDD.t32 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X53 a_8360_n43060.t12 VINP.t9 w_1750_n43456.t24 w_1750_n43456.t23 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X54 a_2044_n43060.t14 VINN.t7 w_1750_n43456.t59 w_1750_n43456.t58 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X55 IB.t1 IB.t0 VDD.t29 VDD.t28 pfet_06v0 ad=2.156p pd=7.14u as=0.728p ps=3.32u w=2.8u l=0.56u
X56 w_1750_n43456.t22 VINP.t10 a_8360_n43060.t13 w_1750_n43456.t21 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X57 a_8360_n43060.t8 VINP.t11 w_1750_n43456.t20 w_1750_n43456.t19 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X58 a_2044_n43060.t13 VINN.t8 w_1750_n43456.t61 w_1750_n43456.t60 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X59 w_1750_n43456.t63 VINN.t9 a_2044_n43060.t12 w_1750_n43456.t62 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X60 VDD.t27 IB.t16 OUT.t16 VDD.t26 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X61 OUT.t0 IB.t17 VDD.t25 VDD.t24 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X62 w_1750_n43456.t65 VINN.t10 a_2044_n43060.t11 w_1750_n43456.t64 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X63 a_8360_n43060.t4 VINP.t12 w_1750_n43456.t18 w_1750_n43456.t17 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X64 OUT.t5 IB.t18 VDD.t23 VDD.t22 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X65 OUT.t11 IB.t19 VDD.t21 VDD.t20 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X66 a_2044_n43060.t10 VINN.t11 w_1750_n43456.t67 w_1750_n43456.t66 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X67 OUT.t2 IB.t20 VDD.t19 VDD.t18 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X68 a_8360_n43060.t11 VINP.t13 w_1750_n43456.t16 w_1750_n43456.t15 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X69 a_2044_n43060.t9 VINN.t12 w_1750_n43456.t69 w_1750_n43456.t68 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X70 VDD.t17 IB.t21 a_n1924_n43526.t0 VDD.t16 pfet_06v0 ad=0.728p pd=3.32u as=2.156p ps=7.14u w=2.8u l=0.56u
X71 w_1750_n43456.t14 VINP.t14 a_8360_n43060.t14 w_1750_n43456.t13 pfet_06v0 ad=0.728p pd=3.32u as=2.156p ps=7.14u w=2.8u l=0.56u
X72 w_1750_n43456.t71 VINN.t13 a_2044_n43060.t8 w_1750_n43456.t70 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X73 VDD.t15 IB.t22 w_1750_n43456.t2 VDD.t14 pfet_06v0 ad=0.728p pd=3.32u as=2.156p ps=7.14u w=2.8u l=0.56u
X74 a_8360_n43060.t13 VINP.t15 w_1750_n43456.t12 w_1750_n43456.t11 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X75 OUT.t20 a_8360_n43060.t32 VSS.t15 VSS.t14 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X76 OUT.t39 IB.t23 VDD.t13 VDD.t12 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X77 a_8360_n43060.t0 a_n1924_n43526.t6 a_16582_n43566.t1 VSS.t0 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X78 w_1750_n43456.t10 VINP.t16 a_8360_n43060.t7 w_1750_n43456.t9 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X79 a_2044_n43060.t7 VINN.t14 w_1750_n43456.t73 w_1750_n43456.t72 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X80 OUT.t3 IB.t24 VDD.t11 VDD.t10 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X81 VSS.t13 a_8360_n43060.t33 OUT.t19 VSS.t12 nfet_06v0 ad=2.19p pd=7.46u as=0.78p ps=3.52u w=3u l=0.6u
X82 w_1750_n43456.t75 VINN.t15 a_2044_n43060.t6 w_1750_n43456.t74 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X83 VDD.t9 IB.t25 OUT.t15 VDD.t8 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X84 a_16582_n43566.t0 a_n1924_n43526.t7 a_8360_n43060.t0 VSS.t3 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X85 w_1750_n43456.t8 VINP.t17 a_8360_n43060.t12 w_1750_n43456.t7 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X86 w_1750_n43456.t6 VINP.t18 a_8360_n43060.t6 w_1750_n43456.t5 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X87 VDD.t7 IB.t26 OUT.t12 VDD.t6 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X88 w_1750_n43456.t77 VINN.t16 a_2044_n43060.t5 w_1750_n43456.t76 pfet_06v0 ad=0.728p pd=3.32u as=2.156p ps=7.14u w=2.8u l=0.56u
X89 a_2044_n43060.t4 VINN.t17 w_1750_n43456.t79 w_1750_n43456.t78 pfet_06v0 ad=2.156p pd=7.14u as=0.728p ps=3.32u w=2.8u l=0.56u
X90 VDD.t5 IB.t27 OUT.t4 VDD.t4 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X91 a_2044_n43060.t3 VINN.t18 w_1750_n43456.t81 w_1750_n43456.t80 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X92 w_1750_n43456.t43 IB.t28 VDD.t3 VDD.t2 pfet_06v0 ad=2.156p pd=7.14u as=0.728p ps=3.32u w=2.8u l=0.56u
X93 OUT.t18 a_8360_n43060.t34 VSS.t11 VSS.t10 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.6u
X94 w_1750_n43456.t4 VINP.t19 a_8360_n43060.t9 w_1750_n43456.t3 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X95 VDD.t1 IB.t29 OUT.t13 VDD.t0 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
X96 w_1750_n43456.t83 VINN.t19 a_2044_n43060.t2 w_1750_n43456.t82 pfet_06v0 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.56u
R0 a_8360_n43060.n1 a_8360_n43060.t33 45.7165
R1 a_8360_n43060.n2 a_8360_n43060.t19 45.5905
R2 a_8360_n43060.n2 a_8360_n43060.t26 45.5905
R3 a_8360_n43060.n2 a_8360_n43060.t34 45.5905
R4 a_8360_n43060.n2 a_8360_n43060.t25 45.5905
R5 a_8360_n43060.n2 a_8360_n43060.t29 45.5905
R6 a_8360_n43060.n2 a_8360_n43060.t18 45.5905
R7 a_8360_n43060.n2 a_8360_n43060.t21 45.5905
R8 a_8360_n43060.n2 a_8360_n43060.t31 45.5905
R9 a_8360_n43060.n2 a_8360_n43060.t24 45.5905
R10 a_8360_n43060.n2 a_8360_n43060.t28 45.5905
R11 a_8360_n43060.n2 a_8360_n43060.t17 45.5905
R12 a_8360_n43060.n2 a_8360_n43060.t20 45.5905
R13 a_8360_n43060.n1 a_8360_n43060.t30 45.5905
R14 a_8360_n43060.n1 a_8360_n43060.t23 45.5905
R15 a_8360_n43060.n1 a_8360_n43060.t27 45.5905
R16 a_8360_n43060.n1 a_8360_n43060.t16 45.5905
R17 a_8360_n43060.n1 a_8360_n43060.t22 45.5905
R18 a_8360_n43060.n1 a_8360_n43060.t15 45.5905
R19 a_8360_n43060.n1 a_8360_n43060.t32 45.5905
R20 a_8360_n43060.n0 a_8360_n43060.t1 10.3183
R21 a_8360_n43060.n0 a_8360_n43060.t10 9.50526
R22 a_8360_n43060.n0 a_8360_n43060.t14 9.32226
R23 a_8360_n43060.t4 a_8360_n43060.n0 7.97226
R24 a_8360_n43060.n0 a_8360_n43060.t9 7.97226
R25 a_8360_n43060.n0 a_8360_n43060.t13 7.97226
R26 a_8360_n43060.n0 a_8360_n43060.t6 7.97226
R27 a_8360_n43060.n0 a_8360_n43060.t11 7.97226
R28 a_8360_n43060.n0 a_8360_n43060.t8 7.97226
R29 a_8360_n43060.n0 a_8360_n43060.t7 7.97226
R30 a_8360_n43060.n0 a_8360_n43060.t5 7.97226
R31 a_8360_n43060.n0 a_8360_n43060.t12 7.97226
R32 a_8360_n43060.n3 a_8360_n43060.t3 7.22176
R33 a_8360_n43060.n3 a_8360_n43060.t2 7.03426
R34 a_8360_n43060.n3 a_8360_n43060.t0 5.94226
R35 a_8360_n43060.n0 a_8360_n43060.n4 5.34326
R36 a_8360_n43060.n4 a_8360_n43060.n3 2.51291
R37 a_8360_n43060.n2 a_8360_n43060.n1 2.26567
R38 a_8360_n43060.n4 a_8360_n43060.n2 2.24658
R39 OUT.n39 OUT.n38 17.1003
R40 OUT.n1 OUT.t9 9.50526
R41 OUT.n18 OUT.t14 9.32226
R42 OUT.n22 OUT.n20 8.35926
R43 OUT.n22 OUT.n21 8.19126
R44 OUT.n24 OUT.n23 8.19126
R45 OUT.n26 OUT.n25 8.19126
R46 OUT.n28 OUT.n27 8.19126
R47 OUT.n32 OUT.n31 8.19126
R48 OUT.n34 OUT.n33 8.19126
R49 OUT.n36 OUT.n35 8.19126
R50 OUT.n38 OUT.n37 8.19126
R51 OUT.n30 OUT.n29 8.18938
R52 OUT.n1 OUT.n0 7.97226
R53 OUT.n3 OUT.n2 7.97226
R54 OUT.n5 OUT.n4 7.97226
R55 OUT.n7 OUT.n6 7.97226
R56 OUT.n9 OUT.n8 7.97226
R57 OUT.n11 OUT.n10 7.97226
R58 OUT.n13 OUT.n12 7.97226
R59 OUT.n15 OUT.n14 7.97226
R60 OUT.n17 OUT.n16 7.97226
R61 OUT.n19 OUT.n18 3.98467
R62 OUT.n39 OUT.n19 3.4289
R63 OUT.n0 OUT.t1 0.6505
R64 OUT.n0 OUT.t6 0.6505
R65 OUT.n2 OUT.t38 0.6505
R66 OUT.n2 OUT.t11 0.6505
R67 OUT.n4 OUT.t17 0.6505
R68 OUT.n4 OUT.t2 0.6505
R69 OUT.n6 OUT.t15 0.6505
R70 OUT.n6 OUT.t39 0.6505
R71 OUT.n8 OUT.t12 0.6505
R72 OUT.n8 OUT.t0 0.6505
R73 OUT.n10 OUT.t7 0.6505
R74 OUT.n10 OUT.t5 0.6505
R75 OUT.n12 OUT.t4 0.6505
R76 OUT.n12 OUT.t8 0.6505
R77 OUT.n14 OUT.t13 0.6505
R78 OUT.n14 OUT.t10 0.6505
R79 OUT.n16 OUT.t16 0.6505
R80 OUT.n16 OUT.t3 0.6505
R81 OUT.n20 OUT.t26 0.5465
R82 OUT.n20 OUT.t33 0.5465
R83 OUT.n21 OUT.t27 0.5465
R84 OUT.n21 OUT.t18 0.5465
R85 OUT.n23 OUT.t34 0.5465
R86 OUT.n23 OUT.t23 0.5465
R87 OUT.n25 OUT.t21 0.5465
R88 OUT.n25 OUT.t31 0.5465
R89 OUT.n27 OUT.t24 0.5465
R90 OUT.n27 OUT.t28 0.5465
R91 OUT.n29 OUT.t32 0.5465
R92 OUT.n29 OUT.t35 0.5465
R93 OUT.n31 OUT.t29 0.5465
R94 OUT.n31 OUT.t22 0.5465
R95 OUT.n33 OUT.t36 0.5465
R96 OUT.n33 OUT.t25 0.5465
R97 OUT.n35 OUT.t37 0.5465
R98 OUT.n35 OUT.t30 0.5465
R99 OUT.n37 OUT.t19 0.5465
R100 OUT.n37 OUT.t20 0.5465
R101 OUT.n18 OUT.n17 0.1835
R102 OUT.n32 OUT.n30 0.16925
R103 OUT.n38 OUT.n36 0.1685
R104 OUT.n36 OUT.n34 0.1685
R105 OUT.n34 OUT.n32 0.1685
R106 OUT.n28 OUT.n26 0.1685
R107 OUT.n26 OUT.n24 0.1685
R108 OUT.n24 OUT.n22 0.1685
R109 OUT.n30 OUT.n28 0.16775
R110 OUT.n17 OUT.n15 0.1625
R111 OUT.n15 OUT.n13 0.1625
R112 OUT.n13 OUT.n11 0.1625
R113 OUT.n11 OUT.n9 0.1625
R114 OUT.n9 OUT.n7 0.1625
R115 OUT.n7 OUT.n5 0.1625
R116 OUT.n5 OUT.n3 0.1625
R117 OUT.n3 OUT.n1 0.1625
R118 OUT OUT.n39 0.04406
R119 OUT.n19 OUT.t40 0.00626923
R120 VSS.n1653 VSS.n895 69723.4
R121 VSS.n1755 VSS.n1654 6559.61
R122 VSS.n1653 VSS.n774 5526.89
R123 VSS.n3422 VSS.n895 1647.74
R124 VSS.n1654 VSS.n1653 947.068
R125 VSS.n3422 VSS.n896 549.845
R126 VSS.n1756 VSS.n1755 519.331
R127 VSS.n3405 VSS.t1 446.337
R128 VSS.n3508 VSS.n775 427.789
R129 VSS.t7 VSS.n775 415.824
R130 VSS.n3405 VSS.n774 396.079
R131 VSS.n4029 VSS.n705 324.303
R132 VSS.n705 VSS.n606 289.947
R133 VSS.n4158 VSS.n458 271.067
R134 VSS.n4026 VSS.n471 256.421
R135 VSS.n4144 VSS.n471 256.421
R136 VSS.n1756 VSS.n1699 226.161
R137 VSS.n3402 VSS.n896 195.647
R138 VSS.t1 VSS.n3402 183.083
R139 VSS.n1699 VSS.t7 183.083
R140 VSS.n895 VSS.n708 180.463
R141 VSS.n3424 VSS.n893 173.712
R142 VSS.n2187 VSS.n1622 169.013
R143 VSS.n1757 VSS.n1698 169.013
R144 VSS.n2238 VSS.n1623 154.922
R145 VSS.n4158 VSS.n459 147.554
R146 VSS.n3801 VSS.n3559 131.619
R147 VSS.n1925 VSS.n1621 127.013
R148 VSS.n2238 VSS.n1622 127.013
R149 VSS.n2106 VSS.n1619 127.013
R150 VSS.n3406 VSS.n897 127.013
R151 VSS.n1702 VSS.n1701 127.013
R152 VSS.n3404 VSS.n893 127.013
R153 VSS.n1758 VSS.n1757 127.013
R154 VSS.n2097 VSS.n1623 126.921
R155 VSS.n3509 VSS.n773 126.921
R156 VSS.n1703 VSS.n1698 126.921
R157 VSS.n4026 VSS.n710 126.921
R158 VSS.n3852 VSS.n3803 126.921
R159 VSS.n4160 VSS.n457 116.626
R160 VSS.n3421 VSS.n897 98.6452
R161 VSS.n3853 VSS.n3801 96.8952
R162 VSS.n1925 VSS.n1656 93.9479
R163 VSS.n1753 VSS.n1702 93.9479
R164 VSS.n3853 VSS.n3852 89.6189
R165 VSS.n1880 VSS.n1657 89.0663
R166 VSS.n2125 VSS.n2006 89.0663
R167 VSS.n3509 VSS.n772 89.0663
R168 VSS.n2185 VSS.n1618 81.2458
R169 VSS.n2106 VSS.n1657 79.9479
R170 VSS.n2005 VSS.n1621 79.8558
R171 VSS.n2185 VSS.n1654 78.625
R172 VSS.n4029 VSS.n706 78.5663
R173 VSS.n2239 VSS.n1620 66.9249
R174 VSS.n2006 VSS.n1619 65.8558
R175 VSS.n1701 VSS.n776 65.8558
R176 VSS.n1758 VSS.n772 65.8558
R177 VSS.n4028 VSS.n4027 65.0529
R178 VSS.t4 VSS.n2239 65.0529
R179 VSS.n3406 VSS.n776 61.1584
R180 VSS.n3404 VSS.n772 61.1584
R181 VSS.n3797 VSS.n3559 61.0663
R182 VSS.n1866 VSS.n1656 51.6716
R183 VSS.n2127 VSS.n2005 51.6716
R184 VSS.n2184 VSS.n1652 51.6716
R185 VSS.n3421 VSS.n894 51.6716
R186 VSS.n616 VSS.n606 51.6716
R187 VSS.n4147 VSS.n470 51.6716
R188 VSS.n3797 VSS.n459 45.1321
R189 VSS.n2242 VSS.n1618 35.3815
R190 VSS.n4028 VSS.n707 33.4159
R191 VSS.t40 VSS.n707 32.9479
R192 VSS.n4160 VSS.t12 28.6423
R193 VSS.n2242 VSS.t4 28.6423
R194 VSS.t12 VSS.t14 20.967
R195 VSS.t34 VSS.t48 20.967
R196 VSS.t46 VSS.t34 20.967
R197 VSS.t24 VSS.t46 20.967
R198 VSS.t32 VSS.t24 20.967
R199 VSS.t18 VSS.t38 20.967
R200 VSS.t38 VSS.t44 20.967
R201 VSS.t30 VSS.t22 20.967
R202 VSS.t16 VSS.t36 20.967
R203 VSS.t36 VSS.t42 20.967
R204 VSS.t20 VSS.t9 20.4054
R205 VSS.t28 VSS.t3 20.4054
R206 VSS.t26 VSS.t6 20.4054
R207 VSS.n4146 VSS.t22 20.031
R208 VSS.t14 VSS.n4159 18.7206
R209 VSS.n3560 VSS.t0 17.1294
R210 VSS.n3796 VSS.t16 16.0998
R211 VSS.n2099 VSS.n2006 14.0005
R212 VSS.n2184 VSS.n1657 14.0005
R213 VSS.n3506 VSS.n776 14.0005
R214 VSS.n3854 VSS.n3853 14.0005
R215 VSS.n4147 VSS.n459 14.0005
R216 VSS.n704 VSS.t18 11.607
R217 VSS.n3206 VSS.n1375 9.92188
R218 VSS.n2243 VSS.n1375 9.86
R219 VSS.n704 VSS.t32 9.36056
R220 VSS.n3795 VSS.n3794 8.70536
R221 VSS.n3794 VSS.t20 8.23735
R222 VSS.n4162 VSS.t41 7.22413
R223 VSS.n4162 VSS.n4161 5.94463
R224 VSS.n4164 VSS.n4163 5.94463
R225 VSS.n4166 VSS.n4165 5.94463
R226 VSS.n4168 VSS.n4167 5.94463
R227 VSS.n4170 VSS.n4169 5.94463
R228 VSS.n4174 VSS.n4173 5.94463
R229 VSS.n4176 VSS.n4175 5.94463
R230 VSS.n4178 VSS.n4177 5.94463
R231 VSS.n4172 VSS.n4171 5.94275
R232 VSS.n2241 VSS.t5 4.96786
R233 VSS.n3796 VSS.t30 4.86773
R234 VSS.n4179 VSS.t13 4.75524
R235 VSS.n1030 VSS.t8 4.74785
R236 VSS.n3401 VSS.t2 4.74752
R237 VSS.n4503 VSS.n4502 4.5005
R238 VSS.n4504 VSS.n4503 4.5005
R239 VSS.n4504 VSS.n383 4.5005
R240 VSS.n193 VSS.n69 4.5005
R241 VSS.n195 VSS.n69 4.5005
R242 VSS.n192 VSS.n69 4.5005
R243 VSS.n196 VSS.n69 4.5005
R244 VSS.n191 VSS.n69 4.5005
R245 VSS.n197 VSS.n69 4.5005
R246 VSS.n190 VSS.n69 4.5005
R247 VSS.n198 VSS.n69 4.5005
R248 VSS.n189 VSS.n69 4.5005
R249 VSS.n199 VSS.n69 4.5005
R250 VSS.n188 VSS.n69 4.5005
R251 VSS.n200 VSS.n69 4.5005
R252 VSS.n187 VSS.n69 4.5005
R253 VSS.n201 VSS.n69 4.5005
R254 VSS.n186 VSS.n69 4.5005
R255 VSS.n202 VSS.n69 4.5005
R256 VSS.n185 VSS.n69 4.5005
R257 VSS.n203 VSS.n69 4.5005
R258 VSS.n184 VSS.n69 4.5005
R259 VSS.n204 VSS.n69 4.5005
R260 VSS.n183 VSS.n69 4.5005
R261 VSS.n205 VSS.n69 4.5005
R262 VSS.n182 VSS.n69 4.5005
R263 VSS.n206 VSS.n69 4.5005
R264 VSS.n181 VSS.n69 4.5005
R265 VSS.n207 VSS.n69 4.5005
R266 VSS.n180 VSS.n69 4.5005
R267 VSS.n208 VSS.n69 4.5005
R268 VSS.n179 VSS.n69 4.5005
R269 VSS.n209 VSS.n69 4.5005
R270 VSS.n178 VSS.n69 4.5005
R271 VSS.n210 VSS.n69 4.5005
R272 VSS.n177 VSS.n69 4.5005
R273 VSS.n211 VSS.n69 4.5005
R274 VSS.n176 VSS.n69 4.5005
R275 VSS.n212 VSS.n69 4.5005
R276 VSS.n175 VSS.n69 4.5005
R277 VSS.n213 VSS.n69 4.5005
R278 VSS.n174 VSS.n69 4.5005
R279 VSS.n214 VSS.n69 4.5005
R280 VSS.n173 VSS.n69 4.5005
R281 VSS.n215 VSS.n69 4.5005
R282 VSS.n172 VSS.n69 4.5005
R283 VSS.n216 VSS.n69 4.5005
R284 VSS.n171 VSS.n69 4.5005
R285 VSS.n217 VSS.n69 4.5005
R286 VSS.n170 VSS.n69 4.5005
R287 VSS.n218 VSS.n69 4.5005
R288 VSS.n169 VSS.n69 4.5005
R289 VSS.n219 VSS.n69 4.5005
R290 VSS.n168 VSS.n69 4.5005
R291 VSS.n220 VSS.n69 4.5005
R292 VSS.n167 VSS.n69 4.5005
R293 VSS.n221 VSS.n69 4.5005
R294 VSS.n166 VSS.n69 4.5005
R295 VSS.n222 VSS.n69 4.5005
R296 VSS.n165 VSS.n69 4.5005
R297 VSS.n223 VSS.n69 4.5005
R298 VSS.n164 VSS.n69 4.5005
R299 VSS.n224 VSS.n69 4.5005
R300 VSS.n163 VSS.n69 4.5005
R301 VSS.n225 VSS.n69 4.5005
R302 VSS.n162 VSS.n69 4.5005
R303 VSS.n226 VSS.n69 4.5005
R304 VSS.n161 VSS.n69 4.5005
R305 VSS.n227 VSS.n69 4.5005
R306 VSS.n160 VSS.n69 4.5005
R307 VSS.n228 VSS.n69 4.5005
R308 VSS.n159 VSS.n69 4.5005
R309 VSS.n229 VSS.n69 4.5005
R310 VSS.n158 VSS.n69 4.5005
R311 VSS.n230 VSS.n69 4.5005
R312 VSS.n157 VSS.n69 4.5005
R313 VSS.n231 VSS.n69 4.5005
R314 VSS.n156 VSS.n69 4.5005
R315 VSS.n232 VSS.n69 4.5005
R316 VSS.n155 VSS.n69 4.5005
R317 VSS.n233 VSS.n69 4.5005
R318 VSS.n154 VSS.n69 4.5005
R319 VSS.n234 VSS.n69 4.5005
R320 VSS.n153 VSS.n69 4.5005
R321 VSS.n235 VSS.n69 4.5005
R322 VSS.n4506 VSS.n69 4.5005
R323 VSS.n236 VSS.n69 4.5005
R324 VSS.n152 VSS.n69 4.5005
R325 VSS.n237 VSS.n69 4.5005
R326 VSS.n151 VSS.n69 4.5005
R327 VSS.n238 VSS.n69 4.5005
R328 VSS.n150 VSS.n69 4.5005
R329 VSS.n239 VSS.n69 4.5005
R330 VSS.n149 VSS.n69 4.5005
R331 VSS.n240 VSS.n69 4.5005
R332 VSS.n148 VSS.n69 4.5005
R333 VSS.n241 VSS.n69 4.5005
R334 VSS.n147 VSS.n69 4.5005
R335 VSS.n242 VSS.n69 4.5005
R336 VSS.n146 VSS.n69 4.5005
R337 VSS.n243 VSS.n69 4.5005
R338 VSS.n145 VSS.n69 4.5005
R339 VSS.n244 VSS.n69 4.5005
R340 VSS.n144 VSS.n69 4.5005
R341 VSS.n245 VSS.n69 4.5005
R342 VSS.n143 VSS.n69 4.5005
R343 VSS.n246 VSS.n69 4.5005
R344 VSS.n142 VSS.n69 4.5005
R345 VSS.n247 VSS.n69 4.5005
R346 VSS.n141 VSS.n69 4.5005
R347 VSS.n248 VSS.n69 4.5005
R348 VSS.n140 VSS.n69 4.5005
R349 VSS.n249 VSS.n69 4.5005
R350 VSS.n139 VSS.n69 4.5005
R351 VSS.n250 VSS.n69 4.5005
R352 VSS.n138 VSS.n69 4.5005
R353 VSS.n251 VSS.n69 4.5005
R354 VSS.n137 VSS.n69 4.5005
R355 VSS.n252 VSS.n69 4.5005
R356 VSS.n136 VSS.n69 4.5005
R357 VSS.n253 VSS.n69 4.5005
R358 VSS.n135 VSS.n69 4.5005
R359 VSS.n254 VSS.n69 4.5005
R360 VSS.n134 VSS.n69 4.5005
R361 VSS.n255 VSS.n69 4.5005
R362 VSS.n133 VSS.n69 4.5005
R363 VSS.n256 VSS.n69 4.5005
R364 VSS.n132 VSS.n69 4.5005
R365 VSS.n4502 VSS.n69 4.5005
R366 VSS.n4504 VSS.n69 4.5005
R367 VSS.n193 VSS.n67 4.5005
R368 VSS.n195 VSS.n67 4.5005
R369 VSS.n192 VSS.n67 4.5005
R370 VSS.n196 VSS.n67 4.5005
R371 VSS.n191 VSS.n67 4.5005
R372 VSS.n197 VSS.n67 4.5005
R373 VSS.n190 VSS.n67 4.5005
R374 VSS.n198 VSS.n67 4.5005
R375 VSS.n189 VSS.n67 4.5005
R376 VSS.n199 VSS.n67 4.5005
R377 VSS.n188 VSS.n67 4.5005
R378 VSS.n200 VSS.n67 4.5005
R379 VSS.n187 VSS.n67 4.5005
R380 VSS.n201 VSS.n67 4.5005
R381 VSS.n186 VSS.n67 4.5005
R382 VSS.n202 VSS.n67 4.5005
R383 VSS.n185 VSS.n67 4.5005
R384 VSS.n203 VSS.n67 4.5005
R385 VSS.n184 VSS.n67 4.5005
R386 VSS.n204 VSS.n67 4.5005
R387 VSS.n183 VSS.n67 4.5005
R388 VSS.n205 VSS.n67 4.5005
R389 VSS.n182 VSS.n67 4.5005
R390 VSS.n206 VSS.n67 4.5005
R391 VSS.n181 VSS.n67 4.5005
R392 VSS.n207 VSS.n67 4.5005
R393 VSS.n180 VSS.n67 4.5005
R394 VSS.n208 VSS.n67 4.5005
R395 VSS.n179 VSS.n67 4.5005
R396 VSS.n209 VSS.n67 4.5005
R397 VSS.n178 VSS.n67 4.5005
R398 VSS.n210 VSS.n67 4.5005
R399 VSS.n177 VSS.n67 4.5005
R400 VSS.n211 VSS.n67 4.5005
R401 VSS.n176 VSS.n67 4.5005
R402 VSS.n212 VSS.n67 4.5005
R403 VSS.n175 VSS.n67 4.5005
R404 VSS.n213 VSS.n67 4.5005
R405 VSS.n174 VSS.n67 4.5005
R406 VSS.n214 VSS.n67 4.5005
R407 VSS.n173 VSS.n67 4.5005
R408 VSS.n215 VSS.n67 4.5005
R409 VSS.n172 VSS.n67 4.5005
R410 VSS.n216 VSS.n67 4.5005
R411 VSS.n171 VSS.n67 4.5005
R412 VSS.n217 VSS.n67 4.5005
R413 VSS.n170 VSS.n67 4.5005
R414 VSS.n218 VSS.n67 4.5005
R415 VSS.n169 VSS.n67 4.5005
R416 VSS.n219 VSS.n67 4.5005
R417 VSS.n168 VSS.n67 4.5005
R418 VSS.n220 VSS.n67 4.5005
R419 VSS.n167 VSS.n67 4.5005
R420 VSS.n221 VSS.n67 4.5005
R421 VSS.n166 VSS.n67 4.5005
R422 VSS.n222 VSS.n67 4.5005
R423 VSS.n165 VSS.n67 4.5005
R424 VSS.n223 VSS.n67 4.5005
R425 VSS.n164 VSS.n67 4.5005
R426 VSS.n224 VSS.n67 4.5005
R427 VSS.n163 VSS.n67 4.5005
R428 VSS.n225 VSS.n67 4.5005
R429 VSS.n162 VSS.n67 4.5005
R430 VSS.n226 VSS.n67 4.5005
R431 VSS.n161 VSS.n67 4.5005
R432 VSS.n227 VSS.n67 4.5005
R433 VSS.n160 VSS.n67 4.5005
R434 VSS.n228 VSS.n67 4.5005
R435 VSS.n159 VSS.n67 4.5005
R436 VSS.n229 VSS.n67 4.5005
R437 VSS.n158 VSS.n67 4.5005
R438 VSS.n230 VSS.n67 4.5005
R439 VSS.n157 VSS.n67 4.5005
R440 VSS.n231 VSS.n67 4.5005
R441 VSS.n156 VSS.n67 4.5005
R442 VSS.n232 VSS.n67 4.5005
R443 VSS.n155 VSS.n67 4.5005
R444 VSS.n233 VSS.n67 4.5005
R445 VSS.n154 VSS.n67 4.5005
R446 VSS.n234 VSS.n67 4.5005
R447 VSS.n153 VSS.n67 4.5005
R448 VSS.n235 VSS.n67 4.5005
R449 VSS.n4506 VSS.n67 4.5005
R450 VSS.n236 VSS.n67 4.5005
R451 VSS.n152 VSS.n67 4.5005
R452 VSS.n237 VSS.n67 4.5005
R453 VSS.n151 VSS.n67 4.5005
R454 VSS.n238 VSS.n67 4.5005
R455 VSS.n150 VSS.n67 4.5005
R456 VSS.n239 VSS.n67 4.5005
R457 VSS.n149 VSS.n67 4.5005
R458 VSS.n240 VSS.n67 4.5005
R459 VSS.n148 VSS.n67 4.5005
R460 VSS.n241 VSS.n67 4.5005
R461 VSS.n147 VSS.n67 4.5005
R462 VSS.n242 VSS.n67 4.5005
R463 VSS.n146 VSS.n67 4.5005
R464 VSS.n243 VSS.n67 4.5005
R465 VSS.n145 VSS.n67 4.5005
R466 VSS.n244 VSS.n67 4.5005
R467 VSS.n144 VSS.n67 4.5005
R468 VSS.n245 VSS.n67 4.5005
R469 VSS.n143 VSS.n67 4.5005
R470 VSS.n246 VSS.n67 4.5005
R471 VSS.n142 VSS.n67 4.5005
R472 VSS.n247 VSS.n67 4.5005
R473 VSS.n141 VSS.n67 4.5005
R474 VSS.n248 VSS.n67 4.5005
R475 VSS.n140 VSS.n67 4.5005
R476 VSS.n249 VSS.n67 4.5005
R477 VSS.n139 VSS.n67 4.5005
R478 VSS.n250 VSS.n67 4.5005
R479 VSS.n138 VSS.n67 4.5005
R480 VSS.n251 VSS.n67 4.5005
R481 VSS.n137 VSS.n67 4.5005
R482 VSS.n252 VSS.n67 4.5005
R483 VSS.n136 VSS.n67 4.5005
R484 VSS.n253 VSS.n67 4.5005
R485 VSS.n135 VSS.n67 4.5005
R486 VSS.n254 VSS.n67 4.5005
R487 VSS.n134 VSS.n67 4.5005
R488 VSS.n255 VSS.n67 4.5005
R489 VSS.n133 VSS.n67 4.5005
R490 VSS.n256 VSS.n67 4.5005
R491 VSS.n132 VSS.n67 4.5005
R492 VSS.n4502 VSS.n67 4.5005
R493 VSS.n4504 VSS.n67 4.5005
R494 VSS.n193 VSS.n70 4.5005
R495 VSS.n195 VSS.n70 4.5005
R496 VSS.n192 VSS.n70 4.5005
R497 VSS.n196 VSS.n70 4.5005
R498 VSS.n191 VSS.n70 4.5005
R499 VSS.n197 VSS.n70 4.5005
R500 VSS.n190 VSS.n70 4.5005
R501 VSS.n198 VSS.n70 4.5005
R502 VSS.n189 VSS.n70 4.5005
R503 VSS.n199 VSS.n70 4.5005
R504 VSS.n188 VSS.n70 4.5005
R505 VSS.n200 VSS.n70 4.5005
R506 VSS.n187 VSS.n70 4.5005
R507 VSS.n201 VSS.n70 4.5005
R508 VSS.n186 VSS.n70 4.5005
R509 VSS.n202 VSS.n70 4.5005
R510 VSS.n185 VSS.n70 4.5005
R511 VSS.n203 VSS.n70 4.5005
R512 VSS.n184 VSS.n70 4.5005
R513 VSS.n204 VSS.n70 4.5005
R514 VSS.n183 VSS.n70 4.5005
R515 VSS.n205 VSS.n70 4.5005
R516 VSS.n182 VSS.n70 4.5005
R517 VSS.n206 VSS.n70 4.5005
R518 VSS.n181 VSS.n70 4.5005
R519 VSS.n207 VSS.n70 4.5005
R520 VSS.n180 VSS.n70 4.5005
R521 VSS.n208 VSS.n70 4.5005
R522 VSS.n179 VSS.n70 4.5005
R523 VSS.n209 VSS.n70 4.5005
R524 VSS.n178 VSS.n70 4.5005
R525 VSS.n210 VSS.n70 4.5005
R526 VSS.n177 VSS.n70 4.5005
R527 VSS.n211 VSS.n70 4.5005
R528 VSS.n176 VSS.n70 4.5005
R529 VSS.n212 VSS.n70 4.5005
R530 VSS.n175 VSS.n70 4.5005
R531 VSS.n213 VSS.n70 4.5005
R532 VSS.n174 VSS.n70 4.5005
R533 VSS.n214 VSS.n70 4.5005
R534 VSS.n173 VSS.n70 4.5005
R535 VSS.n215 VSS.n70 4.5005
R536 VSS.n172 VSS.n70 4.5005
R537 VSS.n216 VSS.n70 4.5005
R538 VSS.n171 VSS.n70 4.5005
R539 VSS.n217 VSS.n70 4.5005
R540 VSS.n170 VSS.n70 4.5005
R541 VSS.n218 VSS.n70 4.5005
R542 VSS.n169 VSS.n70 4.5005
R543 VSS.n219 VSS.n70 4.5005
R544 VSS.n168 VSS.n70 4.5005
R545 VSS.n220 VSS.n70 4.5005
R546 VSS.n167 VSS.n70 4.5005
R547 VSS.n221 VSS.n70 4.5005
R548 VSS.n166 VSS.n70 4.5005
R549 VSS.n222 VSS.n70 4.5005
R550 VSS.n165 VSS.n70 4.5005
R551 VSS.n223 VSS.n70 4.5005
R552 VSS.n164 VSS.n70 4.5005
R553 VSS.n224 VSS.n70 4.5005
R554 VSS.n163 VSS.n70 4.5005
R555 VSS.n225 VSS.n70 4.5005
R556 VSS.n162 VSS.n70 4.5005
R557 VSS.n226 VSS.n70 4.5005
R558 VSS.n161 VSS.n70 4.5005
R559 VSS.n227 VSS.n70 4.5005
R560 VSS.n160 VSS.n70 4.5005
R561 VSS.n228 VSS.n70 4.5005
R562 VSS.n159 VSS.n70 4.5005
R563 VSS.n229 VSS.n70 4.5005
R564 VSS.n158 VSS.n70 4.5005
R565 VSS.n230 VSS.n70 4.5005
R566 VSS.n157 VSS.n70 4.5005
R567 VSS.n231 VSS.n70 4.5005
R568 VSS.n156 VSS.n70 4.5005
R569 VSS.n232 VSS.n70 4.5005
R570 VSS.n155 VSS.n70 4.5005
R571 VSS.n233 VSS.n70 4.5005
R572 VSS.n154 VSS.n70 4.5005
R573 VSS.n234 VSS.n70 4.5005
R574 VSS.n153 VSS.n70 4.5005
R575 VSS.n235 VSS.n70 4.5005
R576 VSS.n4506 VSS.n70 4.5005
R577 VSS.n236 VSS.n70 4.5005
R578 VSS.n152 VSS.n70 4.5005
R579 VSS.n237 VSS.n70 4.5005
R580 VSS.n151 VSS.n70 4.5005
R581 VSS.n238 VSS.n70 4.5005
R582 VSS.n150 VSS.n70 4.5005
R583 VSS.n239 VSS.n70 4.5005
R584 VSS.n149 VSS.n70 4.5005
R585 VSS.n240 VSS.n70 4.5005
R586 VSS.n148 VSS.n70 4.5005
R587 VSS.n241 VSS.n70 4.5005
R588 VSS.n147 VSS.n70 4.5005
R589 VSS.n242 VSS.n70 4.5005
R590 VSS.n146 VSS.n70 4.5005
R591 VSS.n243 VSS.n70 4.5005
R592 VSS.n145 VSS.n70 4.5005
R593 VSS.n244 VSS.n70 4.5005
R594 VSS.n144 VSS.n70 4.5005
R595 VSS.n245 VSS.n70 4.5005
R596 VSS.n143 VSS.n70 4.5005
R597 VSS.n246 VSS.n70 4.5005
R598 VSS.n142 VSS.n70 4.5005
R599 VSS.n247 VSS.n70 4.5005
R600 VSS.n141 VSS.n70 4.5005
R601 VSS.n248 VSS.n70 4.5005
R602 VSS.n140 VSS.n70 4.5005
R603 VSS.n249 VSS.n70 4.5005
R604 VSS.n139 VSS.n70 4.5005
R605 VSS.n250 VSS.n70 4.5005
R606 VSS.n138 VSS.n70 4.5005
R607 VSS.n251 VSS.n70 4.5005
R608 VSS.n137 VSS.n70 4.5005
R609 VSS.n252 VSS.n70 4.5005
R610 VSS.n136 VSS.n70 4.5005
R611 VSS.n253 VSS.n70 4.5005
R612 VSS.n135 VSS.n70 4.5005
R613 VSS.n254 VSS.n70 4.5005
R614 VSS.n134 VSS.n70 4.5005
R615 VSS.n255 VSS.n70 4.5005
R616 VSS.n133 VSS.n70 4.5005
R617 VSS.n256 VSS.n70 4.5005
R618 VSS.n132 VSS.n70 4.5005
R619 VSS.n4502 VSS.n70 4.5005
R620 VSS.n4504 VSS.n70 4.5005
R621 VSS.n193 VSS.n66 4.5005
R622 VSS.n195 VSS.n66 4.5005
R623 VSS.n192 VSS.n66 4.5005
R624 VSS.n196 VSS.n66 4.5005
R625 VSS.n191 VSS.n66 4.5005
R626 VSS.n197 VSS.n66 4.5005
R627 VSS.n190 VSS.n66 4.5005
R628 VSS.n198 VSS.n66 4.5005
R629 VSS.n189 VSS.n66 4.5005
R630 VSS.n199 VSS.n66 4.5005
R631 VSS.n188 VSS.n66 4.5005
R632 VSS.n200 VSS.n66 4.5005
R633 VSS.n187 VSS.n66 4.5005
R634 VSS.n201 VSS.n66 4.5005
R635 VSS.n186 VSS.n66 4.5005
R636 VSS.n202 VSS.n66 4.5005
R637 VSS.n185 VSS.n66 4.5005
R638 VSS.n203 VSS.n66 4.5005
R639 VSS.n184 VSS.n66 4.5005
R640 VSS.n204 VSS.n66 4.5005
R641 VSS.n183 VSS.n66 4.5005
R642 VSS.n205 VSS.n66 4.5005
R643 VSS.n182 VSS.n66 4.5005
R644 VSS.n206 VSS.n66 4.5005
R645 VSS.n181 VSS.n66 4.5005
R646 VSS.n207 VSS.n66 4.5005
R647 VSS.n180 VSS.n66 4.5005
R648 VSS.n208 VSS.n66 4.5005
R649 VSS.n179 VSS.n66 4.5005
R650 VSS.n209 VSS.n66 4.5005
R651 VSS.n178 VSS.n66 4.5005
R652 VSS.n210 VSS.n66 4.5005
R653 VSS.n177 VSS.n66 4.5005
R654 VSS.n211 VSS.n66 4.5005
R655 VSS.n176 VSS.n66 4.5005
R656 VSS.n212 VSS.n66 4.5005
R657 VSS.n175 VSS.n66 4.5005
R658 VSS.n213 VSS.n66 4.5005
R659 VSS.n174 VSS.n66 4.5005
R660 VSS.n214 VSS.n66 4.5005
R661 VSS.n173 VSS.n66 4.5005
R662 VSS.n215 VSS.n66 4.5005
R663 VSS.n172 VSS.n66 4.5005
R664 VSS.n216 VSS.n66 4.5005
R665 VSS.n171 VSS.n66 4.5005
R666 VSS.n217 VSS.n66 4.5005
R667 VSS.n170 VSS.n66 4.5005
R668 VSS.n218 VSS.n66 4.5005
R669 VSS.n169 VSS.n66 4.5005
R670 VSS.n219 VSS.n66 4.5005
R671 VSS.n168 VSS.n66 4.5005
R672 VSS.n220 VSS.n66 4.5005
R673 VSS.n167 VSS.n66 4.5005
R674 VSS.n221 VSS.n66 4.5005
R675 VSS.n166 VSS.n66 4.5005
R676 VSS.n222 VSS.n66 4.5005
R677 VSS.n165 VSS.n66 4.5005
R678 VSS.n223 VSS.n66 4.5005
R679 VSS.n164 VSS.n66 4.5005
R680 VSS.n224 VSS.n66 4.5005
R681 VSS.n163 VSS.n66 4.5005
R682 VSS.n225 VSS.n66 4.5005
R683 VSS.n162 VSS.n66 4.5005
R684 VSS.n226 VSS.n66 4.5005
R685 VSS.n161 VSS.n66 4.5005
R686 VSS.n227 VSS.n66 4.5005
R687 VSS.n160 VSS.n66 4.5005
R688 VSS.n228 VSS.n66 4.5005
R689 VSS.n159 VSS.n66 4.5005
R690 VSS.n229 VSS.n66 4.5005
R691 VSS.n158 VSS.n66 4.5005
R692 VSS.n230 VSS.n66 4.5005
R693 VSS.n157 VSS.n66 4.5005
R694 VSS.n231 VSS.n66 4.5005
R695 VSS.n156 VSS.n66 4.5005
R696 VSS.n232 VSS.n66 4.5005
R697 VSS.n155 VSS.n66 4.5005
R698 VSS.n233 VSS.n66 4.5005
R699 VSS.n154 VSS.n66 4.5005
R700 VSS.n234 VSS.n66 4.5005
R701 VSS.n153 VSS.n66 4.5005
R702 VSS.n235 VSS.n66 4.5005
R703 VSS.n4506 VSS.n66 4.5005
R704 VSS.n236 VSS.n66 4.5005
R705 VSS.n152 VSS.n66 4.5005
R706 VSS.n237 VSS.n66 4.5005
R707 VSS.n151 VSS.n66 4.5005
R708 VSS.n238 VSS.n66 4.5005
R709 VSS.n150 VSS.n66 4.5005
R710 VSS.n239 VSS.n66 4.5005
R711 VSS.n149 VSS.n66 4.5005
R712 VSS.n240 VSS.n66 4.5005
R713 VSS.n148 VSS.n66 4.5005
R714 VSS.n241 VSS.n66 4.5005
R715 VSS.n147 VSS.n66 4.5005
R716 VSS.n242 VSS.n66 4.5005
R717 VSS.n146 VSS.n66 4.5005
R718 VSS.n243 VSS.n66 4.5005
R719 VSS.n145 VSS.n66 4.5005
R720 VSS.n244 VSS.n66 4.5005
R721 VSS.n144 VSS.n66 4.5005
R722 VSS.n245 VSS.n66 4.5005
R723 VSS.n143 VSS.n66 4.5005
R724 VSS.n246 VSS.n66 4.5005
R725 VSS.n142 VSS.n66 4.5005
R726 VSS.n247 VSS.n66 4.5005
R727 VSS.n141 VSS.n66 4.5005
R728 VSS.n248 VSS.n66 4.5005
R729 VSS.n140 VSS.n66 4.5005
R730 VSS.n249 VSS.n66 4.5005
R731 VSS.n139 VSS.n66 4.5005
R732 VSS.n250 VSS.n66 4.5005
R733 VSS.n138 VSS.n66 4.5005
R734 VSS.n251 VSS.n66 4.5005
R735 VSS.n137 VSS.n66 4.5005
R736 VSS.n252 VSS.n66 4.5005
R737 VSS.n136 VSS.n66 4.5005
R738 VSS.n253 VSS.n66 4.5005
R739 VSS.n135 VSS.n66 4.5005
R740 VSS.n254 VSS.n66 4.5005
R741 VSS.n134 VSS.n66 4.5005
R742 VSS.n255 VSS.n66 4.5005
R743 VSS.n133 VSS.n66 4.5005
R744 VSS.n256 VSS.n66 4.5005
R745 VSS.n132 VSS.n66 4.5005
R746 VSS.n4502 VSS.n66 4.5005
R747 VSS.n4504 VSS.n66 4.5005
R748 VSS.n193 VSS.n71 4.5005
R749 VSS.n195 VSS.n71 4.5005
R750 VSS.n192 VSS.n71 4.5005
R751 VSS.n196 VSS.n71 4.5005
R752 VSS.n191 VSS.n71 4.5005
R753 VSS.n197 VSS.n71 4.5005
R754 VSS.n190 VSS.n71 4.5005
R755 VSS.n198 VSS.n71 4.5005
R756 VSS.n189 VSS.n71 4.5005
R757 VSS.n199 VSS.n71 4.5005
R758 VSS.n188 VSS.n71 4.5005
R759 VSS.n200 VSS.n71 4.5005
R760 VSS.n187 VSS.n71 4.5005
R761 VSS.n201 VSS.n71 4.5005
R762 VSS.n186 VSS.n71 4.5005
R763 VSS.n202 VSS.n71 4.5005
R764 VSS.n185 VSS.n71 4.5005
R765 VSS.n203 VSS.n71 4.5005
R766 VSS.n184 VSS.n71 4.5005
R767 VSS.n204 VSS.n71 4.5005
R768 VSS.n183 VSS.n71 4.5005
R769 VSS.n205 VSS.n71 4.5005
R770 VSS.n182 VSS.n71 4.5005
R771 VSS.n206 VSS.n71 4.5005
R772 VSS.n181 VSS.n71 4.5005
R773 VSS.n207 VSS.n71 4.5005
R774 VSS.n180 VSS.n71 4.5005
R775 VSS.n208 VSS.n71 4.5005
R776 VSS.n179 VSS.n71 4.5005
R777 VSS.n209 VSS.n71 4.5005
R778 VSS.n178 VSS.n71 4.5005
R779 VSS.n210 VSS.n71 4.5005
R780 VSS.n177 VSS.n71 4.5005
R781 VSS.n211 VSS.n71 4.5005
R782 VSS.n176 VSS.n71 4.5005
R783 VSS.n212 VSS.n71 4.5005
R784 VSS.n175 VSS.n71 4.5005
R785 VSS.n213 VSS.n71 4.5005
R786 VSS.n174 VSS.n71 4.5005
R787 VSS.n214 VSS.n71 4.5005
R788 VSS.n173 VSS.n71 4.5005
R789 VSS.n215 VSS.n71 4.5005
R790 VSS.n172 VSS.n71 4.5005
R791 VSS.n216 VSS.n71 4.5005
R792 VSS.n171 VSS.n71 4.5005
R793 VSS.n217 VSS.n71 4.5005
R794 VSS.n170 VSS.n71 4.5005
R795 VSS.n218 VSS.n71 4.5005
R796 VSS.n169 VSS.n71 4.5005
R797 VSS.n219 VSS.n71 4.5005
R798 VSS.n168 VSS.n71 4.5005
R799 VSS.n220 VSS.n71 4.5005
R800 VSS.n167 VSS.n71 4.5005
R801 VSS.n221 VSS.n71 4.5005
R802 VSS.n166 VSS.n71 4.5005
R803 VSS.n222 VSS.n71 4.5005
R804 VSS.n165 VSS.n71 4.5005
R805 VSS.n223 VSS.n71 4.5005
R806 VSS.n164 VSS.n71 4.5005
R807 VSS.n224 VSS.n71 4.5005
R808 VSS.n163 VSS.n71 4.5005
R809 VSS.n225 VSS.n71 4.5005
R810 VSS.n162 VSS.n71 4.5005
R811 VSS.n226 VSS.n71 4.5005
R812 VSS.n161 VSS.n71 4.5005
R813 VSS.n227 VSS.n71 4.5005
R814 VSS.n160 VSS.n71 4.5005
R815 VSS.n228 VSS.n71 4.5005
R816 VSS.n159 VSS.n71 4.5005
R817 VSS.n229 VSS.n71 4.5005
R818 VSS.n158 VSS.n71 4.5005
R819 VSS.n230 VSS.n71 4.5005
R820 VSS.n157 VSS.n71 4.5005
R821 VSS.n231 VSS.n71 4.5005
R822 VSS.n156 VSS.n71 4.5005
R823 VSS.n232 VSS.n71 4.5005
R824 VSS.n155 VSS.n71 4.5005
R825 VSS.n233 VSS.n71 4.5005
R826 VSS.n154 VSS.n71 4.5005
R827 VSS.n234 VSS.n71 4.5005
R828 VSS.n153 VSS.n71 4.5005
R829 VSS.n235 VSS.n71 4.5005
R830 VSS.n4506 VSS.n71 4.5005
R831 VSS.n236 VSS.n71 4.5005
R832 VSS.n152 VSS.n71 4.5005
R833 VSS.n237 VSS.n71 4.5005
R834 VSS.n151 VSS.n71 4.5005
R835 VSS.n238 VSS.n71 4.5005
R836 VSS.n150 VSS.n71 4.5005
R837 VSS.n239 VSS.n71 4.5005
R838 VSS.n149 VSS.n71 4.5005
R839 VSS.n240 VSS.n71 4.5005
R840 VSS.n148 VSS.n71 4.5005
R841 VSS.n241 VSS.n71 4.5005
R842 VSS.n147 VSS.n71 4.5005
R843 VSS.n242 VSS.n71 4.5005
R844 VSS.n146 VSS.n71 4.5005
R845 VSS.n243 VSS.n71 4.5005
R846 VSS.n145 VSS.n71 4.5005
R847 VSS.n244 VSS.n71 4.5005
R848 VSS.n144 VSS.n71 4.5005
R849 VSS.n245 VSS.n71 4.5005
R850 VSS.n143 VSS.n71 4.5005
R851 VSS.n246 VSS.n71 4.5005
R852 VSS.n142 VSS.n71 4.5005
R853 VSS.n247 VSS.n71 4.5005
R854 VSS.n141 VSS.n71 4.5005
R855 VSS.n248 VSS.n71 4.5005
R856 VSS.n140 VSS.n71 4.5005
R857 VSS.n249 VSS.n71 4.5005
R858 VSS.n139 VSS.n71 4.5005
R859 VSS.n250 VSS.n71 4.5005
R860 VSS.n138 VSS.n71 4.5005
R861 VSS.n251 VSS.n71 4.5005
R862 VSS.n137 VSS.n71 4.5005
R863 VSS.n252 VSS.n71 4.5005
R864 VSS.n136 VSS.n71 4.5005
R865 VSS.n253 VSS.n71 4.5005
R866 VSS.n135 VSS.n71 4.5005
R867 VSS.n254 VSS.n71 4.5005
R868 VSS.n134 VSS.n71 4.5005
R869 VSS.n255 VSS.n71 4.5005
R870 VSS.n133 VSS.n71 4.5005
R871 VSS.n256 VSS.n71 4.5005
R872 VSS.n132 VSS.n71 4.5005
R873 VSS.n4502 VSS.n71 4.5005
R874 VSS.n4504 VSS.n71 4.5005
R875 VSS.n193 VSS.n65 4.5005
R876 VSS.n195 VSS.n65 4.5005
R877 VSS.n192 VSS.n65 4.5005
R878 VSS.n196 VSS.n65 4.5005
R879 VSS.n191 VSS.n65 4.5005
R880 VSS.n197 VSS.n65 4.5005
R881 VSS.n190 VSS.n65 4.5005
R882 VSS.n198 VSS.n65 4.5005
R883 VSS.n189 VSS.n65 4.5005
R884 VSS.n199 VSS.n65 4.5005
R885 VSS.n188 VSS.n65 4.5005
R886 VSS.n200 VSS.n65 4.5005
R887 VSS.n187 VSS.n65 4.5005
R888 VSS.n201 VSS.n65 4.5005
R889 VSS.n186 VSS.n65 4.5005
R890 VSS.n202 VSS.n65 4.5005
R891 VSS.n185 VSS.n65 4.5005
R892 VSS.n203 VSS.n65 4.5005
R893 VSS.n184 VSS.n65 4.5005
R894 VSS.n204 VSS.n65 4.5005
R895 VSS.n183 VSS.n65 4.5005
R896 VSS.n205 VSS.n65 4.5005
R897 VSS.n182 VSS.n65 4.5005
R898 VSS.n206 VSS.n65 4.5005
R899 VSS.n181 VSS.n65 4.5005
R900 VSS.n207 VSS.n65 4.5005
R901 VSS.n180 VSS.n65 4.5005
R902 VSS.n208 VSS.n65 4.5005
R903 VSS.n179 VSS.n65 4.5005
R904 VSS.n209 VSS.n65 4.5005
R905 VSS.n178 VSS.n65 4.5005
R906 VSS.n210 VSS.n65 4.5005
R907 VSS.n177 VSS.n65 4.5005
R908 VSS.n211 VSS.n65 4.5005
R909 VSS.n176 VSS.n65 4.5005
R910 VSS.n212 VSS.n65 4.5005
R911 VSS.n175 VSS.n65 4.5005
R912 VSS.n213 VSS.n65 4.5005
R913 VSS.n174 VSS.n65 4.5005
R914 VSS.n214 VSS.n65 4.5005
R915 VSS.n173 VSS.n65 4.5005
R916 VSS.n215 VSS.n65 4.5005
R917 VSS.n172 VSS.n65 4.5005
R918 VSS.n216 VSS.n65 4.5005
R919 VSS.n171 VSS.n65 4.5005
R920 VSS.n217 VSS.n65 4.5005
R921 VSS.n170 VSS.n65 4.5005
R922 VSS.n218 VSS.n65 4.5005
R923 VSS.n169 VSS.n65 4.5005
R924 VSS.n219 VSS.n65 4.5005
R925 VSS.n168 VSS.n65 4.5005
R926 VSS.n220 VSS.n65 4.5005
R927 VSS.n167 VSS.n65 4.5005
R928 VSS.n221 VSS.n65 4.5005
R929 VSS.n166 VSS.n65 4.5005
R930 VSS.n222 VSS.n65 4.5005
R931 VSS.n165 VSS.n65 4.5005
R932 VSS.n223 VSS.n65 4.5005
R933 VSS.n164 VSS.n65 4.5005
R934 VSS.n224 VSS.n65 4.5005
R935 VSS.n163 VSS.n65 4.5005
R936 VSS.n225 VSS.n65 4.5005
R937 VSS.n162 VSS.n65 4.5005
R938 VSS.n226 VSS.n65 4.5005
R939 VSS.n161 VSS.n65 4.5005
R940 VSS.n227 VSS.n65 4.5005
R941 VSS.n160 VSS.n65 4.5005
R942 VSS.n228 VSS.n65 4.5005
R943 VSS.n159 VSS.n65 4.5005
R944 VSS.n229 VSS.n65 4.5005
R945 VSS.n158 VSS.n65 4.5005
R946 VSS.n230 VSS.n65 4.5005
R947 VSS.n157 VSS.n65 4.5005
R948 VSS.n231 VSS.n65 4.5005
R949 VSS.n156 VSS.n65 4.5005
R950 VSS.n232 VSS.n65 4.5005
R951 VSS.n155 VSS.n65 4.5005
R952 VSS.n233 VSS.n65 4.5005
R953 VSS.n154 VSS.n65 4.5005
R954 VSS.n234 VSS.n65 4.5005
R955 VSS.n153 VSS.n65 4.5005
R956 VSS.n235 VSS.n65 4.5005
R957 VSS.n4506 VSS.n65 4.5005
R958 VSS.n236 VSS.n65 4.5005
R959 VSS.n152 VSS.n65 4.5005
R960 VSS.n237 VSS.n65 4.5005
R961 VSS.n151 VSS.n65 4.5005
R962 VSS.n238 VSS.n65 4.5005
R963 VSS.n150 VSS.n65 4.5005
R964 VSS.n239 VSS.n65 4.5005
R965 VSS.n149 VSS.n65 4.5005
R966 VSS.n240 VSS.n65 4.5005
R967 VSS.n148 VSS.n65 4.5005
R968 VSS.n241 VSS.n65 4.5005
R969 VSS.n147 VSS.n65 4.5005
R970 VSS.n242 VSS.n65 4.5005
R971 VSS.n146 VSS.n65 4.5005
R972 VSS.n243 VSS.n65 4.5005
R973 VSS.n145 VSS.n65 4.5005
R974 VSS.n244 VSS.n65 4.5005
R975 VSS.n144 VSS.n65 4.5005
R976 VSS.n245 VSS.n65 4.5005
R977 VSS.n143 VSS.n65 4.5005
R978 VSS.n246 VSS.n65 4.5005
R979 VSS.n142 VSS.n65 4.5005
R980 VSS.n247 VSS.n65 4.5005
R981 VSS.n141 VSS.n65 4.5005
R982 VSS.n248 VSS.n65 4.5005
R983 VSS.n140 VSS.n65 4.5005
R984 VSS.n249 VSS.n65 4.5005
R985 VSS.n139 VSS.n65 4.5005
R986 VSS.n250 VSS.n65 4.5005
R987 VSS.n138 VSS.n65 4.5005
R988 VSS.n251 VSS.n65 4.5005
R989 VSS.n137 VSS.n65 4.5005
R990 VSS.n252 VSS.n65 4.5005
R991 VSS.n136 VSS.n65 4.5005
R992 VSS.n253 VSS.n65 4.5005
R993 VSS.n135 VSS.n65 4.5005
R994 VSS.n254 VSS.n65 4.5005
R995 VSS.n134 VSS.n65 4.5005
R996 VSS.n255 VSS.n65 4.5005
R997 VSS.n133 VSS.n65 4.5005
R998 VSS.n256 VSS.n65 4.5005
R999 VSS.n132 VSS.n65 4.5005
R1000 VSS.n4502 VSS.n65 4.5005
R1001 VSS.n4504 VSS.n65 4.5005
R1002 VSS.n193 VSS.n72 4.5005
R1003 VSS.n195 VSS.n72 4.5005
R1004 VSS.n192 VSS.n72 4.5005
R1005 VSS.n196 VSS.n72 4.5005
R1006 VSS.n191 VSS.n72 4.5005
R1007 VSS.n197 VSS.n72 4.5005
R1008 VSS.n190 VSS.n72 4.5005
R1009 VSS.n198 VSS.n72 4.5005
R1010 VSS.n189 VSS.n72 4.5005
R1011 VSS.n199 VSS.n72 4.5005
R1012 VSS.n188 VSS.n72 4.5005
R1013 VSS.n200 VSS.n72 4.5005
R1014 VSS.n187 VSS.n72 4.5005
R1015 VSS.n201 VSS.n72 4.5005
R1016 VSS.n186 VSS.n72 4.5005
R1017 VSS.n202 VSS.n72 4.5005
R1018 VSS.n185 VSS.n72 4.5005
R1019 VSS.n203 VSS.n72 4.5005
R1020 VSS.n184 VSS.n72 4.5005
R1021 VSS.n204 VSS.n72 4.5005
R1022 VSS.n183 VSS.n72 4.5005
R1023 VSS.n205 VSS.n72 4.5005
R1024 VSS.n182 VSS.n72 4.5005
R1025 VSS.n206 VSS.n72 4.5005
R1026 VSS.n181 VSS.n72 4.5005
R1027 VSS.n207 VSS.n72 4.5005
R1028 VSS.n180 VSS.n72 4.5005
R1029 VSS.n208 VSS.n72 4.5005
R1030 VSS.n179 VSS.n72 4.5005
R1031 VSS.n209 VSS.n72 4.5005
R1032 VSS.n178 VSS.n72 4.5005
R1033 VSS.n210 VSS.n72 4.5005
R1034 VSS.n177 VSS.n72 4.5005
R1035 VSS.n211 VSS.n72 4.5005
R1036 VSS.n176 VSS.n72 4.5005
R1037 VSS.n212 VSS.n72 4.5005
R1038 VSS.n175 VSS.n72 4.5005
R1039 VSS.n213 VSS.n72 4.5005
R1040 VSS.n174 VSS.n72 4.5005
R1041 VSS.n214 VSS.n72 4.5005
R1042 VSS.n173 VSS.n72 4.5005
R1043 VSS.n215 VSS.n72 4.5005
R1044 VSS.n172 VSS.n72 4.5005
R1045 VSS.n216 VSS.n72 4.5005
R1046 VSS.n171 VSS.n72 4.5005
R1047 VSS.n217 VSS.n72 4.5005
R1048 VSS.n170 VSS.n72 4.5005
R1049 VSS.n218 VSS.n72 4.5005
R1050 VSS.n169 VSS.n72 4.5005
R1051 VSS.n219 VSS.n72 4.5005
R1052 VSS.n168 VSS.n72 4.5005
R1053 VSS.n220 VSS.n72 4.5005
R1054 VSS.n167 VSS.n72 4.5005
R1055 VSS.n221 VSS.n72 4.5005
R1056 VSS.n166 VSS.n72 4.5005
R1057 VSS.n222 VSS.n72 4.5005
R1058 VSS.n165 VSS.n72 4.5005
R1059 VSS.n223 VSS.n72 4.5005
R1060 VSS.n164 VSS.n72 4.5005
R1061 VSS.n224 VSS.n72 4.5005
R1062 VSS.n163 VSS.n72 4.5005
R1063 VSS.n225 VSS.n72 4.5005
R1064 VSS.n162 VSS.n72 4.5005
R1065 VSS.n226 VSS.n72 4.5005
R1066 VSS.n161 VSS.n72 4.5005
R1067 VSS.n227 VSS.n72 4.5005
R1068 VSS.n160 VSS.n72 4.5005
R1069 VSS.n228 VSS.n72 4.5005
R1070 VSS.n159 VSS.n72 4.5005
R1071 VSS.n229 VSS.n72 4.5005
R1072 VSS.n158 VSS.n72 4.5005
R1073 VSS.n230 VSS.n72 4.5005
R1074 VSS.n157 VSS.n72 4.5005
R1075 VSS.n231 VSS.n72 4.5005
R1076 VSS.n156 VSS.n72 4.5005
R1077 VSS.n232 VSS.n72 4.5005
R1078 VSS.n155 VSS.n72 4.5005
R1079 VSS.n233 VSS.n72 4.5005
R1080 VSS.n154 VSS.n72 4.5005
R1081 VSS.n234 VSS.n72 4.5005
R1082 VSS.n153 VSS.n72 4.5005
R1083 VSS.n235 VSS.n72 4.5005
R1084 VSS.n4506 VSS.n72 4.5005
R1085 VSS.n236 VSS.n72 4.5005
R1086 VSS.n152 VSS.n72 4.5005
R1087 VSS.n237 VSS.n72 4.5005
R1088 VSS.n151 VSS.n72 4.5005
R1089 VSS.n238 VSS.n72 4.5005
R1090 VSS.n150 VSS.n72 4.5005
R1091 VSS.n239 VSS.n72 4.5005
R1092 VSS.n149 VSS.n72 4.5005
R1093 VSS.n240 VSS.n72 4.5005
R1094 VSS.n148 VSS.n72 4.5005
R1095 VSS.n241 VSS.n72 4.5005
R1096 VSS.n147 VSS.n72 4.5005
R1097 VSS.n242 VSS.n72 4.5005
R1098 VSS.n146 VSS.n72 4.5005
R1099 VSS.n243 VSS.n72 4.5005
R1100 VSS.n145 VSS.n72 4.5005
R1101 VSS.n244 VSS.n72 4.5005
R1102 VSS.n144 VSS.n72 4.5005
R1103 VSS.n245 VSS.n72 4.5005
R1104 VSS.n143 VSS.n72 4.5005
R1105 VSS.n246 VSS.n72 4.5005
R1106 VSS.n142 VSS.n72 4.5005
R1107 VSS.n247 VSS.n72 4.5005
R1108 VSS.n141 VSS.n72 4.5005
R1109 VSS.n248 VSS.n72 4.5005
R1110 VSS.n140 VSS.n72 4.5005
R1111 VSS.n249 VSS.n72 4.5005
R1112 VSS.n139 VSS.n72 4.5005
R1113 VSS.n250 VSS.n72 4.5005
R1114 VSS.n138 VSS.n72 4.5005
R1115 VSS.n251 VSS.n72 4.5005
R1116 VSS.n137 VSS.n72 4.5005
R1117 VSS.n252 VSS.n72 4.5005
R1118 VSS.n136 VSS.n72 4.5005
R1119 VSS.n253 VSS.n72 4.5005
R1120 VSS.n135 VSS.n72 4.5005
R1121 VSS.n254 VSS.n72 4.5005
R1122 VSS.n134 VSS.n72 4.5005
R1123 VSS.n255 VSS.n72 4.5005
R1124 VSS.n133 VSS.n72 4.5005
R1125 VSS.n256 VSS.n72 4.5005
R1126 VSS.n132 VSS.n72 4.5005
R1127 VSS.n4502 VSS.n72 4.5005
R1128 VSS.n4504 VSS.n72 4.5005
R1129 VSS.n193 VSS.n64 4.5005
R1130 VSS.n195 VSS.n64 4.5005
R1131 VSS.n192 VSS.n64 4.5005
R1132 VSS.n196 VSS.n64 4.5005
R1133 VSS.n191 VSS.n64 4.5005
R1134 VSS.n197 VSS.n64 4.5005
R1135 VSS.n190 VSS.n64 4.5005
R1136 VSS.n198 VSS.n64 4.5005
R1137 VSS.n189 VSS.n64 4.5005
R1138 VSS.n199 VSS.n64 4.5005
R1139 VSS.n188 VSS.n64 4.5005
R1140 VSS.n200 VSS.n64 4.5005
R1141 VSS.n187 VSS.n64 4.5005
R1142 VSS.n201 VSS.n64 4.5005
R1143 VSS.n186 VSS.n64 4.5005
R1144 VSS.n202 VSS.n64 4.5005
R1145 VSS.n185 VSS.n64 4.5005
R1146 VSS.n203 VSS.n64 4.5005
R1147 VSS.n184 VSS.n64 4.5005
R1148 VSS.n204 VSS.n64 4.5005
R1149 VSS.n183 VSS.n64 4.5005
R1150 VSS.n205 VSS.n64 4.5005
R1151 VSS.n182 VSS.n64 4.5005
R1152 VSS.n206 VSS.n64 4.5005
R1153 VSS.n181 VSS.n64 4.5005
R1154 VSS.n207 VSS.n64 4.5005
R1155 VSS.n180 VSS.n64 4.5005
R1156 VSS.n208 VSS.n64 4.5005
R1157 VSS.n179 VSS.n64 4.5005
R1158 VSS.n209 VSS.n64 4.5005
R1159 VSS.n178 VSS.n64 4.5005
R1160 VSS.n210 VSS.n64 4.5005
R1161 VSS.n177 VSS.n64 4.5005
R1162 VSS.n211 VSS.n64 4.5005
R1163 VSS.n176 VSS.n64 4.5005
R1164 VSS.n212 VSS.n64 4.5005
R1165 VSS.n175 VSS.n64 4.5005
R1166 VSS.n213 VSS.n64 4.5005
R1167 VSS.n174 VSS.n64 4.5005
R1168 VSS.n214 VSS.n64 4.5005
R1169 VSS.n173 VSS.n64 4.5005
R1170 VSS.n215 VSS.n64 4.5005
R1171 VSS.n172 VSS.n64 4.5005
R1172 VSS.n216 VSS.n64 4.5005
R1173 VSS.n171 VSS.n64 4.5005
R1174 VSS.n217 VSS.n64 4.5005
R1175 VSS.n170 VSS.n64 4.5005
R1176 VSS.n218 VSS.n64 4.5005
R1177 VSS.n169 VSS.n64 4.5005
R1178 VSS.n219 VSS.n64 4.5005
R1179 VSS.n168 VSS.n64 4.5005
R1180 VSS.n220 VSS.n64 4.5005
R1181 VSS.n167 VSS.n64 4.5005
R1182 VSS.n221 VSS.n64 4.5005
R1183 VSS.n166 VSS.n64 4.5005
R1184 VSS.n222 VSS.n64 4.5005
R1185 VSS.n165 VSS.n64 4.5005
R1186 VSS.n223 VSS.n64 4.5005
R1187 VSS.n164 VSS.n64 4.5005
R1188 VSS.n224 VSS.n64 4.5005
R1189 VSS.n163 VSS.n64 4.5005
R1190 VSS.n225 VSS.n64 4.5005
R1191 VSS.n162 VSS.n64 4.5005
R1192 VSS.n226 VSS.n64 4.5005
R1193 VSS.n161 VSS.n64 4.5005
R1194 VSS.n227 VSS.n64 4.5005
R1195 VSS.n160 VSS.n64 4.5005
R1196 VSS.n228 VSS.n64 4.5005
R1197 VSS.n159 VSS.n64 4.5005
R1198 VSS.n229 VSS.n64 4.5005
R1199 VSS.n158 VSS.n64 4.5005
R1200 VSS.n230 VSS.n64 4.5005
R1201 VSS.n157 VSS.n64 4.5005
R1202 VSS.n231 VSS.n64 4.5005
R1203 VSS.n156 VSS.n64 4.5005
R1204 VSS.n232 VSS.n64 4.5005
R1205 VSS.n155 VSS.n64 4.5005
R1206 VSS.n233 VSS.n64 4.5005
R1207 VSS.n154 VSS.n64 4.5005
R1208 VSS.n234 VSS.n64 4.5005
R1209 VSS.n153 VSS.n64 4.5005
R1210 VSS.n235 VSS.n64 4.5005
R1211 VSS.n4506 VSS.n64 4.5005
R1212 VSS.n236 VSS.n64 4.5005
R1213 VSS.n152 VSS.n64 4.5005
R1214 VSS.n237 VSS.n64 4.5005
R1215 VSS.n151 VSS.n64 4.5005
R1216 VSS.n238 VSS.n64 4.5005
R1217 VSS.n150 VSS.n64 4.5005
R1218 VSS.n239 VSS.n64 4.5005
R1219 VSS.n149 VSS.n64 4.5005
R1220 VSS.n240 VSS.n64 4.5005
R1221 VSS.n148 VSS.n64 4.5005
R1222 VSS.n241 VSS.n64 4.5005
R1223 VSS.n147 VSS.n64 4.5005
R1224 VSS.n242 VSS.n64 4.5005
R1225 VSS.n146 VSS.n64 4.5005
R1226 VSS.n243 VSS.n64 4.5005
R1227 VSS.n145 VSS.n64 4.5005
R1228 VSS.n244 VSS.n64 4.5005
R1229 VSS.n144 VSS.n64 4.5005
R1230 VSS.n245 VSS.n64 4.5005
R1231 VSS.n143 VSS.n64 4.5005
R1232 VSS.n246 VSS.n64 4.5005
R1233 VSS.n142 VSS.n64 4.5005
R1234 VSS.n247 VSS.n64 4.5005
R1235 VSS.n141 VSS.n64 4.5005
R1236 VSS.n248 VSS.n64 4.5005
R1237 VSS.n140 VSS.n64 4.5005
R1238 VSS.n249 VSS.n64 4.5005
R1239 VSS.n139 VSS.n64 4.5005
R1240 VSS.n250 VSS.n64 4.5005
R1241 VSS.n138 VSS.n64 4.5005
R1242 VSS.n251 VSS.n64 4.5005
R1243 VSS.n137 VSS.n64 4.5005
R1244 VSS.n252 VSS.n64 4.5005
R1245 VSS.n136 VSS.n64 4.5005
R1246 VSS.n253 VSS.n64 4.5005
R1247 VSS.n135 VSS.n64 4.5005
R1248 VSS.n254 VSS.n64 4.5005
R1249 VSS.n134 VSS.n64 4.5005
R1250 VSS.n255 VSS.n64 4.5005
R1251 VSS.n133 VSS.n64 4.5005
R1252 VSS.n256 VSS.n64 4.5005
R1253 VSS.n132 VSS.n64 4.5005
R1254 VSS.n4502 VSS.n64 4.5005
R1255 VSS.n4504 VSS.n64 4.5005
R1256 VSS.n193 VSS.n73 4.5005
R1257 VSS.n195 VSS.n73 4.5005
R1258 VSS.n192 VSS.n73 4.5005
R1259 VSS.n196 VSS.n73 4.5005
R1260 VSS.n191 VSS.n73 4.5005
R1261 VSS.n197 VSS.n73 4.5005
R1262 VSS.n190 VSS.n73 4.5005
R1263 VSS.n198 VSS.n73 4.5005
R1264 VSS.n189 VSS.n73 4.5005
R1265 VSS.n199 VSS.n73 4.5005
R1266 VSS.n188 VSS.n73 4.5005
R1267 VSS.n200 VSS.n73 4.5005
R1268 VSS.n187 VSS.n73 4.5005
R1269 VSS.n201 VSS.n73 4.5005
R1270 VSS.n186 VSS.n73 4.5005
R1271 VSS.n202 VSS.n73 4.5005
R1272 VSS.n185 VSS.n73 4.5005
R1273 VSS.n203 VSS.n73 4.5005
R1274 VSS.n184 VSS.n73 4.5005
R1275 VSS.n204 VSS.n73 4.5005
R1276 VSS.n183 VSS.n73 4.5005
R1277 VSS.n205 VSS.n73 4.5005
R1278 VSS.n182 VSS.n73 4.5005
R1279 VSS.n206 VSS.n73 4.5005
R1280 VSS.n181 VSS.n73 4.5005
R1281 VSS.n207 VSS.n73 4.5005
R1282 VSS.n180 VSS.n73 4.5005
R1283 VSS.n208 VSS.n73 4.5005
R1284 VSS.n179 VSS.n73 4.5005
R1285 VSS.n209 VSS.n73 4.5005
R1286 VSS.n178 VSS.n73 4.5005
R1287 VSS.n210 VSS.n73 4.5005
R1288 VSS.n177 VSS.n73 4.5005
R1289 VSS.n211 VSS.n73 4.5005
R1290 VSS.n176 VSS.n73 4.5005
R1291 VSS.n212 VSS.n73 4.5005
R1292 VSS.n175 VSS.n73 4.5005
R1293 VSS.n213 VSS.n73 4.5005
R1294 VSS.n174 VSS.n73 4.5005
R1295 VSS.n214 VSS.n73 4.5005
R1296 VSS.n173 VSS.n73 4.5005
R1297 VSS.n215 VSS.n73 4.5005
R1298 VSS.n172 VSS.n73 4.5005
R1299 VSS.n216 VSS.n73 4.5005
R1300 VSS.n171 VSS.n73 4.5005
R1301 VSS.n217 VSS.n73 4.5005
R1302 VSS.n170 VSS.n73 4.5005
R1303 VSS.n218 VSS.n73 4.5005
R1304 VSS.n169 VSS.n73 4.5005
R1305 VSS.n219 VSS.n73 4.5005
R1306 VSS.n168 VSS.n73 4.5005
R1307 VSS.n220 VSS.n73 4.5005
R1308 VSS.n167 VSS.n73 4.5005
R1309 VSS.n221 VSS.n73 4.5005
R1310 VSS.n166 VSS.n73 4.5005
R1311 VSS.n222 VSS.n73 4.5005
R1312 VSS.n165 VSS.n73 4.5005
R1313 VSS.n223 VSS.n73 4.5005
R1314 VSS.n164 VSS.n73 4.5005
R1315 VSS.n224 VSS.n73 4.5005
R1316 VSS.n163 VSS.n73 4.5005
R1317 VSS.n225 VSS.n73 4.5005
R1318 VSS.n162 VSS.n73 4.5005
R1319 VSS.n226 VSS.n73 4.5005
R1320 VSS.n161 VSS.n73 4.5005
R1321 VSS.n227 VSS.n73 4.5005
R1322 VSS.n160 VSS.n73 4.5005
R1323 VSS.n228 VSS.n73 4.5005
R1324 VSS.n159 VSS.n73 4.5005
R1325 VSS.n229 VSS.n73 4.5005
R1326 VSS.n158 VSS.n73 4.5005
R1327 VSS.n230 VSS.n73 4.5005
R1328 VSS.n157 VSS.n73 4.5005
R1329 VSS.n231 VSS.n73 4.5005
R1330 VSS.n156 VSS.n73 4.5005
R1331 VSS.n232 VSS.n73 4.5005
R1332 VSS.n155 VSS.n73 4.5005
R1333 VSS.n233 VSS.n73 4.5005
R1334 VSS.n154 VSS.n73 4.5005
R1335 VSS.n234 VSS.n73 4.5005
R1336 VSS.n153 VSS.n73 4.5005
R1337 VSS.n235 VSS.n73 4.5005
R1338 VSS.n4506 VSS.n73 4.5005
R1339 VSS.n236 VSS.n73 4.5005
R1340 VSS.n152 VSS.n73 4.5005
R1341 VSS.n237 VSS.n73 4.5005
R1342 VSS.n151 VSS.n73 4.5005
R1343 VSS.n238 VSS.n73 4.5005
R1344 VSS.n150 VSS.n73 4.5005
R1345 VSS.n239 VSS.n73 4.5005
R1346 VSS.n149 VSS.n73 4.5005
R1347 VSS.n240 VSS.n73 4.5005
R1348 VSS.n148 VSS.n73 4.5005
R1349 VSS.n241 VSS.n73 4.5005
R1350 VSS.n147 VSS.n73 4.5005
R1351 VSS.n242 VSS.n73 4.5005
R1352 VSS.n146 VSS.n73 4.5005
R1353 VSS.n243 VSS.n73 4.5005
R1354 VSS.n145 VSS.n73 4.5005
R1355 VSS.n244 VSS.n73 4.5005
R1356 VSS.n144 VSS.n73 4.5005
R1357 VSS.n245 VSS.n73 4.5005
R1358 VSS.n143 VSS.n73 4.5005
R1359 VSS.n246 VSS.n73 4.5005
R1360 VSS.n142 VSS.n73 4.5005
R1361 VSS.n247 VSS.n73 4.5005
R1362 VSS.n141 VSS.n73 4.5005
R1363 VSS.n248 VSS.n73 4.5005
R1364 VSS.n140 VSS.n73 4.5005
R1365 VSS.n249 VSS.n73 4.5005
R1366 VSS.n139 VSS.n73 4.5005
R1367 VSS.n250 VSS.n73 4.5005
R1368 VSS.n138 VSS.n73 4.5005
R1369 VSS.n251 VSS.n73 4.5005
R1370 VSS.n137 VSS.n73 4.5005
R1371 VSS.n252 VSS.n73 4.5005
R1372 VSS.n136 VSS.n73 4.5005
R1373 VSS.n253 VSS.n73 4.5005
R1374 VSS.n135 VSS.n73 4.5005
R1375 VSS.n254 VSS.n73 4.5005
R1376 VSS.n134 VSS.n73 4.5005
R1377 VSS.n255 VSS.n73 4.5005
R1378 VSS.n133 VSS.n73 4.5005
R1379 VSS.n256 VSS.n73 4.5005
R1380 VSS.n132 VSS.n73 4.5005
R1381 VSS.n4502 VSS.n73 4.5005
R1382 VSS.n4504 VSS.n73 4.5005
R1383 VSS.n193 VSS.n63 4.5005
R1384 VSS.n195 VSS.n63 4.5005
R1385 VSS.n192 VSS.n63 4.5005
R1386 VSS.n196 VSS.n63 4.5005
R1387 VSS.n191 VSS.n63 4.5005
R1388 VSS.n197 VSS.n63 4.5005
R1389 VSS.n190 VSS.n63 4.5005
R1390 VSS.n198 VSS.n63 4.5005
R1391 VSS.n189 VSS.n63 4.5005
R1392 VSS.n199 VSS.n63 4.5005
R1393 VSS.n188 VSS.n63 4.5005
R1394 VSS.n200 VSS.n63 4.5005
R1395 VSS.n187 VSS.n63 4.5005
R1396 VSS.n201 VSS.n63 4.5005
R1397 VSS.n186 VSS.n63 4.5005
R1398 VSS.n202 VSS.n63 4.5005
R1399 VSS.n185 VSS.n63 4.5005
R1400 VSS.n203 VSS.n63 4.5005
R1401 VSS.n184 VSS.n63 4.5005
R1402 VSS.n204 VSS.n63 4.5005
R1403 VSS.n183 VSS.n63 4.5005
R1404 VSS.n205 VSS.n63 4.5005
R1405 VSS.n182 VSS.n63 4.5005
R1406 VSS.n206 VSS.n63 4.5005
R1407 VSS.n181 VSS.n63 4.5005
R1408 VSS.n207 VSS.n63 4.5005
R1409 VSS.n180 VSS.n63 4.5005
R1410 VSS.n208 VSS.n63 4.5005
R1411 VSS.n179 VSS.n63 4.5005
R1412 VSS.n209 VSS.n63 4.5005
R1413 VSS.n178 VSS.n63 4.5005
R1414 VSS.n210 VSS.n63 4.5005
R1415 VSS.n177 VSS.n63 4.5005
R1416 VSS.n211 VSS.n63 4.5005
R1417 VSS.n176 VSS.n63 4.5005
R1418 VSS.n212 VSS.n63 4.5005
R1419 VSS.n175 VSS.n63 4.5005
R1420 VSS.n213 VSS.n63 4.5005
R1421 VSS.n174 VSS.n63 4.5005
R1422 VSS.n214 VSS.n63 4.5005
R1423 VSS.n173 VSS.n63 4.5005
R1424 VSS.n215 VSS.n63 4.5005
R1425 VSS.n172 VSS.n63 4.5005
R1426 VSS.n216 VSS.n63 4.5005
R1427 VSS.n171 VSS.n63 4.5005
R1428 VSS.n217 VSS.n63 4.5005
R1429 VSS.n170 VSS.n63 4.5005
R1430 VSS.n218 VSS.n63 4.5005
R1431 VSS.n169 VSS.n63 4.5005
R1432 VSS.n219 VSS.n63 4.5005
R1433 VSS.n168 VSS.n63 4.5005
R1434 VSS.n220 VSS.n63 4.5005
R1435 VSS.n167 VSS.n63 4.5005
R1436 VSS.n221 VSS.n63 4.5005
R1437 VSS.n166 VSS.n63 4.5005
R1438 VSS.n222 VSS.n63 4.5005
R1439 VSS.n165 VSS.n63 4.5005
R1440 VSS.n223 VSS.n63 4.5005
R1441 VSS.n164 VSS.n63 4.5005
R1442 VSS.n224 VSS.n63 4.5005
R1443 VSS.n163 VSS.n63 4.5005
R1444 VSS.n225 VSS.n63 4.5005
R1445 VSS.n162 VSS.n63 4.5005
R1446 VSS.n226 VSS.n63 4.5005
R1447 VSS.n161 VSS.n63 4.5005
R1448 VSS.n227 VSS.n63 4.5005
R1449 VSS.n160 VSS.n63 4.5005
R1450 VSS.n228 VSS.n63 4.5005
R1451 VSS.n159 VSS.n63 4.5005
R1452 VSS.n229 VSS.n63 4.5005
R1453 VSS.n158 VSS.n63 4.5005
R1454 VSS.n230 VSS.n63 4.5005
R1455 VSS.n157 VSS.n63 4.5005
R1456 VSS.n231 VSS.n63 4.5005
R1457 VSS.n156 VSS.n63 4.5005
R1458 VSS.n232 VSS.n63 4.5005
R1459 VSS.n155 VSS.n63 4.5005
R1460 VSS.n233 VSS.n63 4.5005
R1461 VSS.n154 VSS.n63 4.5005
R1462 VSS.n234 VSS.n63 4.5005
R1463 VSS.n153 VSS.n63 4.5005
R1464 VSS.n235 VSS.n63 4.5005
R1465 VSS.n4506 VSS.n63 4.5005
R1466 VSS.n236 VSS.n63 4.5005
R1467 VSS.n152 VSS.n63 4.5005
R1468 VSS.n237 VSS.n63 4.5005
R1469 VSS.n151 VSS.n63 4.5005
R1470 VSS.n238 VSS.n63 4.5005
R1471 VSS.n150 VSS.n63 4.5005
R1472 VSS.n239 VSS.n63 4.5005
R1473 VSS.n149 VSS.n63 4.5005
R1474 VSS.n240 VSS.n63 4.5005
R1475 VSS.n148 VSS.n63 4.5005
R1476 VSS.n241 VSS.n63 4.5005
R1477 VSS.n147 VSS.n63 4.5005
R1478 VSS.n242 VSS.n63 4.5005
R1479 VSS.n146 VSS.n63 4.5005
R1480 VSS.n243 VSS.n63 4.5005
R1481 VSS.n145 VSS.n63 4.5005
R1482 VSS.n244 VSS.n63 4.5005
R1483 VSS.n144 VSS.n63 4.5005
R1484 VSS.n245 VSS.n63 4.5005
R1485 VSS.n143 VSS.n63 4.5005
R1486 VSS.n246 VSS.n63 4.5005
R1487 VSS.n142 VSS.n63 4.5005
R1488 VSS.n247 VSS.n63 4.5005
R1489 VSS.n141 VSS.n63 4.5005
R1490 VSS.n248 VSS.n63 4.5005
R1491 VSS.n140 VSS.n63 4.5005
R1492 VSS.n249 VSS.n63 4.5005
R1493 VSS.n139 VSS.n63 4.5005
R1494 VSS.n250 VSS.n63 4.5005
R1495 VSS.n138 VSS.n63 4.5005
R1496 VSS.n251 VSS.n63 4.5005
R1497 VSS.n137 VSS.n63 4.5005
R1498 VSS.n252 VSS.n63 4.5005
R1499 VSS.n136 VSS.n63 4.5005
R1500 VSS.n253 VSS.n63 4.5005
R1501 VSS.n135 VSS.n63 4.5005
R1502 VSS.n254 VSS.n63 4.5005
R1503 VSS.n134 VSS.n63 4.5005
R1504 VSS.n255 VSS.n63 4.5005
R1505 VSS.n133 VSS.n63 4.5005
R1506 VSS.n256 VSS.n63 4.5005
R1507 VSS.n132 VSS.n63 4.5005
R1508 VSS.n4502 VSS.n63 4.5005
R1509 VSS.n4504 VSS.n63 4.5005
R1510 VSS.n193 VSS.n74 4.5005
R1511 VSS.n195 VSS.n74 4.5005
R1512 VSS.n192 VSS.n74 4.5005
R1513 VSS.n196 VSS.n74 4.5005
R1514 VSS.n191 VSS.n74 4.5005
R1515 VSS.n197 VSS.n74 4.5005
R1516 VSS.n190 VSS.n74 4.5005
R1517 VSS.n198 VSS.n74 4.5005
R1518 VSS.n189 VSS.n74 4.5005
R1519 VSS.n199 VSS.n74 4.5005
R1520 VSS.n188 VSS.n74 4.5005
R1521 VSS.n200 VSS.n74 4.5005
R1522 VSS.n187 VSS.n74 4.5005
R1523 VSS.n201 VSS.n74 4.5005
R1524 VSS.n186 VSS.n74 4.5005
R1525 VSS.n202 VSS.n74 4.5005
R1526 VSS.n185 VSS.n74 4.5005
R1527 VSS.n203 VSS.n74 4.5005
R1528 VSS.n184 VSS.n74 4.5005
R1529 VSS.n204 VSS.n74 4.5005
R1530 VSS.n183 VSS.n74 4.5005
R1531 VSS.n205 VSS.n74 4.5005
R1532 VSS.n182 VSS.n74 4.5005
R1533 VSS.n206 VSS.n74 4.5005
R1534 VSS.n181 VSS.n74 4.5005
R1535 VSS.n207 VSS.n74 4.5005
R1536 VSS.n180 VSS.n74 4.5005
R1537 VSS.n208 VSS.n74 4.5005
R1538 VSS.n179 VSS.n74 4.5005
R1539 VSS.n209 VSS.n74 4.5005
R1540 VSS.n178 VSS.n74 4.5005
R1541 VSS.n210 VSS.n74 4.5005
R1542 VSS.n177 VSS.n74 4.5005
R1543 VSS.n211 VSS.n74 4.5005
R1544 VSS.n176 VSS.n74 4.5005
R1545 VSS.n212 VSS.n74 4.5005
R1546 VSS.n175 VSS.n74 4.5005
R1547 VSS.n213 VSS.n74 4.5005
R1548 VSS.n174 VSS.n74 4.5005
R1549 VSS.n214 VSS.n74 4.5005
R1550 VSS.n173 VSS.n74 4.5005
R1551 VSS.n215 VSS.n74 4.5005
R1552 VSS.n172 VSS.n74 4.5005
R1553 VSS.n216 VSS.n74 4.5005
R1554 VSS.n171 VSS.n74 4.5005
R1555 VSS.n217 VSS.n74 4.5005
R1556 VSS.n170 VSS.n74 4.5005
R1557 VSS.n218 VSS.n74 4.5005
R1558 VSS.n169 VSS.n74 4.5005
R1559 VSS.n219 VSS.n74 4.5005
R1560 VSS.n168 VSS.n74 4.5005
R1561 VSS.n220 VSS.n74 4.5005
R1562 VSS.n167 VSS.n74 4.5005
R1563 VSS.n221 VSS.n74 4.5005
R1564 VSS.n166 VSS.n74 4.5005
R1565 VSS.n222 VSS.n74 4.5005
R1566 VSS.n165 VSS.n74 4.5005
R1567 VSS.n223 VSS.n74 4.5005
R1568 VSS.n164 VSS.n74 4.5005
R1569 VSS.n224 VSS.n74 4.5005
R1570 VSS.n163 VSS.n74 4.5005
R1571 VSS.n225 VSS.n74 4.5005
R1572 VSS.n162 VSS.n74 4.5005
R1573 VSS.n226 VSS.n74 4.5005
R1574 VSS.n161 VSS.n74 4.5005
R1575 VSS.n227 VSS.n74 4.5005
R1576 VSS.n160 VSS.n74 4.5005
R1577 VSS.n228 VSS.n74 4.5005
R1578 VSS.n159 VSS.n74 4.5005
R1579 VSS.n229 VSS.n74 4.5005
R1580 VSS.n158 VSS.n74 4.5005
R1581 VSS.n230 VSS.n74 4.5005
R1582 VSS.n157 VSS.n74 4.5005
R1583 VSS.n231 VSS.n74 4.5005
R1584 VSS.n156 VSS.n74 4.5005
R1585 VSS.n232 VSS.n74 4.5005
R1586 VSS.n155 VSS.n74 4.5005
R1587 VSS.n233 VSS.n74 4.5005
R1588 VSS.n154 VSS.n74 4.5005
R1589 VSS.n234 VSS.n74 4.5005
R1590 VSS.n153 VSS.n74 4.5005
R1591 VSS.n235 VSS.n74 4.5005
R1592 VSS.n4506 VSS.n74 4.5005
R1593 VSS.n236 VSS.n74 4.5005
R1594 VSS.n152 VSS.n74 4.5005
R1595 VSS.n237 VSS.n74 4.5005
R1596 VSS.n151 VSS.n74 4.5005
R1597 VSS.n238 VSS.n74 4.5005
R1598 VSS.n150 VSS.n74 4.5005
R1599 VSS.n239 VSS.n74 4.5005
R1600 VSS.n149 VSS.n74 4.5005
R1601 VSS.n240 VSS.n74 4.5005
R1602 VSS.n148 VSS.n74 4.5005
R1603 VSS.n241 VSS.n74 4.5005
R1604 VSS.n147 VSS.n74 4.5005
R1605 VSS.n242 VSS.n74 4.5005
R1606 VSS.n146 VSS.n74 4.5005
R1607 VSS.n243 VSS.n74 4.5005
R1608 VSS.n145 VSS.n74 4.5005
R1609 VSS.n244 VSS.n74 4.5005
R1610 VSS.n144 VSS.n74 4.5005
R1611 VSS.n245 VSS.n74 4.5005
R1612 VSS.n143 VSS.n74 4.5005
R1613 VSS.n246 VSS.n74 4.5005
R1614 VSS.n142 VSS.n74 4.5005
R1615 VSS.n247 VSS.n74 4.5005
R1616 VSS.n141 VSS.n74 4.5005
R1617 VSS.n248 VSS.n74 4.5005
R1618 VSS.n140 VSS.n74 4.5005
R1619 VSS.n249 VSS.n74 4.5005
R1620 VSS.n139 VSS.n74 4.5005
R1621 VSS.n250 VSS.n74 4.5005
R1622 VSS.n138 VSS.n74 4.5005
R1623 VSS.n251 VSS.n74 4.5005
R1624 VSS.n137 VSS.n74 4.5005
R1625 VSS.n252 VSS.n74 4.5005
R1626 VSS.n136 VSS.n74 4.5005
R1627 VSS.n253 VSS.n74 4.5005
R1628 VSS.n135 VSS.n74 4.5005
R1629 VSS.n254 VSS.n74 4.5005
R1630 VSS.n134 VSS.n74 4.5005
R1631 VSS.n255 VSS.n74 4.5005
R1632 VSS.n133 VSS.n74 4.5005
R1633 VSS.n256 VSS.n74 4.5005
R1634 VSS.n132 VSS.n74 4.5005
R1635 VSS.n4502 VSS.n74 4.5005
R1636 VSS.n4504 VSS.n74 4.5005
R1637 VSS.n193 VSS.n62 4.5005
R1638 VSS.n195 VSS.n62 4.5005
R1639 VSS.n192 VSS.n62 4.5005
R1640 VSS.n196 VSS.n62 4.5005
R1641 VSS.n191 VSS.n62 4.5005
R1642 VSS.n197 VSS.n62 4.5005
R1643 VSS.n190 VSS.n62 4.5005
R1644 VSS.n198 VSS.n62 4.5005
R1645 VSS.n189 VSS.n62 4.5005
R1646 VSS.n199 VSS.n62 4.5005
R1647 VSS.n188 VSS.n62 4.5005
R1648 VSS.n200 VSS.n62 4.5005
R1649 VSS.n187 VSS.n62 4.5005
R1650 VSS.n201 VSS.n62 4.5005
R1651 VSS.n186 VSS.n62 4.5005
R1652 VSS.n202 VSS.n62 4.5005
R1653 VSS.n185 VSS.n62 4.5005
R1654 VSS.n203 VSS.n62 4.5005
R1655 VSS.n184 VSS.n62 4.5005
R1656 VSS.n204 VSS.n62 4.5005
R1657 VSS.n183 VSS.n62 4.5005
R1658 VSS.n205 VSS.n62 4.5005
R1659 VSS.n182 VSS.n62 4.5005
R1660 VSS.n206 VSS.n62 4.5005
R1661 VSS.n181 VSS.n62 4.5005
R1662 VSS.n207 VSS.n62 4.5005
R1663 VSS.n180 VSS.n62 4.5005
R1664 VSS.n208 VSS.n62 4.5005
R1665 VSS.n179 VSS.n62 4.5005
R1666 VSS.n209 VSS.n62 4.5005
R1667 VSS.n178 VSS.n62 4.5005
R1668 VSS.n210 VSS.n62 4.5005
R1669 VSS.n177 VSS.n62 4.5005
R1670 VSS.n211 VSS.n62 4.5005
R1671 VSS.n176 VSS.n62 4.5005
R1672 VSS.n212 VSS.n62 4.5005
R1673 VSS.n175 VSS.n62 4.5005
R1674 VSS.n213 VSS.n62 4.5005
R1675 VSS.n174 VSS.n62 4.5005
R1676 VSS.n214 VSS.n62 4.5005
R1677 VSS.n173 VSS.n62 4.5005
R1678 VSS.n215 VSS.n62 4.5005
R1679 VSS.n172 VSS.n62 4.5005
R1680 VSS.n216 VSS.n62 4.5005
R1681 VSS.n171 VSS.n62 4.5005
R1682 VSS.n217 VSS.n62 4.5005
R1683 VSS.n170 VSS.n62 4.5005
R1684 VSS.n218 VSS.n62 4.5005
R1685 VSS.n169 VSS.n62 4.5005
R1686 VSS.n219 VSS.n62 4.5005
R1687 VSS.n168 VSS.n62 4.5005
R1688 VSS.n220 VSS.n62 4.5005
R1689 VSS.n167 VSS.n62 4.5005
R1690 VSS.n221 VSS.n62 4.5005
R1691 VSS.n166 VSS.n62 4.5005
R1692 VSS.n222 VSS.n62 4.5005
R1693 VSS.n165 VSS.n62 4.5005
R1694 VSS.n223 VSS.n62 4.5005
R1695 VSS.n164 VSS.n62 4.5005
R1696 VSS.n224 VSS.n62 4.5005
R1697 VSS.n163 VSS.n62 4.5005
R1698 VSS.n225 VSS.n62 4.5005
R1699 VSS.n162 VSS.n62 4.5005
R1700 VSS.n226 VSS.n62 4.5005
R1701 VSS.n161 VSS.n62 4.5005
R1702 VSS.n227 VSS.n62 4.5005
R1703 VSS.n160 VSS.n62 4.5005
R1704 VSS.n228 VSS.n62 4.5005
R1705 VSS.n159 VSS.n62 4.5005
R1706 VSS.n229 VSS.n62 4.5005
R1707 VSS.n158 VSS.n62 4.5005
R1708 VSS.n230 VSS.n62 4.5005
R1709 VSS.n157 VSS.n62 4.5005
R1710 VSS.n231 VSS.n62 4.5005
R1711 VSS.n156 VSS.n62 4.5005
R1712 VSS.n232 VSS.n62 4.5005
R1713 VSS.n155 VSS.n62 4.5005
R1714 VSS.n233 VSS.n62 4.5005
R1715 VSS.n154 VSS.n62 4.5005
R1716 VSS.n234 VSS.n62 4.5005
R1717 VSS.n153 VSS.n62 4.5005
R1718 VSS.n235 VSS.n62 4.5005
R1719 VSS.n4506 VSS.n62 4.5005
R1720 VSS.n236 VSS.n62 4.5005
R1721 VSS.n152 VSS.n62 4.5005
R1722 VSS.n237 VSS.n62 4.5005
R1723 VSS.n151 VSS.n62 4.5005
R1724 VSS.n238 VSS.n62 4.5005
R1725 VSS.n150 VSS.n62 4.5005
R1726 VSS.n239 VSS.n62 4.5005
R1727 VSS.n149 VSS.n62 4.5005
R1728 VSS.n240 VSS.n62 4.5005
R1729 VSS.n148 VSS.n62 4.5005
R1730 VSS.n241 VSS.n62 4.5005
R1731 VSS.n147 VSS.n62 4.5005
R1732 VSS.n242 VSS.n62 4.5005
R1733 VSS.n146 VSS.n62 4.5005
R1734 VSS.n243 VSS.n62 4.5005
R1735 VSS.n145 VSS.n62 4.5005
R1736 VSS.n244 VSS.n62 4.5005
R1737 VSS.n144 VSS.n62 4.5005
R1738 VSS.n245 VSS.n62 4.5005
R1739 VSS.n143 VSS.n62 4.5005
R1740 VSS.n246 VSS.n62 4.5005
R1741 VSS.n142 VSS.n62 4.5005
R1742 VSS.n247 VSS.n62 4.5005
R1743 VSS.n141 VSS.n62 4.5005
R1744 VSS.n248 VSS.n62 4.5005
R1745 VSS.n140 VSS.n62 4.5005
R1746 VSS.n249 VSS.n62 4.5005
R1747 VSS.n139 VSS.n62 4.5005
R1748 VSS.n250 VSS.n62 4.5005
R1749 VSS.n138 VSS.n62 4.5005
R1750 VSS.n251 VSS.n62 4.5005
R1751 VSS.n137 VSS.n62 4.5005
R1752 VSS.n252 VSS.n62 4.5005
R1753 VSS.n136 VSS.n62 4.5005
R1754 VSS.n253 VSS.n62 4.5005
R1755 VSS.n135 VSS.n62 4.5005
R1756 VSS.n254 VSS.n62 4.5005
R1757 VSS.n134 VSS.n62 4.5005
R1758 VSS.n255 VSS.n62 4.5005
R1759 VSS.n133 VSS.n62 4.5005
R1760 VSS.n256 VSS.n62 4.5005
R1761 VSS.n132 VSS.n62 4.5005
R1762 VSS.n4502 VSS.n62 4.5005
R1763 VSS.n4504 VSS.n62 4.5005
R1764 VSS.n193 VSS.n75 4.5005
R1765 VSS.n195 VSS.n75 4.5005
R1766 VSS.n192 VSS.n75 4.5005
R1767 VSS.n196 VSS.n75 4.5005
R1768 VSS.n191 VSS.n75 4.5005
R1769 VSS.n197 VSS.n75 4.5005
R1770 VSS.n190 VSS.n75 4.5005
R1771 VSS.n198 VSS.n75 4.5005
R1772 VSS.n189 VSS.n75 4.5005
R1773 VSS.n199 VSS.n75 4.5005
R1774 VSS.n188 VSS.n75 4.5005
R1775 VSS.n200 VSS.n75 4.5005
R1776 VSS.n187 VSS.n75 4.5005
R1777 VSS.n201 VSS.n75 4.5005
R1778 VSS.n186 VSS.n75 4.5005
R1779 VSS.n202 VSS.n75 4.5005
R1780 VSS.n185 VSS.n75 4.5005
R1781 VSS.n203 VSS.n75 4.5005
R1782 VSS.n184 VSS.n75 4.5005
R1783 VSS.n204 VSS.n75 4.5005
R1784 VSS.n183 VSS.n75 4.5005
R1785 VSS.n205 VSS.n75 4.5005
R1786 VSS.n182 VSS.n75 4.5005
R1787 VSS.n206 VSS.n75 4.5005
R1788 VSS.n181 VSS.n75 4.5005
R1789 VSS.n207 VSS.n75 4.5005
R1790 VSS.n180 VSS.n75 4.5005
R1791 VSS.n208 VSS.n75 4.5005
R1792 VSS.n179 VSS.n75 4.5005
R1793 VSS.n209 VSS.n75 4.5005
R1794 VSS.n178 VSS.n75 4.5005
R1795 VSS.n210 VSS.n75 4.5005
R1796 VSS.n177 VSS.n75 4.5005
R1797 VSS.n211 VSS.n75 4.5005
R1798 VSS.n176 VSS.n75 4.5005
R1799 VSS.n212 VSS.n75 4.5005
R1800 VSS.n175 VSS.n75 4.5005
R1801 VSS.n213 VSS.n75 4.5005
R1802 VSS.n174 VSS.n75 4.5005
R1803 VSS.n214 VSS.n75 4.5005
R1804 VSS.n173 VSS.n75 4.5005
R1805 VSS.n215 VSS.n75 4.5005
R1806 VSS.n172 VSS.n75 4.5005
R1807 VSS.n216 VSS.n75 4.5005
R1808 VSS.n171 VSS.n75 4.5005
R1809 VSS.n217 VSS.n75 4.5005
R1810 VSS.n170 VSS.n75 4.5005
R1811 VSS.n218 VSS.n75 4.5005
R1812 VSS.n169 VSS.n75 4.5005
R1813 VSS.n219 VSS.n75 4.5005
R1814 VSS.n168 VSS.n75 4.5005
R1815 VSS.n220 VSS.n75 4.5005
R1816 VSS.n167 VSS.n75 4.5005
R1817 VSS.n221 VSS.n75 4.5005
R1818 VSS.n166 VSS.n75 4.5005
R1819 VSS.n222 VSS.n75 4.5005
R1820 VSS.n165 VSS.n75 4.5005
R1821 VSS.n223 VSS.n75 4.5005
R1822 VSS.n164 VSS.n75 4.5005
R1823 VSS.n224 VSS.n75 4.5005
R1824 VSS.n163 VSS.n75 4.5005
R1825 VSS.n225 VSS.n75 4.5005
R1826 VSS.n162 VSS.n75 4.5005
R1827 VSS.n226 VSS.n75 4.5005
R1828 VSS.n161 VSS.n75 4.5005
R1829 VSS.n227 VSS.n75 4.5005
R1830 VSS.n160 VSS.n75 4.5005
R1831 VSS.n228 VSS.n75 4.5005
R1832 VSS.n159 VSS.n75 4.5005
R1833 VSS.n229 VSS.n75 4.5005
R1834 VSS.n158 VSS.n75 4.5005
R1835 VSS.n230 VSS.n75 4.5005
R1836 VSS.n157 VSS.n75 4.5005
R1837 VSS.n231 VSS.n75 4.5005
R1838 VSS.n156 VSS.n75 4.5005
R1839 VSS.n232 VSS.n75 4.5005
R1840 VSS.n155 VSS.n75 4.5005
R1841 VSS.n233 VSS.n75 4.5005
R1842 VSS.n154 VSS.n75 4.5005
R1843 VSS.n234 VSS.n75 4.5005
R1844 VSS.n153 VSS.n75 4.5005
R1845 VSS.n235 VSS.n75 4.5005
R1846 VSS.n4506 VSS.n75 4.5005
R1847 VSS.n236 VSS.n75 4.5005
R1848 VSS.n152 VSS.n75 4.5005
R1849 VSS.n237 VSS.n75 4.5005
R1850 VSS.n151 VSS.n75 4.5005
R1851 VSS.n238 VSS.n75 4.5005
R1852 VSS.n150 VSS.n75 4.5005
R1853 VSS.n239 VSS.n75 4.5005
R1854 VSS.n149 VSS.n75 4.5005
R1855 VSS.n240 VSS.n75 4.5005
R1856 VSS.n148 VSS.n75 4.5005
R1857 VSS.n241 VSS.n75 4.5005
R1858 VSS.n147 VSS.n75 4.5005
R1859 VSS.n242 VSS.n75 4.5005
R1860 VSS.n146 VSS.n75 4.5005
R1861 VSS.n243 VSS.n75 4.5005
R1862 VSS.n145 VSS.n75 4.5005
R1863 VSS.n244 VSS.n75 4.5005
R1864 VSS.n144 VSS.n75 4.5005
R1865 VSS.n245 VSS.n75 4.5005
R1866 VSS.n143 VSS.n75 4.5005
R1867 VSS.n246 VSS.n75 4.5005
R1868 VSS.n142 VSS.n75 4.5005
R1869 VSS.n247 VSS.n75 4.5005
R1870 VSS.n141 VSS.n75 4.5005
R1871 VSS.n248 VSS.n75 4.5005
R1872 VSS.n140 VSS.n75 4.5005
R1873 VSS.n249 VSS.n75 4.5005
R1874 VSS.n139 VSS.n75 4.5005
R1875 VSS.n250 VSS.n75 4.5005
R1876 VSS.n138 VSS.n75 4.5005
R1877 VSS.n251 VSS.n75 4.5005
R1878 VSS.n137 VSS.n75 4.5005
R1879 VSS.n252 VSS.n75 4.5005
R1880 VSS.n136 VSS.n75 4.5005
R1881 VSS.n253 VSS.n75 4.5005
R1882 VSS.n135 VSS.n75 4.5005
R1883 VSS.n254 VSS.n75 4.5005
R1884 VSS.n134 VSS.n75 4.5005
R1885 VSS.n255 VSS.n75 4.5005
R1886 VSS.n133 VSS.n75 4.5005
R1887 VSS.n256 VSS.n75 4.5005
R1888 VSS.n132 VSS.n75 4.5005
R1889 VSS.n4502 VSS.n75 4.5005
R1890 VSS.n4504 VSS.n75 4.5005
R1891 VSS.n193 VSS.n61 4.5005
R1892 VSS.n195 VSS.n61 4.5005
R1893 VSS.n192 VSS.n61 4.5005
R1894 VSS.n196 VSS.n61 4.5005
R1895 VSS.n191 VSS.n61 4.5005
R1896 VSS.n197 VSS.n61 4.5005
R1897 VSS.n190 VSS.n61 4.5005
R1898 VSS.n198 VSS.n61 4.5005
R1899 VSS.n189 VSS.n61 4.5005
R1900 VSS.n199 VSS.n61 4.5005
R1901 VSS.n188 VSS.n61 4.5005
R1902 VSS.n200 VSS.n61 4.5005
R1903 VSS.n187 VSS.n61 4.5005
R1904 VSS.n201 VSS.n61 4.5005
R1905 VSS.n186 VSS.n61 4.5005
R1906 VSS.n202 VSS.n61 4.5005
R1907 VSS.n185 VSS.n61 4.5005
R1908 VSS.n203 VSS.n61 4.5005
R1909 VSS.n184 VSS.n61 4.5005
R1910 VSS.n204 VSS.n61 4.5005
R1911 VSS.n183 VSS.n61 4.5005
R1912 VSS.n205 VSS.n61 4.5005
R1913 VSS.n182 VSS.n61 4.5005
R1914 VSS.n206 VSS.n61 4.5005
R1915 VSS.n181 VSS.n61 4.5005
R1916 VSS.n207 VSS.n61 4.5005
R1917 VSS.n180 VSS.n61 4.5005
R1918 VSS.n208 VSS.n61 4.5005
R1919 VSS.n179 VSS.n61 4.5005
R1920 VSS.n209 VSS.n61 4.5005
R1921 VSS.n178 VSS.n61 4.5005
R1922 VSS.n210 VSS.n61 4.5005
R1923 VSS.n177 VSS.n61 4.5005
R1924 VSS.n211 VSS.n61 4.5005
R1925 VSS.n176 VSS.n61 4.5005
R1926 VSS.n212 VSS.n61 4.5005
R1927 VSS.n175 VSS.n61 4.5005
R1928 VSS.n213 VSS.n61 4.5005
R1929 VSS.n174 VSS.n61 4.5005
R1930 VSS.n214 VSS.n61 4.5005
R1931 VSS.n173 VSS.n61 4.5005
R1932 VSS.n215 VSS.n61 4.5005
R1933 VSS.n172 VSS.n61 4.5005
R1934 VSS.n216 VSS.n61 4.5005
R1935 VSS.n171 VSS.n61 4.5005
R1936 VSS.n217 VSS.n61 4.5005
R1937 VSS.n170 VSS.n61 4.5005
R1938 VSS.n218 VSS.n61 4.5005
R1939 VSS.n169 VSS.n61 4.5005
R1940 VSS.n219 VSS.n61 4.5005
R1941 VSS.n168 VSS.n61 4.5005
R1942 VSS.n220 VSS.n61 4.5005
R1943 VSS.n167 VSS.n61 4.5005
R1944 VSS.n221 VSS.n61 4.5005
R1945 VSS.n166 VSS.n61 4.5005
R1946 VSS.n222 VSS.n61 4.5005
R1947 VSS.n165 VSS.n61 4.5005
R1948 VSS.n223 VSS.n61 4.5005
R1949 VSS.n164 VSS.n61 4.5005
R1950 VSS.n224 VSS.n61 4.5005
R1951 VSS.n163 VSS.n61 4.5005
R1952 VSS.n225 VSS.n61 4.5005
R1953 VSS.n162 VSS.n61 4.5005
R1954 VSS.n226 VSS.n61 4.5005
R1955 VSS.n161 VSS.n61 4.5005
R1956 VSS.n227 VSS.n61 4.5005
R1957 VSS.n160 VSS.n61 4.5005
R1958 VSS.n228 VSS.n61 4.5005
R1959 VSS.n159 VSS.n61 4.5005
R1960 VSS.n229 VSS.n61 4.5005
R1961 VSS.n158 VSS.n61 4.5005
R1962 VSS.n230 VSS.n61 4.5005
R1963 VSS.n157 VSS.n61 4.5005
R1964 VSS.n231 VSS.n61 4.5005
R1965 VSS.n156 VSS.n61 4.5005
R1966 VSS.n232 VSS.n61 4.5005
R1967 VSS.n155 VSS.n61 4.5005
R1968 VSS.n233 VSS.n61 4.5005
R1969 VSS.n154 VSS.n61 4.5005
R1970 VSS.n234 VSS.n61 4.5005
R1971 VSS.n153 VSS.n61 4.5005
R1972 VSS.n235 VSS.n61 4.5005
R1973 VSS.n4506 VSS.n61 4.5005
R1974 VSS.n236 VSS.n61 4.5005
R1975 VSS.n152 VSS.n61 4.5005
R1976 VSS.n237 VSS.n61 4.5005
R1977 VSS.n151 VSS.n61 4.5005
R1978 VSS.n238 VSS.n61 4.5005
R1979 VSS.n150 VSS.n61 4.5005
R1980 VSS.n239 VSS.n61 4.5005
R1981 VSS.n149 VSS.n61 4.5005
R1982 VSS.n240 VSS.n61 4.5005
R1983 VSS.n148 VSS.n61 4.5005
R1984 VSS.n241 VSS.n61 4.5005
R1985 VSS.n147 VSS.n61 4.5005
R1986 VSS.n242 VSS.n61 4.5005
R1987 VSS.n146 VSS.n61 4.5005
R1988 VSS.n243 VSS.n61 4.5005
R1989 VSS.n145 VSS.n61 4.5005
R1990 VSS.n244 VSS.n61 4.5005
R1991 VSS.n144 VSS.n61 4.5005
R1992 VSS.n245 VSS.n61 4.5005
R1993 VSS.n143 VSS.n61 4.5005
R1994 VSS.n246 VSS.n61 4.5005
R1995 VSS.n142 VSS.n61 4.5005
R1996 VSS.n247 VSS.n61 4.5005
R1997 VSS.n141 VSS.n61 4.5005
R1998 VSS.n248 VSS.n61 4.5005
R1999 VSS.n140 VSS.n61 4.5005
R2000 VSS.n249 VSS.n61 4.5005
R2001 VSS.n139 VSS.n61 4.5005
R2002 VSS.n250 VSS.n61 4.5005
R2003 VSS.n138 VSS.n61 4.5005
R2004 VSS.n251 VSS.n61 4.5005
R2005 VSS.n137 VSS.n61 4.5005
R2006 VSS.n252 VSS.n61 4.5005
R2007 VSS.n136 VSS.n61 4.5005
R2008 VSS.n253 VSS.n61 4.5005
R2009 VSS.n135 VSS.n61 4.5005
R2010 VSS.n254 VSS.n61 4.5005
R2011 VSS.n134 VSS.n61 4.5005
R2012 VSS.n255 VSS.n61 4.5005
R2013 VSS.n133 VSS.n61 4.5005
R2014 VSS.n256 VSS.n61 4.5005
R2015 VSS.n132 VSS.n61 4.5005
R2016 VSS.n4502 VSS.n61 4.5005
R2017 VSS.n4504 VSS.n61 4.5005
R2018 VSS.n193 VSS.n76 4.5005
R2019 VSS.n195 VSS.n76 4.5005
R2020 VSS.n192 VSS.n76 4.5005
R2021 VSS.n196 VSS.n76 4.5005
R2022 VSS.n191 VSS.n76 4.5005
R2023 VSS.n197 VSS.n76 4.5005
R2024 VSS.n190 VSS.n76 4.5005
R2025 VSS.n198 VSS.n76 4.5005
R2026 VSS.n189 VSS.n76 4.5005
R2027 VSS.n199 VSS.n76 4.5005
R2028 VSS.n188 VSS.n76 4.5005
R2029 VSS.n200 VSS.n76 4.5005
R2030 VSS.n187 VSS.n76 4.5005
R2031 VSS.n201 VSS.n76 4.5005
R2032 VSS.n186 VSS.n76 4.5005
R2033 VSS.n202 VSS.n76 4.5005
R2034 VSS.n185 VSS.n76 4.5005
R2035 VSS.n203 VSS.n76 4.5005
R2036 VSS.n184 VSS.n76 4.5005
R2037 VSS.n204 VSS.n76 4.5005
R2038 VSS.n183 VSS.n76 4.5005
R2039 VSS.n205 VSS.n76 4.5005
R2040 VSS.n182 VSS.n76 4.5005
R2041 VSS.n206 VSS.n76 4.5005
R2042 VSS.n181 VSS.n76 4.5005
R2043 VSS.n207 VSS.n76 4.5005
R2044 VSS.n180 VSS.n76 4.5005
R2045 VSS.n208 VSS.n76 4.5005
R2046 VSS.n179 VSS.n76 4.5005
R2047 VSS.n209 VSS.n76 4.5005
R2048 VSS.n178 VSS.n76 4.5005
R2049 VSS.n210 VSS.n76 4.5005
R2050 VSS.n177 VSS.n76 4.5005
R2051 VSS.n211 VSS.n76 4.5005
R2052 VSS.n176 VSS.n76 4.5005
R2053 VSS.n212 VSS.n76 4.5005
R2054 VSS.n175 VSS.n76 4.5005
R2055 VSS.n213 VSS.n76 4.5005
R2056 VSS.n174 VSS.n76 4.5005
R2057 VSS.n214 VSS.n76 4.5005
R2058 VSS.n173 VSS.n76 4.5005
R2059 VSS.n215 VSS.n76 4.5005
R2060 VSS.n172 VSS.n76 4.5005
R2061 VSS.n216 VSS.n76 4.5005
R2062 VSS.n171 VSS.n76 4.5005
R2063 VSS.n217 VSS.n76 4.5005
R2064 VSS.n170 VSS.n76 4.5005
R2065 VSS.n218 VSS.n76 4.5005
R2066 VSS.n169 VSS.n76 4.5005
R2067 VSS.n219 VSS.n76 4.5005
R2068 VSS.n168 VSS.n76 4.5005
R2069 VSS.n220 VSS.n76 4.5005
R2070 VSS.n167 VSS.n76 4.5005
R2071 VSS.n221 VSS.n76 4.5005
R2072 VSS.n166 VSS.n76 4.5005
R2073 VSS.n222 VSS.n76 4.5005
R2074 VSS.n165 VSS.n76 4.5005
R2075 VSS.n223 VSS.n76 4.5005
R2076 VSS.n164 VSS.n76 4.5005
R2077 VSS.n224 VSS.n76 4.5005
R2078 VSS.n163 VSS.n76 4.5005
R2079 VSS.n225 VSS.n76 4.5005
R2080 VSS.n162 VSS.n76 4.5005
R2081 VSS.n226 VSS.n76 4.5005
R2082 VSS.n161 VSS.n76 4.5005
R2083 VSS.n227 VSS.n76 4.5005
R2084 VSS.n160 VSS.n76 4.5005
R2085 VSS.n228 VSS.n76 4.5005
R2086 VSS.n159 VSS.n76 4.5005
R2087 VSS.n229 VSS.n76 4.5005
R2088 VSS.n158 VSS.n76 4.5005
R2089 VSS.n230 VSS.n76 4.5005
R2090 VSS.n157 VSS.n76 4.5005
R2091 VSS.n231 VSS.n76 4.5005
R2092 VSS.n156 VSS.n76 4.5005
R2093 VSS.n232 VSS.n76 4.5005
R2094 VSS.n155 VSS.n76 4.5005
R2095 VSS.n233 VSS.n76 4.5005
R2096 VSS.n154 VSS.n76 4.5005
R2097 VSS.n234 VSS.n76 4.5005
R2098 VSS.n153 VSS.n76 4.5005
R2099 VSS.n235 VSS.n76 4.5005
R2100 VSS.n4506 VSS.n76 4.5005
R2101 VSS.n236 VSS.n76 4.5005
R2102 VSS.n152 VSS.n76 4.5005
R2103 VSS.n237 VSS.n76 4.5005
R2104 VSS.n151 VSS.n76 4.5005
R2105 VSS.n238 VSS.n76 4.5005
R2106 VSS.n150 VSS.n76 4.5005
R2107 VSS.n239 VSS.n76 4.5005
R2108 VSS.n149 VSS.n76 4.5005
R2109 VSS.n240 VSS.n76 4.5005
R2110 VSS.n148 VSS.n76 4.5005
R2111 VSS.n241 VSS.n76 4.5005
R2112 VSS.n147 VSS.n76 4.5005
R2113 VSS.n242 VSS.n76 4.5005
R2114 VSS.n146 VSS.n76 4.5005
R2115 VSS.n243 VSS.n76 4.5005
R2116 VSS.n145 VSS.n76 4.5005
R2117 VSS.n244 VSS.n76 4.5005
R2118 VSS.n144 VSS.n76 4.5005
R2119 VSS.n245 VSS.n76 4.5005
R2120 VSS.n143 VSS.n76 4.5005
R2121 VSS.n246 VSS.n76 4.5005
R2122 VSS.n142 VSS.n76 4.5005
R2123 VSS.n247 VSS.n76 4.5005
R2124 VSS.n141 VSS.n76 4.5005
R2125 VSS.n248 VSS.n76 4.5005
R2126 VSS.n140 VSS.n76 4.5005
R2127 VSS.n249 VSS.n76 4.5005
R2128 VSS.n139 VSS.n76 4.5005
R2129 VSS.n250 VSS.n76 4.5005
R2130 VSS.n138 VSS.n76 4.5005
R2131 VSS.n251 VSS.n76 4.5005
R2132 VSS.n137 VSS.n76 4.5005
R2133 VSS.n252 VSS.n76 4.5005
R2134 VSS.n136 VSS.n76 4.5005
R2135 VSS.n253 VSS.n76 4.5005
R2136 VSS.n135 VSS.n76 4.5005
R2137 VSS.n254 VSS.n76 4.5005
R2138 VSS.n134 VSS.n76 4.5005
R2139 VSS.n255 VSS.n76 4.5005
R2140 VSS.n133 VSS.n76 4.5005
R2141 VSS.n256 VSS.n76 4.5005
R2142 VSS.n132 VSS.n76 4.5005
R2143 VSS.n4502 VSS.n76 4.5005
R2144 VSS.n4504 VSS.n76 4.5005
R2145 VSS.n193 VSS.n60 4.5005
R2146 VSS.n195 VSS.n60 4.5005
R2147 VSS.n192 VSS.n60 4.5005
R2148 VSS.n196 VSS.n60 4.5005
R2149 VSS.n191 VSS.n60 4.5005
R2150 VSS.n197 VSS.n60 4.5005
R2151 VSS.n190 VSS.n60 4.5005
R2152 VSS.n198 VSS.n60 4.5005
R2153 VSS.n189 VSS.n60 4.5005
R2154 VSS.n199 VSS.n60 4.5005
R2155 VSS.n188 VSS.n60 4.5005
R2156 VSS.n200 VSS.n60 4.5005
R2157 VSS.n187 VSS.n60 4.5005
R2158 VSS.n201 VSS.n60 4.5005
R2159 VSS.n186 VSS.n60 4.5005
R2160 VSS.n202 VSS.n60 4.5005
R2161 VSS.n185 VSS.n60 4.5005
R2162 VSS.n203 VSS.n60 4.5005
R2163 VSS.n184 VSS.n60 4.5005
R2164 VSS.n204 VSS.n60 4.5005
R2165 VSS.n183 VSS.n60 4.5005
R2166 VSS.n205 VSS.n60 4.5005
R2167 VSS.n182 VSS.n60 4.5005
R2168 VSS.n206 VSS.n60 4.5005
R2169 VSS.n181 VSS.n60 4.5005
R2170 VSS.n207 VSS.n60 4.5005
R2171 VSS.n180 VSS.n60 4.5005
R2172 VSS.n208 VSS.n60 4.5005
R2173 VSS.n179 VSS.n60 4.5005
R2174 VSS.n209 VSS.n60 4.5005
R2175 VSS.n178 VSS.n60 4.5005
R2176 VSS.n210 VSS.n60 4.5005
R2177 VSS.n177 VSS.n60 4.5005
R2178 VSS.n211 VSS.n60 4.5005
R2179 VSS.n176 VSS.n60 4.5005
R2180 VSS.n212 VSS.n60 4.5005
R2181 VSS.n175 VSS.n60 4.5005
R2182 VSS.n213 VSS.n60 4.5005
R2183 VSS.n174 VSS.n60 4.5005
R2184 VSS.n214 VSS.n60 4.5005
R2185 VSS.n173 VSS.n60 4.5005
R2186 VSS.n215 VSS.n60 4.5005
R2187 VSS.n172 VSS.n60 4.5005
R2188 VSS.n216 VSS.n60 4.5005
R2189 VSS.n171 VSS.n60 4.5005
R2190 VSS.n217 VSS.n60 4.5005
R2191 VSS.n170 VSS.n60 4.5005
R2192 VSS.n218 VSS.n60 4.5005
R2193 VSS.n169 VSS.n60 4.5005
R2194 VSS.n219 VSS.n60 4.5005
R2195 VSS.n168 VSS.n60 4.5005
R2196 VSS.n220 VSS.n60 4.5005
R2197 VSS.n167 VSS.n60 4.5005
R2198 VSS.n221 VSS.n60 4.5005
R2199 VSS.n166 VSS.n60 4.5005
R2200 VSS.n222 VSS.n60 4.5005
R2201 VSS.n165 VSS.n60 4.5005
R2202 VSS.n223 VSS.n60 4.5005
R2203 VSS.n164 VSS.n60 4.5005
R2204 VSS.n224 VSS.n60 4.5005
R2205 VSS.n163 VSS.n60 4.5005
R2206 VSS.n225 VSS.n60 4.5005
R2207 VSS.n162 VSS.n60 4.5005
R2208 VSS.n226 VSS.n60 4.5005
R2209 VSS.n161 VSS.n60 4.5005
R2210 VSS.n227 VSS.n60 4.5005
R2211 VSS.n160 VSS.n60 4.5005
R2212 VSS.n228 VSS.n60 4.5005
R2213 VSS.n159 VSS.n60 4.5005
R2214 VSS.n229 VSS.n60 4.5005
R2215 VSS.n158 VSS.n60 4.5005
R2216 VSS.n230 VSS.n60 4.5005
R2217 VSS.n157 VSS.n60 4.5005
R2218 VSS.n231 VSS.n60 4.5005
R2219 VSS.n156 VSS.n60 4.5005
R2220 VSS.n232 VSS.n60 4.5005
R2221 VSS.n155 VSS.n60 4.5005
R2222 VSS.n233 VSS.n60 4.5005
R2223 VSS.n154 VSS.n60 4.5005
R2224 VSS.n234 VSS.n60 4.5005
R2225 VSS.n153 VSS.n60 4.5005
R2226 VSS.n235 VSS.n60 4.5005
R2227 VSS.n4506 VSS.n60 4.5005
R2228 VSS.n236 VSS.n60 4.5005
R2229 VSS.n152 VSS.n60 4.5005
R2230 VSS.n237 VSS.n60 4.5005
R2231 VSS.n151 VSS.n60 4.5005
R2232 VSS.n238 VSS.n60 4.5005
R2233 VSS.n150 VSS.n60 4.5005
R2234 VSS.n239 VSS.n60 4.5005
R2235 VSS.n149 VSS.n60 4.5005
R2236 VSS.n240 VSS.n60 4.5005
R2237 VSS.n148 VSS.n60 4.5005
R2238 VSS.n241 VSS.n60 4.5005
R2239 VSS.n147 VSS.n60 4.5005
R2240 VSS.n242 VSS.n60 4.5005
R2241 VSS.n146 VSS.n60 4.5005
R2242 VSS.n243 VSS.n60 4.5005
R2243 VSS.n145 VSS.n60 4.5005
R2244 VSS.n244 VSS.n60 4.5005
R2245 VSS.n144 VSS.n60 4.5005
R2246 VSS.n245 VSS.n60 4.5005
R2247 VSS.n143 VSS.n60 4.5005
R2248 VSS.n246 VSS.n60 4.5005
R2249 VSS.n142 VSS.n60 4.5005
R2250 VSS.n247 VSS.n60 4.5005
R2251 VSS.n141 VSS.n60 4.5005
R2252 VSS.n248 VSS.n60 4.5005
R2253 VSS.n140 VSS.n60 4.5005
R2254 VSS.n249 VSS.n60 4.5005
R2255 VSS.n139 VSS.n60 4.5005
R2256 VSS.n250 VSS.n60 4.5005
R2257 VSS.n138 VSS.n60 4.5005
R2258 VSS.n251 VSS.n60 4.5005
R2259 VSS.n137 VSS.n60 4.5005
R2260 VSS.n252 VSS.n60 4.5005
R2261 VSS.n136 VSS.n60 4.5005
R2262 VSS.n253 VSS.n60 4.5005
R2263 VSS.n135 VSS.n60 4.5005
R2264 VSS.n254 VSS.n60 4.5005
R2265 VSS.n134 VSS.n60 4.5005
R2266 VSS.n255 VSS.n60 4.5005
R2267 VSS.n133 VSS.n60 4.5005
R2268 VSS.n256 VSS.n60 4.5005
R2269 VSS.n132 VSS.n60 4.5005
R2270 VSS.n4502 VSS.n60 4.5005
R2271 VSS.n4504 VSS.n60 4.5005
R2272 VSS.n193 VSS.n77 4.5005
R2273 VSS.n195 VSS.n77 4.5005
R2274 VSS.n192 VSS.n77 4.5005
R2275 VSS.n196 VSS.n77 4.5005
R2276 VSS.n191 VSS.n77 4.5005
R2277 VSS.n197 VSS.n77 4.5005
R2278 VSS.n190 VSS.n77 4.5005
R2279 VSS.n198 VSS.n77 4.5005
R2280 VSS.n189 VSS.n77 4.5005
R2281 VSS.n199 VSS.n77 4.5005
R2282 VSS.n188 VSS.n77 4.5005
R2283 VSS.n200 VSS.n77 4.5005
R2284 VSS.n187 VSS.n77 4.5005
R2285 VSS.n201 VSS.n77 4.5005
R2286 VSS.n186 VSS.n77 4.5005
R2287 VSS.n202 VSS.n77 4.5005
R2288 VSS.n185 VSS.n77 4.5005
R2289 VSS.n203 VSS.n77 4.5005
R2290 VSS.n184 VSS.n77 4.5005
R2291 VSS.n204 VSS.n77 4.5005
R2292 VSS.n183 VSS.n77 4.5005
R2293 VSS.n205 VSS.n77 4.5005
R2294 VSS.n182 VSS.n77 4.5005
R2295 VSS.n206 VSS.n77 4.5005
R2296 VSS.n181 VSS.n77 4.5005
R2297 VSS.n207 VSS.n77 4.5005
R2298 VSS.n180 VSS.n77 4.5005
R2299 VSS.n208 VSS.n77 4.5005
R2300 VSS.n179 VSS.n77 4.5005
R2301 VSS.n209 VSS.n77 4.5005
R2302 VSS.n178 VSS.n77 4.5005
R2303 VSS.n210 VSS.n77 4.5005
R2304 VSS.n177 VSS.n77 4.5005
R2305 VSS.n211 VSS.n77 4.5005
R2306 VSS.n176 VSS.n77 4.5005
R2307 VSS.n212 VSS.n77 4.5005
R2308 VSS.n175 VSS.n77 4.5005
R2309 VSS.n213 VSS.n77 4.5005
R2310 VSS.n174 VSS.n77 4.5005
R2311 VSS.n214 VSS.n77 4.5005
R2312 VSS.n173 VSS.n77 4.5005
R2313 VSS.n215 VSS.n77 4.5005
R2314 VSS.n172 VSS.n77 4.5005
R2315 VSS.n216 VSS.n77 4.5005
R2316 VSS.n171 VSS.n77 4.5005
R2317 VSS.n217 VSS.n77 4.5005
R2318 VSS.n170 VSS.n77 4.5005
R2319 VSS.n218 VSS.n77 4.5005
R2320 VSS.n169 VSS.n77 4.5005
R2321 VSS.n219 VSS.n77 4.5005
R2322 VSS.n168 VSS.n77 4.5005
R2323 VSS.n220 VSS.n77 4.5005
R2324 VSS.n167 VSS.n77 4.5005
R2325 VSS.n221 VSS.n77 4.5005
R2326 VSS.n166 VSS.n77 4.5005
R2327 VSS.n222 VSS.n77 4.5005
R2328 VSS.n165 VSS.n77 4.5005
R2329 VSS.n223 VSS.n77 4.5005
R2330 VSS.n164 VSS.n77 4.5005
R2331 VSS.n224 VSS.n77 4.5005
R2332 VSS.n163 VSS.n77 4.5005
R2333 VSS.n225 VSS.n77 4.5005
R2334 VSS.n162 VSS.n77 4.5005
R2335 VSS.n226 VSS.n77 4.5005
R2336 VSS.n161 VSS.n77 4.5005
R2337 VSS.n227 VSS.n77 4.5005
R2338 VSS.n160 VSS.n77 4.5005
R2339 VSS.n228 VSS.n77 4.5005
R2340 VSS.n159 VSS.n77 4.5005
R2341 VSS.n229 VSS.n77 4.5005
R2342 VSS.n158 VSS.n77 4.5005
R2343 VSS.n230 VSS.n77 4.5005
R2344 VSS.n157 VSS.n77 4.5005
R2345 VSS.n231 VSS.n77 4.5005
R2346 VSS.n156 VSS.n77 4.5005
R2347 VSS.n232 VSS.n77 4.5005
R2348 VSS.n155 VSS.n77 4.5005
R2349 VSS.n233 VSS.n77 4.5005
R2350 VSS.n154 VSS.n77 4.5005
R2351 VSS.n234 VSS.n77 4.5005
R2352 VSS.n153 VSS.n77 4.5005
R2353 VSS.n235 VSS.n77 4.5005
R2354 VSS.n4506 VSS.n77 4.5005
R2355 VSS.n236 VSS.n77 4.5005
R2356 VSS.n152 VSS.n77 4.5005
R2357 VSS.n237 VSS.n77 4.5005
R2358 VSS.n151 VSS.n77 4.5005
R2359 VSS.n238 VSS.n77 4.5005
R2360 VSS.n150 VSS.n77 4.5005
R2361 VSS.n239 VSS.n77 4.5005
R2362 VSS.n149 VSS.n77 4.5005
R2363 VSS.n240 VSS.n77 4.5005
R2364 VSS.n148 VSS.n77 4.5005
R2365 VSS.n241 VSS.n77 4.5005
R2366 VSS.n147 VSS.n77 4.5005
R2367 VSS.n242 VSS.n77 4.5005
R2368 VSS.n146 VSS.n77 4.5005
R2369 VSS.n243 VSS.n77 4.5005
R2370 VSS.n145 VSS.n77 4.5005
R2371 VSS.n244 VSS.n77 4.5005
R2372 VSS.n144 VSS.n77 4.5005
R2373 VSS.n245 VSS.n77 4.5005
R2374 VSS.n143 VSS.n77 4.5005
R2375 VSS.n246 VSS.n77 4.5005
R2376 VSS.n142 VSS.n77 4.5005
R2377 VSS.n247 VSS.n77 4.5005
R2378 VSS.n141 VSS.n77 4.5005
R2379 VSS.n248 VSS.n77 4.5005
R2380 VSS.n140 VSS.n77 4.5005
R2381 VSS.n249 VSS.n77 4.5005
R2382 VSS.n139 VSS.n77 4.5005
R2383 VSS.n250 VSS.n77 4.5005
R2384 VSS.n138 VSS.n77 4.5005
R2385 VSS.n251 VSS.n77 4.5005
R2386 VSS.n137 VSS.n77 4.5005
R2387 VSS.n252 VSS.n77 4.5005
R2388 VSS.n136 VSS.n77 4.5005
R2389 VSS.n253 VSS.n77 4.5005
R2390 VSS.n135 VSS.n77 4.5005
R2391 VSS.n254 VSS.n77 4.5005
R2392 VSS.n134 VSS.n77 4.5005
R2393 VSS.n255 VSS.n77 4.5005
R2394 VSS.n133 VSS.n77 4.5005
R2395 VSS.n256 VSS.n77 4.5005
R2396 VSS.n132 VSS.n77 4.5005
R2397 VSS.n4502 VSS.n77 4.5005
R2398 VSS.n4504 VSS.n77 4.5005
R2399 VSS.n193 VSS.n59 4.5005
R2400 VSS.n195 VSS.n59 4.5005
R2401 VSS.n192 VSS.n59 4.5005
R2402 VSS.n196 VSS.n59 4.5005
R2403 VSS.n191 VSS.n59 4.5005
R2404 VSS.n197 VSS.n59 4.5005
R2405 VSS.n190 VSS.n59 4.5005
R2406 VSS.n198 VSS.n59 4.5005
R2407 VSS.n189 VSS.n59 4.5005
R2408 VSS.n199 VSS.n59 4.5005
R2409 VSS.n188 VSS.n59 4.5005
R2410 VSS.n200 VSS.n59 4.5005
R2411 VSS.n187 VSS.n59 4.5005
R2412 VSS.n201 VSS.n59 4.5005
R2413 VSS.n186 VSS.n59 4.5005
R2414 VSS.n202 VSS.n59 4.5005
R2415 VSS.n185 VSS.n59 4.5005
R2416 VSS.n203 VSS.n59 4.5005
R2417 VSS.n184 VSS.n59 4.5005
R2418 VSS.n204 VSS.n59 4.5005
R2419 VSS.n183 VSS.n59 4.5005
R2420 VSS.n205 VSS.n59 4.5005
R2421 VSS.n182 VSS.n59 4.5005
R2422 VSS.n206 VSS.n59 4.5005
R2423 VSS.n181 VSS.n59 4.5005
R2424 VSS.n207 VSS.n59 4.5005
R2425 VSS.n180 VSS.n59 4.5005
R2426 VSS.n208 VSS.n59 4.5005
R2427 VSS.n179 VSS.n59 4.5005
R2428 VSS.n209 VSS.n59 4.5005
R2429 VSS.n178 VSS.n59 4.5005
R2430 VSS.n210 VSS.n59 4.5005
R2431 VSS.n177 VSS.n59 4.5005
R2432 VSS.n211 VSS.n59 4.5005
R2433 VSS.n176 VSS.n59 4.5005
R2434 VSS.n212 VSS.n59 4.5005
R2435 VSS.n175 VSS.n59 4.5005
R2436 VSS.n213 VSS.n59 4.5005
R2437 VSS.n174 VSS.n59 4.5005
R2438 VSS.n214 VSS.n59 4.5005
R2439 VSS.n173 VSS.n59 4.5005
R2440 VSS.n215 VSS.n59 4.5005
R2441 VSS.n172 VSS.n59 4.5005
R2442 VSS.n216 VSS.n59 4.5005
R2443 VSS.n171 VSS.n59 4.5005
R2444 VSS.n217 VSS.n59 4.5005
R2445 VSS.n170 VSS.n59 4.5005
R2446 VSS.n218 VSS.n59 4.5005
R2447 VSS.n169 VSS.n59 4.5005
R2448 VSS.n219 VSS.n59 4.5005
R2449 VSS.n168 VSS.n59 4.5005
R2450 VSS.n220 VSS.n59 4.5005
R2451 VSS.n167 VSS.n59 4.5005
R2452 VSS.n221 VSS.n59 4.5005
R2453 VSS.n166 VSS.n59 4.5005
R2454 VSS.n222 VSS.n59 4.5005
R2455 VSS.n165 VSS.n59 4.5005
R2456 VSS.n223 VSS.n59 4.5005
R2457 VSS.n164 VSS.n59 4.5005
R2458 VSS.n224 VSS.n59 4.5005
R2459 VSS.n163 VSS.n59 4.5005
R2460 VSS.n225 VSS.n59 4.5005
R2461 VSS.n162 VSS.n59 4.5005
R2462 VSS.n226 VSS.n59 4.5005
R2463 VSS.n161 VSS.n59 4.5005
R2464 VSS.n227 VSS.n59 4.5005
R2465 VSS.n160 VSS.n59 4.5005
R2466 VSS.n228 VSS.n59 4.5005
R2467 VSS.n159 VSS.n59 4.5005
R2468 VSS.n229 VSS.n59 4.5005
R2469 VSS.n158 VSS.n59 4.5005
R2470 VSS.n230 VSS.n59 4.5005
R2471 VSS.n157 VSS.n59 4.5005
R2472 VSS.n231 VSS.n59 4.5005
R2473 VSS.n156 VSS.n59 4.5005
R2474 VSS.n232 VSS.n59 4.5005
R2475 VSS.n155 VSS.n59 4.5005
R2476 VSS.n233 VSS.n59 4.5005
R2477 VSS.n154 VSS.n59 4.5005
R2478 VSS.n234 VSS.n59 4.5005
R2479 VSS.n153 VSS.n59 4.5005
R2480 VSS.n235 VSS.n59 4.5005
R2481 VSS.n4506 VSS.n59 4.5005
R2482 VSS.n236 VSS.n59 4.5005
R2483 VSS.n152 VSS.n59 4.5005
R2484 VSS.n237 VSS.n59 4.5005
R2485 VSS.n151 VSS.n59 4.5005
R2486 VSS.n238 VSS.n59 4.5005
R2487 VSS.n150 VSS.n59 4.5005
R2488 VSS.n239 VSS.n59 4.5005
R2489 VSS.n149 VSS.n59 4.5005
R2490 VSS.n240 VSS.n59 4.5005
R2491 VSS.n148 VSS.n59 4.5005
R2492 VSS.n241 VSS.n59 4.5005
R2493 VSS.n147 VSS.n59 4.5005
R2494 VSS.n242 VSS.n59 4.5005
R2495 VSS.n146 VSS.n59 4.5005
R2496 VSS.n243 VSS.n59 4.5005
R2497 VSS.n145 VSS.n59 4.5005
R2498 VSS.n244 VSS.n59 4.5005
R2499 VSS.n144 VSS.n59 4.5005
R2500 VSS.n245 VSS.n59 4.5005
R2501 VSS.n143 VSS.n59 4.5005
R2502 VSS.n246 VSS.n59 4.5005
R2503 VSS.n142 VSS.n59 4.5005
R2504 VSS.n247 VSS.n59 4.5005
R2505 VSS.n141 VSS.n59 4.5005
R2506 VSS.n248 VSS.n59 4.5005
R2507 VSS.n140 VSS.n59 4.5005
R2508 VSS.n249 VSS.n59 4.5005
R2509 VSS.n139 VSS.n59 4.5005
R2510 VSS.n250 VSS.n59 4.5005
R2511 VSS.n138 VSS.n59 4.5005
R2512 VSS.n251 VSS.n59 4.5005
R2513 VSS.n137 VSS.n59 4.5005
R2514 VSS.n252 VSS.n59 4.5005
R2515 VSS.n136 VSS.n59 4.5005
R2516 VSS.n253 VSS.n59 4.5005
R2517 VSS.n135 VSS.n59 4.5005
R2518 VSS.n254 VSS.n59 4.5005
R2519 VSS.n134 VSS.n59 4.5005
R2520 VSS.n255 VSS.n59 4.5005
R2521 VSS.n133 VSS.n59 4.5005
R2522 VSS.n256 VSS.n59 4.5005
R2523 VSS.n132 VSS.n59 4.5005
R2524 VSS.n4502 VSS.n59 4.5005
R2525 VSS.n4504 VSS.n59 4.5005
R2526 VSS.n193 VSS.n78 4.5005
R2527 VSS.n195 VSS.n78 4.5005
R2528 VSS.n192 VSS.n78 4.5005
R2529 VSS.n196 VSS.n78 4.5005
R2530 VSS.n191 VSS.n78 4.5005
R2531 VSS.n197 VSS.n78 4.5005
R2532 VSS.n190 VSS.n78 4.5005
R2533 VSS.n198 VSS.n78 4.5005
R2534 VSS.n189 VSS.n78 4.5005
R2535 VSS.n199 VSS.n78 4.5005
R2536 VSS.n188 VSS.n78 4.5005
R2537 VSS.n200 VSS.n78 4.5005
R2538 VSS.n187 VSS.n78 4.5005
R2539 VSS.n201 VSS.n78 4.5005
R2540 VSS.n186 VSS.n78 4.5005
R2541 VSS.n202 VSS.n78 4.5005
R2542 VSS.n185 VSS.n78 4.5005
R2543 VSS.n203 VSS.n78 4.5005
R2544 VSS.n184 VSS.n78 4.5005
R2545 VSS.n204 VSS.n78 4.5005
R2546 VSS.n183 VSS.n78 4.5005
R2547 VSS.n205 VSS.n78 4.5005
R2548 VSS.n182 VSS.n78 4.5005
R2549 VSS.n206 VSS.n78 4.5005
R2550 VSS.n181 VSS.n78 4.5005
R2551 VSS.n207 VSS.n78 4.5005
R2552 VSS.n180 VSS.n78 4.5005
R2553 VSS.n208 VSS.n78 4.5005
R2554 VSS.n179 VSS.n78 4.5005
R2555 VSS.n209 VSS.n78 4.5005
R2556 VSS.n178 VSS.n78 4.5005
R2557 VSS.n210 VSS.n78 4.5005
R2558 VSS.n177 VSS.n78 4.5005
R2559 VSS.n211 VSS.n78 4.5005
R2560 VSS.n176 VSS.n78 4.5005
R2561 VSS.n212 VSS.n78 4.5005
R2562 VSS.n175 VSS.n78 4.5005
R2563 VSS.n213 VSS.n78 4.5005
R2564 VSS.n174 VSS.n78 4.5005
R2565 VSS.n214 VSS.n78 4.5005
R2566 VSS.n173 VSS.n78 4.5005
R2567 VSS.n215 VSS.n78 4.5005
R2568 VSS.n172 VSS.n78 4.5005
R2569 VSS.n216 VSS.n78 4.5005
R2570 VSS.n171 VSS.n78 4.5005
R2571 VSS.n217 VSS.n78 4.5005
R2572 VSS.n170 VSS.n78 4.5005
R2573 VSS.n218 VSS.n78 4.5005
R2574 VSS.n169 VSS.n78 4.5005
R2575 VSS.n219 VSS.n78 4.5005
R2576 VSS.n168 VSS.n78 4.5005
R2577 VSS.n220 VSS.n78 4.5005
R2578 VSS.n167 VSS.n78 4.5005
R2579 VSS.n221 VSS.n78 4.5005
R2580 VSS.n166 VSS.n78 4.5005
R2581 VSS.n222 VSS.n78 4.5005
R2582 VSS.n165 VSS.n78 4.5005
R2583 VSS.n223 VSS.n78 4.5005
R2584 VSS.n164 VSS.n78 4.5005
R2585 VSS.n224 VSS.n78 4.5005
R2586 VSS.n163 VSS.n78 4.5005
R2587 VSS.n225 VSS.n78 4.5005
R2588 VSS.n162 VSS.n78 4.5005
R2589 VSS.n226 VSS.n78 4.5005
R2590 VSS.n161 VSS.n78 4.5005
R2591 VSS.n227 VSS.n78 4.5005
R2592 VSS.n160 VSS.n78 4.5005
R2593 VSS.n228 VSS.n78 4.5005
R2594 VSS.n159 VSS.n78 4.5005
R2595 VSS.n229 VSS.n78 4.5005
R2596 VSS.n158 VSS.n78 4.5005
R2597 VSS.n230 VSS.n78 4.5005
R2598 VSS.n157 VSS.n78 4.5005
R2599 VSS.n231 VSS.n78 4.5005
R2600 VSS.n156 VSS.n78 4.5005
R2601 VSS.n232 VSS.n78 4.5005
R2602 VSS.n155 VSS.n78 4.5005
R2603 VSS.n233 VSS.n78 4.5005
R2604 VSS.n154 VSS.n78 4.5005
R2605 VSS.n234 VSS.n78 4.5005
R2606 VSS.n153 VSS.n78 4.5005
R2607 VSS.n235 VSS.n78 4.5005
R2608 VSS.n4506 VSS.n78 4.5005
R2609 VSS.n236 VSS.n78 4.5005
R2610 VSS.n152 VSS.n78 4.5005
R2611 VSS.n237 VSS.n78 4.5005
R2612 VSS.n151 VSS.n78 4.5005
R2613 VSS.n238 VSS.n78 4.5005
R2614 VSS.n150 VSS.n78 4.5005
R2615 VSS.n239 VSS.n78 4.5005
R2616 VSS.n149 VSS.n78 4.5005
R2617 VSS.n240 VSS.n78 4.5005
R2618 VSS.n148 VSS.n78 4.5005
R2619 VSS.n241 VSS.n78 4.5005
R2620 VSS.n147 VSS.n78 4.5005
R2621 VSS.n242 VSS.n78 4.5005
R2622 VSS.n146 VSS.n78 4.5005
R2623 VSS.n243 VSS.n78 4.5005
R2624 VSS.n145 VSS.n78 4.5005
R2625 VSS.n244 VSS.n78 4.5005
R2626 VSS.n144 VSS.n78 4.5005
R2627 VSS.n245 VSS.n78 4.5005
R2628 VSS.n143 VSS.n78 4.5005
R2629 VSS.n246 VSS.n78 4.5005
R2630 VSS.n142 VSS.n78 4.5005
R2631 VSS.n247 VSS.n78 4.5005
R2632 VSS.n141 VSS.n78 4.5005
R2633 VSS.n248 VSS.n78 4.5005
R2634 VSS.n140 VSS.n78 4.5005
R2635 VSS.n249 VSS.n78 4.5005
R2636 VSS.n139 VSS.n78 4.5005
R2637 VSS.n250 VSS.n78 4.5005
R2638 VSS.n138 VSS.n78 4.5005
R2639 VSS.n251 VSS.n78 4.5005
R2640 VSS.n137 VSS.n78 4.5005
R2641 VSS.n252 VSS.n78 4.5005
R2642 VSS.n136 VSS.n78 4.5005
R2643 VSS.n253 VSS.n78 4.5005
R2644 VSS.n135 VSS.n78 4.5005
R2645 VSS.n254 VSS.n78 4.5005
R2646 VSS.n134 VSS.n78 4.5005
R2647 VSS.n255 VSS.n78 4.5005
R2648 VSS.n133 VSS.n78 4.5005
R2649 VSS.n256 VSS.n78 4.5005
R2650 VSS.n132 VSS.n78 4.5005
R2651 VSS.n4502 VSS.n78 4.5005
R2652 VSS.n4504 VSS.n78 4.5005
R2653 VSS.n193 VSS.n58 4.5005
R2654 VSS.n195 VSS.n58 4.5005
R2655 VSS.n192 VSS.n58 4.5005
R2656 VSS.n196 VSS.n58 4.5005
R2657 VSS.n191 VSS.n58 4.5005
R2658 VSS.n197 VSS.n58 4.5005
R2659 VSS.n190 VSS.n58 4.5005
R2660 VSS.n198 VSS.n58 4.5005
R2661 VSS.n189 VSS.n58 4.5005
R2662 VSS.n199 VSS.n58 4.5005
R2663 VSS.n188 VSS.n58 4.5005
R2664 VSS.n200 VSS.n58 4.5005
R2665 VSS.n187 VSS.n58 4.5005
R2666 VSS.n201 VSS.n58 4.5005
R2667 VSS.n186 VSS.n58 4.5005
R2668 VSS.n202 VSS.n58 4.5005
R2669 VSS.n185 VSS.n58 4.5005
R2670 VSS.n203 VSS.n58 4.5005
R2671 VSS.n184 VSS.n58 4.5005
R2672 VSS.n204 VSS.n58 4.5005
R2673 VSS.n183 VSS.n58 4.5005
R2674 VSS.n205 VSS.n58 4.5005
R2675 VSS.n182 VSS.n58 4.5005
R2676 VSS.n206 VSS.n58 4.5005
R2677 VSS.n181 VSS.n58 4.5005
R2678 VSS.n207 VSS.n58 4.5005
R2679 VSS.n180 VSS.n58 4.5005
R2680 VSS.n208 VSS.n58 4.5005
R2681 VSS.n179 VSS.n58 4.5005
R2682 VSS.n209 VSS.n58 4.5005
R2683 VSS.n178 VSS.n58 4.5005
R2684 VSS.n210 VSS.n58 4.5005
R2685 VSS.n177 VSS.n58 4.5005
R2686 VSS.n211 VSS.n58 4.5005
R2687 VSS.n176 VSS.n58 4.5005
R2688 VSS.n212 VSS.n58 4.5005
R2689 VSS.n175 VSS.n58 4.5005
R2690 VSS.n213 VSS.n58 4.5005
R2691 VSS.n174 VSS.n58 4.5005
R2692 VSS.n214 VSS.n58 4.5005
R2693 VSS.n173 VSS.n58 4.5005
R2694 VSS.n215 VSS.n58 4.5005
R2695 VSS.n172 VSS.n58 4.5005
R2696 VSS.n216 VSS.n58 4.5005
R2697 VSS.n171 VSS.n58 4.5005
R2698 VSS.n217 VSS.n58 4.5005
R2699 VSS.n170 VSS.n58 4.5005
R2700 VSS.n218 VSS.n58 4.5005
R2701 VSS.n169 VSS.n58 4.5005
R2702 VSS.n219 VSS.n58 4.5005
R2703 VSS.n168 VSS.n58 4.5005
R2704 VSS.n220 VSS.n58 4.5005
R2705 VSS.n167 VSS.n58 4.5005
R2706 VSS.n221 VSS.n58 4.5005
R2707 VSS.n166 VSS.n58 4.5005
R2708 VSS.n222 VSS.n58 4.5005
R2709 VSS.n165 VSS.n58 4.5005
R2710 VSS.n223 VSS.n58 4.5005
R2711 VSS.n164 VSS.n58 4.5005
R2712 VSS.n224 VSS.n58 4.5005
R2713 VSS.n163 VSS.n58 4.5005
R2714 VSS.n225 VSS.n58 4.5005
R2715 VSS.n162 VSS.n58 4.5005
R2716 VSS.n226 VSS.n58 4.5005
R2717 VSS.n161 VSS.n58 4.5005
R2718 VSS.n227 VSS.n58 4.5005
R2719 VSS.n160 VSS.n58 4.5005
R2720 VSS.n228 VSS.n58 4.5005
R2721 VSS.n159 VSS.n58 4.5005
R2722 VSS.n229 VSS.n58 4.5005
R2723 VSS.n158 VSS.n58 4.5005
R2724 VSS.n230 VSS.n58 4.5005
R2725 VSS.n157 VSS.n58 4.5005
R2726 VSS.n231 VSS.n58 4.5005
R2727 VSS.n156 VSS.n58 4.5005
R2728 VSS.n232 VSS.n58 4.5005
R2729 VSS.n155 VSS.n58 4.5005
R2730 VSS.n233 VSS.n58 4.5005
R2731 VSS.n154 VSS.n58 4.5005
R2732 VSS.n234 VSS.n58 4.5005
R2733 VSS.n153 VSS.n58 4.5005
R2734 VSS.n235 VSS.n58 4.5005
R2735 VSS.n4506 VSS.n58 4.5005
R2736 VSS.n236 VSS.n58 4.5005
R2737 VSS.n152 VSS.n58 4.5005
R2738 VSS.n237 VSS.n58 4.5005
R2739 VSS.n151 VSS.n58 4.5005
R2740 VSS.n238 VSS.n58 4.5005
R2741 VSS.n150 VSS.n58 4.5005
R2742 VSS.n239 VSS.n58 4.5005
R2743 VSS.n149 VSS.n58 4.5005
R2744 VSS.n240 VSS.n58 4.5005
R2745 VSS.n148 VSS.n58 4.5005
R2746 VSS.n241 VSS.n58 4.5005
R2747 VSS.n147 VSS.n58 4.5005
R2748 VSS.n242 VSS.n58 4.5005
R2749 VSS.n146 VSS.n58 4.5005
R2750 VSS.n243 VSS.n58 4.5005
R2751 VSS.n145 VSS.n58 4.5005
R2752 VSS.n244 VSS.n58 4.5005
R2753 VSS.n144 VSS.n58 4.5005
R2754 VSS.n245 VSS.n58 4.5005
R2755 VSS.n143 VSS.n58 4.5005
R2756 VSS.n246 VSS.n58 4.5005
R2757 VSS.n142 VSS.n58 4.5005
R2758 VSS.n247 VSS.n58 4.5005
R2759 VSS.n141 VSS.n58 4.5005
R2760 VSS.n248 VSS.n58 4.5005
R2761 VSS.n140 VSS.n58 4.5005
R2762 VSS.n249 VSS.n58 4.5005
R2763 VSS.n139 VSS.n58 4.5005
R2764 VSS.n250 VSS.n58 4.5005
R2765 VSS.n138 VSS.n58 4.5005
R2766 VSS.n251 VSS.n58 4.5005
R2767 VSS.n137 VSS.n58 4.5005
R2768 VSS.n252 VSS.n58 4.5005
R2769 VSS.n136 VSS.n58 4.5005
R2770 VSS.n253 VSS.n58 4.5005
R2771 VSS.n135 VSS.n58 4.5005
R2772 VSS.n254 VSS.n58 4.5005
R2773 VSS.n134 VSS.n58 4.5005
R2774 VSS.n255 VSS.n58 4.5005
R2775 VSS.n133 VSS.n58 4.5005
R2776 VSS.n256 VSS.n58 4.5005
R2777 VSS.n132 VSS.n58 4.5005
R2778 VSS.n4502 VSS.n58 4.5005
R2779 VSS.n4504 VSS.n58 4.5005
R2780 VSS.n193 VSS.n79 4.5005
R2781 VSS.n195 VSS.n79 4.5005
R2782 VSS.n192 VSS.n79 4.5005
R2783 VSS.n196 VSS.n79 4.5005
R2784 VSS.n191 VSS.n79 4.5005
R2785 VSS.n197 VSS.n79 4.5005
R2786 VSS.n190 VSS.n79 4.5005
R2787 VSS.n198 VSS.n79 4.5005
R2788 VSS.n189 VSS.n79 4.5005
R2789 VSS.n199 VSS.n79 4.5005
R2790 VSS.n188 VSS.n79 4.5005
R2791 VSS.n200 VSS.n79 4.5005
R2792 VSS.n187 VSS.n79 4.5005
R2793 VSS.n201 VSS.n79 4.5005
R2794 VSS.n186 VSS.n79 4.5005
R2795 VSS.n202 VSS.n79 4.5005
R2796 VSS.n185 VSS.n79 4.5005
R2797 VSS.n203 VSS.n79 4.5005
R2798 VSS.n184 VSS.n79 4.5005
R2799 VSS.n204 VSS.n79 4.5005
R2800 VSS.n183 VSS.n79 4.5005
R2801 VSS.n205 VSS.n79 4.5005
R2802 VSS.n182 VSS.n79 4.5005
R2803 VSS.n206 VSS.n79 4.5005
R2804 VSS.n181 VSS.n79 4.5005
R2805 VSS.n207 VSS.n79 4.5005
R2806 VSS.n180 VSS.n79 4.5005
R2807 VSS.n208 VSS.n79 4.5005
R2808 VSS.n179 VSS.n79 4.5005
R2809 VSS.n209 VSS.n79 4.5005
R2810 VSS.n178 VSS.n79 4.5005
R2811 VSS.n210 VSS.n79 4.5005
R2812 VSS.n177 VSS.n79 4.5005
R2813 VSS.n211 VSS.n79 4.5005
R2814 VSS.n176 VSS.n79 4.5005
R2815 VSS.n212 VSS.n79 4.5005
R2816 VSS.n175 VSS.n79 4.5005
R2817 VSS.n213 VSS.n79 4.5005
R2818 VSS.n174 VSS.n79 4.5005
R2819 VSS.n214 VSS.n79 4.5005
R2820 VSS.n173 VSS.n79 4.5005
R2821 VSS.n215 VSS.n79 4.5005
R2822 VSS.n172 VSS.n79 4.5005
R2823 VSS.n216 VSS.n79 4.5005
R2824 VSS.n171 VSS.n79 4.5005
R2825 VSS.n217 VSS.n79 4.5005
R2826 VSS.n170 VSS.n79 4.5005
R2827 VSS.n218 VSS.n79 4.5005
R2828 VSS.n169 VSS.n79 4.5005
R2829 VSS.n219 VSS.n79 4.5005
R2830 VSS.n168 VSS.n79 4.5005
R2831 VSS.n220 VSS.n79 4.5005
R2832 VSS.n167 VSS.n79 4.5005
R2833 VSS.n221 VSS.n79 4.5005
R2834 VSS.n166 VSS.n79 4.5005
R2835 VSS.n222 VSS.n79 4.5005
R2836 VSS.n165 VSS.n79 4.5005
R2837 VSS.n223 VSS.n79 4.5005
R2838 VSS.n164 VSS.n79 4.5005
R2839 VSS.n224 VSS.n79 4.5005
R2840 VSS.n163 VSS.n79 4.5005
R2841 VSS.n225 VSS.n79 4.5005
R2842 VSS.n162 VSS.n79 4.5005
R2843 VSS.n226 VSS.n79 4.5005
R2844 VSS.n161 VSS.n79 4.5005
R2845 VSS.n227 VSS.n79 4.5005
R2846 VSS.n160 VSS.n79 4.5005
R2847 VSS.n228 VSS.n79 4.5005
R2848 VSS.n159 VSS.n79 4.5005
R2849 VSS.n229 VSS.n79 4.5005
R2850 VSS.n158 VSS.n79 4.5005
R2851 VSS.n230 VSS.n79 4.5005
R2852 VSS.n157 VSS.n79 4.5005
R2853 VSS.n231 VSS.n79 4.5005
R2854 VSS.n156 VSS.n79 4.5005
R2855 VSS.n232 VSS.n79 4.5005
R2856 VSS.n155 VSS.n79 4.5005
R2857 VSS.n233 VSS.n79 4.5005
R2858 VSS.n154 VSS.n79 4.5005
R2859 VSS.n234 VSS.n79 4.5005
R2860 VSS.n153 VSS.n79 4.5005
R2861 VSS.n235 VSS.n79 4.5005
R2862 VSS.n4506 VSS.n79 4.5005
R2863 VSS.n236 VSS.n79 4.5005
R2864 VSS.n152 VSS.n79 4.5005
R2865 VSS.n237 VSS.n79 4.5005
R2866 VSS.n151 VSS.n79 4.5005
R2867 VSS.n238 VSS.n79 4.5005
R2868 VSS.n150 VSS.n79 4.5005
R2869 VSS.n239 VSS.n79 4.5005
R2870 VSS.n149 VSS.n79 4.5005
R2871 VSS.n240 VSS.n79 4.5005
R2872 VSS.n148 VSS.n79 4.5005
R2873 VSS.n241 VSS.n79 4.5005
R2874 VSS.n147 VSS.n79 4.5005
R2875 VSS.n242 VSS.n79 4.5005
R2876 VSS.n146 VSS.n79 4.5005
R2877 VSS.n243 VSS.n79 4.5005
R2878 VSS.n145 VSS.n79 4.5005
R2879 VSS.n244 VSS.n79 4.5005
R2880 VSS.n144 VSS.n79 4.5005
R2881 VSS.n245 VSS.n79 4.5005
R2882 VSS.n143 VSS.n79 4.5005
R2883 VSS.n246 VSS.n79 4.5005
R2884 VSS.n142 VSS.n79 4.5005
R2885 VSS.n247 VSS.n79 4.5005
R2886 VSS.n141 VSS.n79 4.5005
R2887 VSS.n248 VSS.n79 4.5005
R2888 VSS.n140 VSS.n79 4.5005
R2889 VSS.n249 VSS.n79 4.5005
R2890 VSS.n139 VSS.n79 4.5005
R2891 VSS.n250 VSS.n79 4.5005
R2892 VSS.n138 VSS.n79 4.5005
R2893 VSS.n251 VSS.n79 4.5005
R2894 VSS.n137 VSS.n79 4.5005
R2895 VSS.n252 VSS.n79 4.5005
R2896 VSS.n136 VSS.n79 4.5005
R2897 VSS.n253 VSS.n79 4.5005
R2898 VSS.n135 VSS.n79 4.5005
R2899 VSS.n254 VSS.n79 4.5005
R2900 VSS.n134 VSS.n79 4.5005
R2901 VSS.n255 VSS.n79 4.5005
R2902 VSS.n133 VSS.n79 4.5005
R2903 VSS.n256 VSS.n79 4.5005
R2904 VSS.n132 VSS.n79 4.5005
R2905 VSS.n4502 VSS.n79 4.5005
R2906 VSS.n4504 VSS.n79 4.5005
R2907 VSS.n193 VSS.n57 4.5005
R2908 VSS.n195 VSS.n57 4.5005
R2909 VSS.n192 VSS.n57 4.5005
R2910 VSS.n196 VSS.n57 4.5005
R2911 VSS.n191 VSS.n57 4.5005
R2912 VSS.n197 VSS.n57 4.5005
R2913 VSS.n190 VSS.n57 4.5005
R2914 VSS.n198 VSS.n57 4.5005
R2915 VSS.n189 VSS.n57 4.5005
R2916 VSS.n199 VSS.n57 4.5005
R2917 VSS.n188 VSS.n57 4.5005
R2918 VSS.n200 VSS.n57 4.5005
R2919 VSS.n187 VSS.n57 4.5005
R2920 VSS.n201 VSS.n57 4.5005
R2921 VSS.n186 VSS.n57 4.5005
R2922 VSS.n202 VSS.n57 4.5005
R2923 VSS.n185 VSS.n57 4.5005
R2924 VSS.n203 VSS.n57 4.5005
R2925 VSS.n184 VSS.n57 4.5005
R2926 VSS.n204 VSS.n57 4.5005
R2927 VSS.n183 VSS.n57 4.5005
R2928 VSS.n205 VSS.n57 4.5005
R2929 VSS.n182 VSS.n57 4.5005
R2930 VSS.n206 VSS.n57 4.5005
R2931 VSS.n181 VSS.n57 4.5005
R2932 VSS.n207 VSS.n57 4.5005
R2933 VSS.n180 VSS.n57 4.5005
R2934 VSS.n208 VSS.n57 4.5005
R2935 VSS.n179 VSS.n57 4.5005
R2936 VSS.n209 VSS.n57 4.5005
R2937 VSS.n178 VSS.n57 4.5005
R2938 VSS.n210 VSS.n57 4.5005
R2939 VSS.n177 VSS.n57 4.5005
R2940 VSS.n211 VSS.n57 4.5005
R2941 VSS.n176 VSS.n57 4.5005
R2942 VSS.n212 VSS.n57 4.5005
R2943 VSS.n175 VSS.n57 4.5005
R2944 VSS.n213 VSS.n57 4.5005
R2945 VSS.n174 VSS.n57 4.5005
R2946 VSS.n214 VSS.n57 4.5005
R2947 VSS.n173 VSS.n57 4.5005
R2948 VSS.n215 VSS.n57 4.5005
R2949 VSS.n172 VSS.n57 4.5005
R2950 VSS.n216 VSS.n57 4.5005
R2951 VSS.n171 VSS.n57 4.5005
R2952 VSS.n217 VSS.n57 4.5005
R2953 VSS.n170 VSS.n57 4.5005
R2954 VSS.n218 VSS.n57 4.5005
R2955 VSS.n169 VSS.n57 4.5005
R2956 VSS.n219 VSS.n57 4.5005
R2957 VSS.n168 VSS.n57 4.5005
R2958 VSS.n220 VSS.n57 4.5005
R2959 VSS.n167 VSS.n57 4.5005
R2960 VSS.n221 VSS.n57 4.5005
R2961 VSS.n166 VSS.n57 4.5005
R2962 VSS.n222 VSS.n57 4.5005
R2963 VSS.n165 VSS.n57 4.5005
R2964 VSS.n223 VSS.n57 4.5005
R2965 VSS.n164 VSS.n57 4.5005
R2966 VSS.n224 VSS.n57 4.5005
R2967 VSS.n163 VSS.n57 4.5005
R2968 VSS.n225 VSS.n57 4.5005
R2969 VSS.n162 VSS.n57 4.5005
R2970 VSS.n226 VSS.n57 4.5005
R2971 VSS.n161 VSS.n57 4.5005
R2972 VSS.n227 VSS.n57 4.5005
R2973 VSS.n160 VSS.n57 4.5005
R2974 VSS.n228 VSS.n57 4.5005
R2975 VSS.n159 VSS.n57 4.5005
R2976 VSS.n229 VSS.n57 4.5005
R2977 VSS.n158 VSS.n57 4.5005
R2978 VSS.n230 VSS.n57 4.5005
R2979 VSS.n157 VSS.n57 4.5005
R2980 VSS.n231 VSS.n57 4.5005
R2981 VSS.n156 VSS.n57 4.5005
R2982 VSS.n232 VSS.n57 4.5005
R2983 VSS.n155 VSS.n57 4.5005
R2984 VSS.n233 VSS.n57 4.5005
R2985 VSS.n154 VSS.n57 4.5005
R2986 VSS.n234 VSS.n57 4.5005
R2987 VSS.n153 VSS.n57 4.5005
R2988 VSS.n235 VSS.n57 4.5005
R2989 VSS.n4506 VSS.n57 4.5005
R2990 VSS.n236 VSS.n57 4.5005
R2991 VSS.n152 VSS.n57 4.5005
R2992 VSS.n237 VSS.n57 4.5005
R2993 VSS.n151 VSS.n57 4.5005
R2994 VSS.n238 VSS.n57 4.5005
R2995 VSS.n150 VSS.n57 4.5005
R2996 VSS.n239 VSS.n57 4.5005
R2997 VSS.n149 VSS.n57 4.5005
R2998 VSS.n240 VSS.n57 4.5005
R2999 VSS.n148 VSS.n57 4.5005
R3000 VSS.n241 VSS.n57 4.5005
R3001 VSS.n147 VSS.n57 4.5005
R3002 VSS.n242 VSS.n57 4.5005
R3003 VSS.n146 VSS.n57 4.5005
R3004 VSS.n243 VSS.n57 4.5005
R3005 VSS.n145 VSS.n57 4.5005
R3006 VSS.n244 VSS.n57 4.5005
R3007 VSS.n144 VSS.n57 4.5005
R3008 VSS.n245 VSS.n57 4.5005
R3009 VSS.n143 VSS.n57 4.5005
R3010 VSS.n246 VSS.n57 4.5005
R3011 VSS.n142 VSS.n57 4.5005
R3012 VSS.n247 VSS.n57 4.5005
R3013 VSS.n141 VSS.n57 4.5005
R3014 VSS.n248 VSS.n57 4.5005
R3015 VSS.n140 VSS.n57 4.5005
R3016 VSS.n249 VSS.n57 4.5005
R3017 VSS.n139 VSS.n57 4.5005
R3018 VSS.n250 VSS.n57 4.5005
R3019 VSS.n138 VSS.n57 4.5005
R3020 VSS.n251 VSS.n57 4.5005
R3021 VSS.n137 VSS.n57 4.5005
R3022 VSS.n252 VSS.n57 4.5005
R3023 VSS.n136 VSS.n57 4.5005
R3024 VSS.n253 VSS.n57 4.5005
R3025 VSS.n135 VSS.n57 4.5005
R3026 VSS.n254 VSS.n57 4.5005
R3027 VSS.n134 VSS.n57 4.5005
R3028 VSS.n255 VSS.n57 4.5005
R3029 VSS.n133 VSS.n57 4.5005
R3030 VSS.n256 VSS.n57 4.5005
R3031 VSS.n132 VSS.n57 4.5005
R3032 VSS.n4502 VSS.n57 4.5005
R3033 VSS.n4504 VSS.n57 4.5005
R3034 VSS.n193 VSS.n80 4.5005
R3035 VSS.n195 VSS.n80 4.5005
R3036 VSS.n192 VSS.n80 4.5005
R3037 VSS.n196 VSS.n80 4.5005
R3038 VSS.n191 VSS.n80 4.5005
R3039 VSS.n197 VSS.n80 4.5005
R3040 VSS.n190 VSS.n80 4.5005
R3041 VSS.n198 VSS.n80 4.5005
R3042 VSS.n189 VSS.n80 4.5005
R3043 VSS.n199 VSS.n80 4.5005
R3044 VSS.n188 VSS.n80 4.5005
R3045 VSS.n200 VSS.n80 4.5005
R3046 VSS.n187 VSS.n80 4.5005
R3047 VSS.n201 VSS.n80 4.5005
R3048 VSS.n186 VSS.n80 4.5005
R3049 VSS.n202 VSS.n80 4.5005
R3050 VSS.n185 VSS.n80 4.5005
R3051 VSS.n203 VSS.n80 4.5005
R3052 VSS.n184 VSS.n80 4.5005
R3053 VSS.n204 VSS.n80 4.5005
R3054 VSS.n183 VSS.n80 4.5005
R3055 VSS.n205 VSS.n80 4.5005
R3056 VSS.n182 VSS.n80 4.5005
R3057 VSS.n206 VSS.n80 4.5005
R3058 VSS.n181 VSS.n80 4.5005
R3059 VSS.n207 VSS.n80 4.5005
R3060 VSS.n180 VSS.n80 4.5005
R3061 VSS.n208 VSS.n80 4.5005
R3062 VSS.n179 VSS.n80 4.5005
R3063 VSS.n209 VSS.n80 4.5005
R3064 VSS.n178 VSS.n80 4.5005
R3065 VSS.n210 VSS.n80 4.5005
R3066 VSS.n177 VSS.n80 4.5005
R3067 VSS.n211 VSS.n80 4.5005
R3068 VSS.n176 VSS.n80 4.5005
R3069 VSS.n212 VSS.n80 4.5005
R3070 VSS.n175 VSS.n80 4.5005
R3071 VSS.n213 VSS.n80 4.5005
R3072 VSS.n174 VSS.n80 4.5005
R3073 VSS.n214 VSS.n80 4.5005
R3074 VSS.n173 VSS.n80 4.5005
R3075 VSS.n215 VSS.n80 4.5005
R3076 VSS.n172 VSS.n80 4.5005
R3077 VSS.n216 VSS.n80 4.5005
R3078 VSS.n171 VSS.n80 4.5005
R3079 VSS.n217 VSS.n80 4.5005
R3080 VSS.n170 VSS.n80 4.5005
R3081 VSS.n218 VSS.n80 4.5005
R3082 VSS.n169 VSS.n80 4.5005
R3083 VSS.n219 VSS.n80 4.5005
R3084 VSS.n168 VSS.n80 4.5005
R3085 VSS.n220 VSS.n80 4.5005
R3086 VSS.n167 VSS.n80 4.5005
R3087 VSS.n221 VSS.n80 4.5005
R3088 VSS.n166 VSS.n80 4.5005
R3089 VSS.n222 VSS.n80 4.5005
R3090 VSS.n165 VSS.n80 4.5005
R3091 VSS.n223 VSS.n80 4.5005
R3092 VSS.n164 VSS.n80 4.5005
R3093 VSS.n224 VSS.n80 4.5005
R3094 VSS.n163 VSS.n80 4.5005
R3095 VSS.n225 VSS.n80 4.5005
R3096 VSS.n162 VSS.n80 4.5005
R3097 VSS.n226 VSS.n80 4.5005
R3098 VSS.n161 VSS.n80 4.5005
R3099 VSS.n227 VSS.n80 4.5005
R3100 VSS.n160 VSS.n80 4.5005
R3101 VSS.n228 VSS.n80 4.5005
R3102 VSS.n159 VSS.n80 4.5005
R3103 VSS.n229 VSS.n80 4.5005
R3104 VSS.n158 VSS.n80 4.5005
R3105 VSS.n230 VSS.n80 4.5005
R3106 VSS.n157 VSS.n80 4.5005
R3107 VSS.n231 VSS.n80 4.5005
R3108 VSS.n156 VSS.n80 4.5005
R3109 VSS.n232 VSS.n80 4.5005
R3110 VSS.n155 VSS.n80 4.5005
R3111 VSS.n233 VSS.n80 4.5005
R3112 VSS.n154 VSS.n80 4.5005
R3113 VSS.n234 VSS.n80 4.5005
R3114 VSS.n153 VSS.n80 4.5005
R3115 VSS.n235 VSS.n80 4.5005
R3116 VSS.n4506 VSS.n80 4.5005
R3117 VSS.n236 VSS.n80 4.5005
R3118 VSS.n152 VSS.n80 4.5005
R3119 VSS.n237 VSS.n80 4.5005
R3120 VSS.n151 VSS.n80 4.5005
R3121 VSS.n238 VSS.n80 4.5005
R3122 VSS.n150 VSS.n80 4.5005
R3123 VSS.n239 VSS.n80 4.5005
R3124 VSS.n149 VSS.n80 4.5005
R3125 VSS.n240 VSS.n80 4.5005
R3126 VSS.n148 VSS.n80 4.5005
R3127 VSS.n241 VSS.n80 4.5005
R3128 VSS.n147 VSS.n80 4.5005
R3129 VSS.n242 VSS.n80 4.5005
R3130 VSS.n146 VSS.n80 4.5005
R3131 VSS.n243 VSS.n80 4.5005
R3132 VSS.n145 VSS.n80 4.5005
R3133 VSS.n244 VSS.n80 4.5005
R3134 VSS.n144 VSS.n80 4.5005
R3135 VSS.n245 VSS.n80 4.5005
R3136 VSS.n143 VSS.n80 4.5005
R3137 VSS.n246 VSS.n80 4.5005
R3138 VSS.n142 VSS.n80 4.5005
R3139 VSS.n247 VSS.n80 4.5005
R3140 VSS.n141 VSS.n80 4.5005
R3141 VSS.n248 VSS.n80 4.5005
R3142 VSS.n140 VSS.n80 4.5005
R3143 VSS.n249 VSS.n80 4.5005
R3144 VSS.n139 VSS.n80 4.5005
R3145 VSS.n250 VSS.n80 4.5005
R3146 VSS.n138 VSS.n80 4.5005
R3147 VSS.n251 VSS.n80 4.5005
R3148 VSS.n137 VSS.n80 4.5005
R3149 VSS.n252 VSS.n80 4.5005
R3150 VSS.n136 VSS.n80 4.5005
R3151 VSS.n253 VSS.n80 4.5005
R3152 VSS.n135 VSS.n80 4.5005
R3153 VSS.n254 VSS.n80 4.5005
R3154 VSS.n134 VSS.n80 4.5005
R3155 VSS.n255 VSS.n80 4.5005
R3156 VSS.n133 VSS.n80 4.5005
R3157 VSS.n256 VSS.n80 4.5005
R3158 VSS.n132 VSS.n80 4.5005
R3159 VSS.n4502 VSS.n80 4.5005
R3160 VSS.n4504 VSS.n80 4.5005
R3161 VSS.n193 VSS.n56 4.5005
R3162 VSS.n195 VSS.n56 4.5005
R3163 VSS.n192 VSS.n56 4.5005
R3164 VSS.n196 VSS.n56 4.5005
R3165 VSS.n191 VSS.n56 4.5005
R3166 VSS.n197 VSS.n56 4.5005
R3167 VSS.n190 VSS.n56 4.5005
R3168 VSS.n198 VSS.n56 4.5005
R3169 VSS.n189 VSS.n56 4.5005
R3170 VSS.n199 VSS.n56 4.5005
R3171 VSS.n188 VSS.n56 4.5005
R3172 VSS.n200 VSS.n56 4.5005
R3173 VSS.n187 VSS.n56 4.5005
R3174 VSS.n201 VSS.n56 4.5005
R3175 VSS.n186 VSS.n56 4.5005
R3176 VSS.n202 VSS.n56 4.5005
R3177 VSS.n185 VSS.n56 4.5005
R3178 VSS.n203 VSS.n56 4.5005
R3179 VSS.n184 VSS.n56 4.5005
R3180 VSS.n204 VSS.n56 4.5005
R3181 VSS.n183 VSS.n56 4.5005
R3182 VSS.n205 VSS.n56 4.5005
R3183 VSS.n182 VSS.n56 4.5005
R3184 VSS.n206 VSS.n56 4.5005
R3185 VSS.n181 VSS.n56 4.5005
R3186 VSS.n207 VSS.n56 4.5005
R3187 VSS.n180 VSS.n56 4.5005
R3188 VSS.n208 VSS.n56 4.5005
R3189 VSS.n179 VSS.n56 4.5005
R3190 VSS.n209 VSS.n56 4.5005
R3191 VSS.n178 VSS.n56 4.5005
R3192 VSS.n210 VSS.n56 4.5005
R3193 VSS.n177 VSS.n56 4.5005
R3194 VSS.n211 VSS.n56 4.5005
R3195 VSS.n176 VSS.n56 4.5005
R3196 VSS.n212 VSS.n56 4.5005
R3197 VSS.n175 VSS.n56 4.5005
R3198 VSS.n213 VSS.n56 4.5005
R3199 VSS.n174 VSS.n56 4.5005
R3200 VSS.n214 VSS.n56 4.5005
R3201 VSS.n173 VSS.n56 4.5005
R3202 VSS.n215 VSS.n56 4.5005
R3203 VSS.n172 VSS.n56 4.5005
R3204 VSS.n216 VSS.n56 4.5005
R3205 VSS.n171 VSS.n56 4.5005
R3206 VSS.n217 VSS.n56 4.5005
R3207 VSS.n170 VSS.n56 4.5005
R3208 VSS.n218 VSS.n56 4.5005
R3209 VSS.n169 VSS.n56 4.5005
R3210 VSS.n219 VSS.n56 4.5005
R3211 VSS.n168 VSS.n56 4.5005
R3212 VSS.n220 VSS.n56 4.5005
R3213 VSS.n167 VSS.n56 4.5005
R3214 VSS.n221 VSS.n56 4.5005
R3215 VSS.n166 VSS.n56 4.5005
R3216 VSS.n222 VSS.n56 4.5005
R3217 VSS.n165 VSS.n56 4.5005
R3218 VSS.n223 VSS.n56 4.5005
R3219 VSS.n164 VSS.n56 4.5005
R3220 VSS.n224 VSS.n56 4.5005
R3221 VSS.n163 VSS.n56 4.5005
R3222 VSS.n225 VSS.n56 4.5005
R3223 VSS.n162 VSS.n56 4.5005
R3224 VSS.n226 VSS.n56 4.5005
R3225 VSS.n161 VSS.n56 4.5005
R3226 VSS.n227 VSS.n56 4.5005
R3227 VSS.n160 VSS.n56 4.5005
R3228 VSS.n228 VSS.n56 4.5005
R3229 VSS.n159 VSS.n56 4.5005
R3230 VSS.n229 VSS.n56 4.5005
R3231 VSS.n158 VSS.n56 4.5005
R3232 VSS.n230 VSS.n56 4.5005
R3233 VSS.n157 VSS.n56 4.5005
R3234 VSS.n231 VSS.n56 4.5005
R3235 VSS.n156 VSS.n56 4.5005
R3236 VSS.n232 VSS.n56 4.5005
R3237 VSS.n155 VSS.n56 4.5005
R3238 VSS.n233 VSS.n56 4.5005
R3239 VSS.n154 VSS.n56 4.5005
R3240 VSS.n234 VSS.n56 4.5005
R3241 VSS.n153 VSS.n56 4.5005
R3242 VSS.n235 VSS.n56 4.5005
R3243 VSS.n4506 VSS.n56 4.5005
R3244 VSS.n236 VSS.n56 4.5005
R3245 VSS.n152 VSS.n56 4.5005
R3246 VSS.n237 VSS.n56 4.5005
R3247 VSS.n151 VSS.n56 4.5005
R3248 VSS.n238 VSS.n56 4.5005
R3249 VSS.n150 VSS.n56 4.5005
R3250 VSS.n239 VSS.n56 4.5005
R3251 VSS.n149 VSS.n56 4.5005
R3252 VSS.n240 VSS.n56 4.5005
R3253 VSS.n148 VSS.n56 4.5005
R3254 VSS.n241 VSS.n56 4.5005
R3255 VSS.n147 VSS.n56 4.5005
R3256 VSS.n242 VSS.n56 4.5005
R3257 VSS.n146 VSS.n56 4.5005
R3258 VSS.n243 VSS.n56 4.5005
R3259 VSS.n145 VSS.n56 4.5005
R3260 VSS.n244 VSS.n56 4.5005
R3261 VSS.n144 VSS.n56 4.5005
R3262 VSS.n245 VSS.n56 4.5005
R3263 VSS.n143 VSS.n56 4.5005
R3264 VSS.n246 VSS.n56 4.5005
R3265 VSS.n142 VSS.n56 4.5005
R3266 VSS.n247 VSS.n56 4.5005
R3267 VSS.n141 VSS.n56 4.5005
R3268 VSS.n248 VSS.n56 4.5005
R3269 VSS.n140 VSS.n56 4.5005
R3270 VSS.n249 VSS.n56 4.5005
R3271 VSS.n139 VSS.n56 4.5005
R3272 VSS.n250 VSS.n56 4.5005
R3273 VSS.n138 VSS.n56 4.5005
R3274 VSS.n251 VSS.n56 4.5005
R3275 VSS.n137 VSS.n56 4.5005
R3276 VSS.n252 VSS.n56 4.5005
R3277 VSS.n136 VSS.n56 4.5005
R3278 VSS.n253 VSS.n56 4.5005
R3279 VSS.n135 VSS.n56 4.5005
R3280 VSS.n254 VSS.n56 4.5005
R3281 VSS.n134 VSS.n56 4.5005
R3282 VSS.n255 VSS.n56 4.5005
R3283 VSS.n133 VSS.n56 4.5005
R3284 VSS.n256 VSS.n56 4.5005
R3285 VSS.n132 VSS.n56 4.5005
R3286 VSS.n4502 VSS.n56 4.5005
R3287 VSS.n4504 VSS.n56 4.5005
R3288 VSS.n193 VSS.n81 4.5005
R3289 VSS.n195 VSS.n81 4.5005
R3290 VSS.n192 VSS.n81 4.5005
R3291 VSS.n196 VSS.n81 4.5005
R3292 VSS.n191 VSS.n81 4.5005
R3293 VSS.n197 VSS.n81 4.5005
R3294 VSS.n190 VSS.n81 4.5005
R3295 VSS.n198 VSS.n81 4.5005
R3296 VSS.n189 VSS.n81 4.5005
R3297 VSS.n199 VSS.n81 4.5005
R3298 VSS.n188 VSS.n81 4.5005
R3299 VSS.n200 VSS.n81 4.5005
R3300 VSS.n187 VSS.n81 4.5005
R3301 VSS.n201 VSS.n81 4.5005
R3302 VSS.n186 VSS.n81 4.5005
R3303 VSS.n202 VSS.n81 4.5005
R3304 VSS.n185 VSS.n81 4.5005
R3305 VSS.n203 VSS.n81 4.5005
R3306 VSS.n184 VSS.n81 4.5005
R3307 VSS.n204 VSS.n81 4.5005
R3308 VSS.n183 VSS.n81 4.5005
R3309 VSS.n205 VSS.n81 4.5005
R3310 VSS.n182 VSS.n81 4.5005
R3311 VSS.n206 VSS.n81 4.5005
R3312 VSS.n181 VSS.n81 4.5005
R3313 VSS.n207 VSS.n81 4.5005
R3314 VSS.n180 VSS.n81 4.5005
R3315 VSS.n208 VSS.n81 4.5005
R3316 VSS.n179 VSS.n81 4.5005
R3317 VSS.n209 VSS.n81 4.5005
R3318 VSS.n178 VSS.n81 4.5005
R3319 VSS.n210 VSS.n81 4.5005
R3320 VSS.n177 VSS.n81 4.5005
R3321 VSS.n211 VSS.n81 4.5005
R3322 VSS.n176 VSS.n81 4.5005
R3323 VSS.n212 VSS.n81 4.5005
R3324 VSS.n175 VSS.n81 4.5005
R3325 VSS.n213 VSS.n81 4.5005
R3326 VSS.n174 VSS.n81 4.5005
R3327 VSS.n214 VSS.n81 4.5005
R3328 VSS.n173 VSS.n81 4.5005
R3329 VSS.n215 VSS.n81 4.5005
R3330 VSS.n172 VSS.n81 4.5005
R3331 VSS.n216 VSS.n81 4.5005
R3332 VSS.n171 VSS.n81 4.5005
R3333 VSS.n217 VSS.n81 4.5005
R3334 VSS.n170 VSS.n81 4.5005
R3335 VSS.n218 VSS.n81 4.5005
R3336 VSS.n169 VSS.n81 4.5005
R3337 VSS.n219 VSS.n81 4.5005
R3338 VSS.n168 VSS.n81 4.5005
R3339 VSS.n220 VSS.n81 4.5005
R3340 VSS.n167 VSS.n81 4.5005
R3341 VSS.n221 VSS.n81 4.5005
R3342 VSS.n166 VSS.n81 4.5005
R3343 VSS.n222 VSS.n81 4.5005
R3344 VSS.n165 VSS.n81 4.5005
R3345 VSS.n223 VSS.n81 4.5005
R3346 VSS.n164 VSS.n81 4.5005
R3347 VSS.n224 VSS.n81 4.5005
R3348 VSS.n163 VSS.n81 4.5005
R3349 VSS.n225 VSS.n81 4.5005
R3350 VSS.n162 VSS.n81 4.5005
R3351 VSS.n226 VSS.n81 4.5005
R3352 VSS.n161 VSS.n81 4.5005
R3353 VSS.n227 VSS.n81 4.5005
R3354 VSS.n160 VSS.n81 4.5005
R3355 VSS.n228 VSS.n81 4.5005
R3356 VSS.n159 VSS.n81 4.5005
R3357 VSS.n229 VSS.n81 4.5005
R3358 VSS.n158 VSS.n81 4.5005
R3359 VSS.n230 VSS.n81 4.5005
R3360 VSS.n157 VSS.n81 4.5005
R3361 VSS.n231 VSS.n81 4.5005
R3362 VSS.n156 VSS.n81 4.5005
R3363 VSS.n232 VSS.n81 4.5005
R3364 VSS.n155 VSS.n81 4.5005
R3365 VSS.n233 VSS.n81 4.5005
R3366 VSS.n154 VSS.n81 4.5005
R3367 VSS.n234 VSS.n81 4.5005
R3368 VSS.n153 VSS.n81 4.5005
R3369 VSS.n235 VSS.n81 4.5005
R3370 VSS.n4506 VSS.n81 4.5005
R3371 VSS.n236 VSS.n81 4.5005
R3372 VSS.n152 VSS.n81 4.5005
R3373 VSS.n237 VSS.n81 4.5005
R3374 VSS.n151 VSS.n81 4.5005
R3375 VSS.n238 VSS.n81 4.5005
R3376 VSS.n150 VSS.n81 4.5005
R3377 VSS.n239 VSS.n81 4.5005
R3378 VSS.n149 VSS.n81 4.5005
R3379 VSS.n240 VSS.n81 4.5005
R3380 VSS.n148 VSS.n81 4.5005
R3381 VSS.n241 VSS.n81 4.5005
R3382 VSS.n147 VSS.n81 4.5005
R3383 VSS.n242 VSS.n81 4.5005
R3384 VSS.n146 VSS.n81 4.5005
R3385 VSS.n243 VSS.n81 4.5005
R3386 VSS.n145 VSS.n81 4.5005
R3387 VSS.n244 VSS.n81 4.5005
R3388 VSS.n144 VSS.n81 4.5005
R3389 VSS.n245 VSS.n81 4.5005
R3390 VSS.n143 VSS.n81 4.5005
R3391 VSS.n246 VSS.n81 4.5005
R3392 VSS.n142 VSS.n81 4.5005
R3393 VSS.n247 VSS.n81 4.5005
R3394 VSS.n141 VSS.n81 4.5005
R3395 VSS.n248 VSS.n81 4.5005
R3396 VSS.n140 VSS.n81 4.5005
R3397 VSS.n249 VSS.n81 4.5005
R3398 VSS.n139 VSS.n81 4.5005
R3399 VSS.n250 VSS.n81 4.5005
R3400 VSS.n138 VSS.n81 4.5005
R3401 VSS.n251 VSS.n81 4.5005
R3402 VSS.n137 VSS.n81 4.5005
R3403 VSS.n252 VSS.n81 4.5005
R3404 VSS.n136 VSS.n81 4.5005
R3405 VSS.n253 VSS.n81 4.5005
R3406 VSS.n135 VSS.n81 4.5005
R3407 VSS.n254 VSS.n81 4.5005
R3408 VSS.n134 VSS.n81 4.5005
R3409 VSS.n255 VSS.n81 4.5005
R3410 VSS.n133 VSS.n81 4.5005
R3411 VSS.n256 VSS.n81 4.5005
R3412 VSS.n132 VSS.n81 4.5005
R3413 VSS.n4502 VSS.n81 4.5005
R3414 VSS.n4504 VSS.n81 4.5005
R3415 VSS.n193 VSS.n55 4.5005
R3416 VSS.n195 VSS.n55 4.5005
R3417 VSS.n192 VSS.n55 4.5005
R3418 VSS.n196 VSS.n55 4.5005
R3419 VSS.n191 VSS.n55 4.5005
R3420 VSS.n197 VSS.n55 4.5005
R3421 VSS.n190 VSS.n55 4.5005
R3422 VSS.n198 VSS.n55 4.5005
R3423 VSS.n189 VSS.n55 4.5005
R3424 VSS.n199 VSS.n55 4.5005
R3425 VSS.n188 VSS.n55 4.5005
R3426 VSS.n200 VSS.n55 4.5005
R3427 VSS.n187 VSS.n55 4.5005
R3428 VSS.n201 VSS.n55 4.5005
R3429 VSS.n186 VSS.n55 4.5005
R3430 VSS.n202 VSS.n55 4.5005
R3431 VSS.n185 VSS.n55 4.5005
R3432 VSS.n203 VSS.n55 4.5005
R3433 VSS.n184 VSS.n55 4.5005
R3434 VSS.n204 VSS.n55 4.5005
R3435 VSS.n183 VSS.n55 4.5005
R3436 VSS.n205 VSS.n55 4.5005
R3437 VSS.n182 VSS.n55 4.5005
R3438 VSS.n206 VSS.n55 4.5005
R3439 VSS.n181 VSS.n55 4.5005
R3440 VSS.n207 VSS.n55 4.5005
R3441 VSS.n180 VSS.n55 4.5005
R3442 VSS.n208 VSS.n55 4.5005
R3443 VSS.n179 VSS.n55 4.5005
R3444 VSS.n209 VSS.n55 4.5005
R3445 VSS.n178 VSS.n55 4.5005
R3446 VSS.n210 VSS.n55 4.5005
R3447 VSS.n177 VSS.n55 4.5005
R3448 VSS.n211 VSS.n55 4.5005
R3449 VSS.n176 VSS.n55 4.5005
R3450 VSS.n212 VSS.n55 4.5005
R3451 VSS.n175 VSS.n55 4.5005
R3452 VSS.n213 VSS.n55 4.5005
R3453 VSS.n174 VSS.n55 4.5005
R3454 VSS.n214 VSS.n55 4.5005
R3455 VSS.n173 VSS.n55 4.5005
R3456 VSS.n215 VSS.n55 4.5005
R3457 VSS.n172 VSS.n55 4.5005
R3458 VSS.n216 VSS.n55 4.5005
R3459 VSS.n171 VSS.n55 4.5005
R3460 VSS.n217 VSS.n55 4.5005
R3461 VSS.n170 VSS.n55 4.5005
R3462 VSS.n218 VSS.n55 4.5005
R3463 VSS.n169 VSS.n55 4.5005
R3464 VSS.n219 VSS.n55 4.5005
R3465 VSS.n168 VSS.n55 4.5005
R3466 VSS.n220 VSS.n55 4.5005
R3467 VSS.n167 VSS.n55 4.5005
R3468 VSS.n221 VSS.n55 4.5005
R3469 VSS.n166 VSS.n55 4.5005
R3470 VSS.n222 VSS.n55 4.5005
R3471 VSS.n165 VSS.n55 4.5005
R3472 VSS.n223 VSS.n55 4.5005
R3473 VSS.n164 VSS.n55 4.5005
R3474 VSS.n224 VSS.n55 4.5005
R3475 VSS.n163 VSS.n55 4.5005
R3476 VSS.n225 VSS.n55 4.5005
R3477 VSS.n162 VSS.n55 4.5005
R3478 VSS.n226 VSS.n55 4.5005
R3479 VSS.n161 VSS.n55 4.5005
R3480 VSS.n227 VSS.n55 4.5005
R3481 VSS.n160 VSS.n55 4.5005
R3482 VSS.n228 VSS.n55 4.5005
R3483 VSS.n159 VSS.n55 4.5005
R3484 VSS.n229 VSS.n55 4.5005
R3485 VSS.n158 VSS.n55 4.5005
R3486 VSS.n230 VSS.n55 4.5005
R3487 VSS.n157 VSS.n55 4.5005
R3488 VSS.n231 VSS.n55 4.5005
R3489 VSS.n156 VSS.n55 4.5005
R3490 VSS.n232 VSS.n55 4.5005
R3491 VSS.n155 VSS.n55 4.5005
R3492 VSS.n233 VSS.n55 4.5005
R3493 VSS.n154 VSS.n55 4.5005
R3494 VSS.n234 VSS.n55 4.5005
R3495 VSS.n153 VSS.n55 4.5005
R3496 VSS.n235 VSS.n55 4.5005
R3497 VSS.n4506 VSS.n55 4.5005
R3498 VSS.n236 VSS.n55 4.5005
R3499 VSS.n152 VSS.n55 4.5005
R3500 VSS.n237 VSS.n55 4.5005
R3501 VSS.n151 VSS.n55 4.5005
R3502 VSS.n238 VSS.n55 4.5005
R3503 VSS.n150 VSS.n55 4.5005
R3504 VSS.n239 VSS.n55 4.5005
R3505 VSS.n149 VSS.n55 4.5005
R3506 VSS.n240 VSS.n55 4.5005
R3507 VSS.n148 VSS.n55 4.5005
R3508 VSS.n241 VSS.n55 4.5005
R3509 VSS.n147 VSS.n55 4.5005
R3510 VSS.n242 VSS.n55 4.5005
R3511 VSS.n146 VSS.n55 4.5005
R3512 VSS.n243 VSS.n55 4.5005
R3513 VSS.n145 VSS.n55 4.5005
R3514 VSS.n244 VSS.n55 4.5005
R3515 VSS.n144 VSS.n55 4.5005
R3516 VSS.n245 VSS.n55 4.5005
R3517 VSS.n143 VSS.n55 4.5005
R3518 VSS.n246 VSS.n55 4.5005
R3519 VSS.n142 VSS.n55 4.5005
R3520 VSS.n247 VSS.n55 4.5005
R3521 VSS.n141 VSS.n55 4.5005
R3522 VSS.n248 VSS.n55 4.5005
R3523 VSS.n140 VSS.n55 4.5005
R3524 VSS.n249 VSS.n55 4.5005
R3525 VSS.n139 VSS.n55 4.5005
R3526 VSS.n250 VSS.n55 4.5005
R3527 VSS.n138 VSS.n55 4.5005
R3528 VSS.n251 VSS.n55 4.5005
R3529 VSS.n137 VSS.n55 4.5005
R3530 VSS.n252 VSS.n55 4.5005
R3531 VSS.n136 VSS.n55 4.5005
R3532 VSS.n253 VSS.n55 4.5005
R3533 VSS.n135 VSS.n55 4.5005
R3534 VSS.n254 VSS.n55 4.5005
R3535 VSS.n134 VSS.n55 4.5005
R3536 VSS.n255 VSS.n55 4.5005
R3537 VSS.n133 VSS.n55 4.5005
R3538 VSS.n256 VSS.n55 4.5005
R3539 VSS.n132 VSS.n55 4.5005
R3540 VSS.n4502 VSS.n55 4.5005
R3541 VSS.n4504 VSS.n55 4.5005
R3542 VSS.n193 VSS.n82 4.5005
R3543 VSS.n195 VSS.n82 4.5005
R3544 VSS.n192 VSS.n82 4.5005
R3545 VSS.n196 VSS.n82 4.5005
R3546 VSS.n191 VSS.n82 4.5005
R3547 VSS.n197 VSS.n82 4.5005
R3548 VSS.n190 VSS.n82 4.5005
R3549 VSS.n198 VSS.n82 4.5005
R3550 VSS.n189 VSS.n82 4.5005
R3551 VSS.n199 VSS.n82 4.5005
R3552 VSS.n188 VSS.n82 4.5005
R3553 VSS.n200 VSS.n82 4.5005
R3554 VSS.n187 VSS.n82 4.5005
R3555 VSS.n201 VSS.n82 4.5005
R3556 VSS.n186 VSS.n82 4.5005
R3557 VSS.n202 VSS.n82 4.5005
R3558 VSS.n185 VSS.n82 4.5005
R3559 VSS.n203 VSS.n82 4.5005
R3560 VSS.n184 VSS.n82 4.5005
R3561 VSS.n204 VSS.n82 4.5005
R3562 VSS.n183 VSS.n82 4.5005
R3563 VSS.n205 VSS.n82 4.5005
R3564 VSS.n182 VSS.n82 4.5005
R3565 VSS.n206 VSS.n82 4.5005
R3566 VSS.n181 VSS.n82 4.5005
R3567 VSS.n207 VSS.n82 4.5005
R3568 VSS.n180 VSS.n82 4.5005
R3569 VSS.n208 VSS.n82 4.5005
R3570 VSS.n179 VSS.n82 4.5005
R3571 VSS.n209 VSS.n82 4.5005
R3572 VSS.n178 VSS.n82 4.5005
R3573 VSS.n210 VSS.n82 4.5005
R3574 VSS.n177 VSS.n82 4.5005
R3575 VSS.n211 VSS.n82 4.5005
R3576 VSS.n176 VSS.n82 4.5005
R3577 VSS.n212 VSS.n82 4.5005
R3578 VSS.n175 VSS.n82 4.5005
R3579 VSS.n213 VSS.n82 4.5005
R3580 VSS.n174 VSS.n82 4.5005
R3581 VSS.n214 VSS.n82 4.5005
R3582 VSS.n173 VSS.n82 4.5005
R3583 VSS.n215 VSS.n82 4.5005
R3584 VSS.n172 VSS.n82 4.5005
R3585 VSS.n216 VSS.n82 4.5005
R3586 VSS.n171 VSS.n82 4.5005
R3587 VSS.n217 VSS.n82 4.5005
R3588 VSS.n170 VSS.n82 4.5005
R3589 VSS.n218 VSS.n82 4.5005
R3590 VSS.n169 VSS.n82 4.5005
R3591 VSS.n219 VSS.n82 4.5005
R3592 VSS.n168 VSS.n82 4.5005
R3593 VSS.n220 VSS.n82 4.5005
R3594 VSS.n167 VSS.n82 4.5005
R3595 VSS.n221 VSS.n82 4.5005
R3596 VSS.n166 VSS.n82 4.5005
R3597 VSS.n222 VSS.n82 4.5005
R3598 VSS.n165 VSS.n82 4.5005
R3599 VSS.n223 VSS.n82 4.5005
R3600 VSS.n164 VSS.n82 4.5005
R3601 VSS.n224 VSS.n82 4.5005
R3602 VSS.n163 VSS.n82 4.5005
R3603 VSS.n225 VSS.n82 4.5005
R3604 VSS.n162 VSS.n82 4.5005
R3605 VSS.n226 VSS.n82 4.5005
R3606 VSS.n161 VSS.n82 4.5005
R3607 VSS.n227 VSS.n82 4.5005
R3608 VSS.n160 VSS.n82 4.5005
R3609 VSS.n228 VSS.n82 4.5005
R3610 VSS.n159 VSS.n82 4.5005
R3611 VSS.n229 VSS.n82 4.5005
R3612 VSS.n158 VSS.n82 4.5005
R3613 VSS.n230 VSS.n82 4.5005
R3614 VSS.n157 VSS.n82 4.5005
R3615 VSS.n231 VSS.n82 4.5005
R3616 VSS.n156 VSS.n82 4.5005
R3617 VSS.n232 VSS.n82 4.5005
R3618 VSS.n155 VSS.n82 4.5005
R3619 VSS.n233 VSS.n82 4.5005
R3620 VSS.n154 VSS.n82 4.5005
R3621 VSS.n234 VSS.n82 4.5005
R3622 VSS.n153 VSS.n82 4.5005
R3623 VSS.n235 VSS.n82 4.5005
R3624 VSS.n4506 VSS.n82 4.5005
R3625 VSS.n236 VSS.n82 4.5005
R3626 VSS.n152 VSS.n82 4.5005
R3627 VSS.n237 VSS.n82 4.5005
R3628 VSS.n151 VSS.n82 4.5005
R3629 VSS.n238 VSS.n82 4.5005
R3630 VSS.n150 VSS.n82 4.5005
R3631 VSS.n239 VSS.n82 4.5005
R3632 VSS.n149 VSS.n82 4.5005
R3633 VSS.n240 VSS.n82 4.5005
R3634 VSS.n148 VSS.n82 4.5005
R3635 VSS.n241 VSS.n82 4.5005
R3636 VSS.n147 VSS.n82 4.5005
R3637 VSS.n242 VSS.n82 4.5005
R3638 VSS.n146 VSS.n82 4.5005
R3639 VSS.n243 VSS.n82 4.5005
R3640 VSS.n145 VSS.n82 4.5005
R3641 VSS.n244 VSS.n82 4.5005
R3642 VSS.n144 VSS.n82 4.5005
R3643 VSS.n245 VSS.n82 4.5005
R3644 VSS.n143 VSS.n82 4.5005
R3645 VSS.n246 VSS.n82 4.5005
R3646 VSS.n142 VSS.n82 4.5005
R3647 VSS.n247 VSS.n82 4.5005
R3648 VSS.n141 VSS.n82 4.5005
R3649 VSS.n248 VSS.n82 4.5005
R3650 VSS.n140 VSS.n82 4.5005
R3651 VSS.n249 VSS.n82 4.5005
R3652 VSS.n139 VSS.n82 4.5005
R3653 VSS.n250 VSS.n82 4.5005
R3654 VSS.n138 VSS.n82 4.5005
R3655 VSS.n251 VSS.n82 4.5005
R3656 VSS.n137 VSS.n82 4.5005
R3657 VSS.n252 VSS.n82 4.5005
R3658 VSS.n136 VSS.n82 4.5005
R3659 VSS.n253 VSS.n82 4.5005
R3660 VSS.n135 VSS.n82 4.5005
R3661 VSS.n254 VSS.n82 4.5005
R3662 VSS.n134 VSS.n82 4.5005
R3663 VSS.n255 VSS.n82 4.5005
R3664 VSS.n133 VSS.n82 4.5005
R3665 VSS.n256 VSS.n82 4.5005
R3666 VSS.n132 VSS.n82 4.5005
R3667 VSS.n4502 VSS.n82 4.5005
R3668 VSS.n4504 VSS.n82 4.5005
R3669 VSS.n193 VSS.n54 4.5005
R3670 VSS.n195 VSS.n54 4.5005
R3671 VSS.n192 VSS.n54 4.5005
R3672 VSS.n196 VSS.n54 4.5005
R3673 VSS.n191 VSS.n54 4.5005
R3674 VSS.n197 VSS.n54 4.5005
R3675 VSS.n190 VSS.n54 4.5005
R3676 VSS.n198 VSS.n54 4.5005
R3677 VSS.n189 VSS.n54 4.5005
R3678 VSS.n199 VSS.n54 4.5005
R3679 VSS.n188 VSS.n54 4.5005
R3680 VSS.n200 VSS.n54 4.5005
R3681 VSS.n187 VSS.n54 4.5005
R3682 VSS.n201 VSS.n54 4.5005
R3683 VSS.n186 VSS.n54 4.5005
R3684 VSS.n202 VSS.n54 4.5005
R3685 VSS.n185 VSS.n54 4.5005
R3686 VSS.n203 VSS.n54 4.5005
R3687 VSS.n184 VSS.n54 4.5005
R3688 VSS.n204 VSS.n54 4.5005
R3689 VSS.n183 VSS.n54 4.5005
R3690 VSS.n205 VSS.n54 4.5005
R3691 VSS.n182 VSS.n54 4.5005
R3692 VSS.n206 VSS.n54 4.5005
R3693 VSS.n181 VSS.n54 4.5005
R3694 VSS.n207 VSS.n54 4.5005
R3695 VSS.n180 VSS.n54 4.5005
R3696 VSS.n208 VSS.n54 4.5005
R3697 VSS.n179 VSS.n54 4.5005
R3698 VSS.n209 VSS.n54 4.5005
R3699 VSS.n178 VSS.n54 4.5005
R3700 VSS.n210 VSS.n54 4.5005
R3701 VSS.n177 VSS.n54 4.5005
R3702 VSS.n211 VSS.n54 4.5005
R3703 VSS.n176 VSS.n54 4.5005
R3704 VSS.n212 VSS.n54 4.5005
R3705 VSS.n175 VSS.n54 4.5005
R3706 VSS.n213 VSS.n54 4.5005
R3707 VSS.n174 VSS.n54 4.5005
R3708 VSS.n214 VSS.n54 4.5005
R3709 VSS.n173 VSS.n54 4.5005
R3710 VSS.n215 VSS.n54 4.5005
R3711 VSS.n172 VSS.n54 4.5005
R3712 VSS.n216 VSS.n54 4.5005
R3713 VSS.n171 VSS.n54 4.5005
R3714 VSS.n217 VSS.n54 4.5005
R3715 VSS.n170 VSS.n54 4.5005
R3716 VSS.n218 VSS.n54 4.5005
R3717 VSS.n169 VSS.n54 4.5005
R3718 VSS.n219 VSS.n54 4.5005
R3719 VSS.n168 VSS.n54 4.5005
R3720 VSS.n220 VSS.n54 4.5005
R3721 VSS.n167 VSS.n54 4.5005
R3722 VSS.n221 VSS.n54 4.5005
R3723 VSS.n166 VSS.n54 4.5005
R3724 VSS.n222 VSS.n54 4.5005
R3725 VSS.n165 VSS.n54 4.5005
R3726 VSS.n223 VSS.n54 4.5005
R3727 VSS.n164 VSS.n54 4.5005
R3728 VSS.n224 VSS.n54 4.5005
R3729 VSS.n163 VSS.n54 4.5005
R3730 VSS.n225 VSS.n54 4.5005
R3731 VSS.n162 VSS.n54 4.5005
R3732 VSS.n226 VSS.n54 4.5005
R3733 VSS.n161 VSS.n54 4.5005
R3734 VSS.n227 VSS.n54 4.5005
R3735 VSS.n160 VSS.n54 4.5005
R3736 VSS.n228 VSS.n54 4.5005
R3737 VSS.n159 VSS.n54 4.5005
R3738 VSS.n229 VSS.n54 4.5005
R3739 VSS.n158 VSS.n54 4.5005
R3740 VSS.n230 VSS.n54 4.5005
R3741 VSS.n157 VSS.n54 4.5005
R3742 VSS.n231 VSS.n54 4.5005
R3743 VSS.n156 VSS.n54 4.5005
R3744 VSS.n232 VSS.n54 4.5005
R3745 VSS.n155 VSS.n54 4.5005
R3746 VSS.n233 VSS.n54 4.5005
R3747 VSS.n154 VSS.n54 4.5005
R3748 VSS.n234 VSS.n54 4.5005
R3749 VSS.n153 VSS.n54 4.5005
R3750 VSS.n235 VSS.n54 4.5005
R3751 VSS.n4506 VSS.n54 4.5005
R3752 VSS.n236 VSS.n54 4.5005
R3753 VSS.n152 VSS.n54 4.5005
R3754 VSS.n237 VSS.n54 4.5005
R3755 VSS.n151 VSS.n54 4.5005
R3756 VSS.n238 VSS.n54 4.5005
R3757 VSS.n150 VSS.n54 4.5005
R3758 VSS.n239 VSS.n54 4.5005
R3759 VSS.n149 VSS.n54 4.5005
R3760 VSS.n240 VSS.n54 4.5005
R3761 VSS.n148 VSS.n54 4.5005
R3762 VSS.n241 VSS.n54 4.5005
R3763 VSS.n147 VSS.n54 4.5005
R3764 VSS.n242 VSS.n54 4.5005
R3765 VSS.n146 VSS.n54 4.5005
R3766 VSS.n243 VSS.n54 4.5005
R3767 VSS.n145 VSS.n54 4.5005
R3768 VSS.n244 VSS.n54 4.5005
R3769 VSS.n144 VSS.n54 4.5005
R3770 VSS.n245 VSS.n54 4.5005
R3771 VSS.n143 VSS.n54 4.5005
R3772 VSS.n246 VSS.n54 4.5005
R3773 VSS.n142 VSS.n54 4.5005
R3774 VSS.n247 VSS.n54 4.5005
R3775 VSS.n141 VSS.n54 4.5005
R3776 VSS.n248 VSS.n54 4.5005
R3777 VSS.n140 VSS.n54 4.5005
R3778 VSS.n249 VSS.n54 4.5005
R3779 VSS.n139 VSS.n54 4.5005
R3780 VSS.n250 VSS.n54 4.5005
R3781 VSS.n138 VSS.n54 4.5005
R3782 VSS.n251 VSS.n54 4.5005
R3783 VSS.n137 VSS.n54 4.5005
R3784 VSS.n252 VSS.n54 4.5005
R3785 VSS.n136 VSS.n54 4.5005
R3786 VSS.n253 VSS.n54 4.5005
R3787 VSS.n135 VSS.n54 4.5005
R3788 VSS.n254 VSS.n54 4.5005
R3789 VSS.n134 VSS.n54 4.5005
R3790 VSS.n255 VSS.n54 4.5005
R3791 VSS.n133 VSS.n54 4.5005
R3792 VSS.n256 VSS.n54 4.5005
R3793 VSS.n132 VSS.n54 4.5005
R3794 VSS.n4502 VSS.n54 4.5005
R3795 VSS.n4504 VSS.n54 4.5005
R3796 VSS.n193 VSS.n83 4.5005
R3797 VSS.n195 VSS.n83 4.5005
R3798 VSS.n192 VSS.n83 4.5005
R3799 VSS.n196 VSS.n83 4.5005
R3800 VSS.n191 VSS.n83 4.5005
R3801 VSS.n197 VSS.n83 4.5005
R3802 VSS.n190 VSS.n83 4.5005
R3803 VSS.n198 VSS.n83 4.5005
R3804 VSS.n189 VSS.n83 4.5005
R3805 VSS.n199 VSS.n83 4.5005
R3806 VSS.n188 VSS.n83 4.5005
R3807 VSS.n200 VSS.n83 4.5005
R3808 VSS.n187 VSS.n83 4.5005
R3809 VSS.n201 VSS.n83 4.5005
R3810 VSS.n186 VSS.n83 4.5005
R3811 VSS.n202 VSS.n83 4.5005
R3812 VSS.n185 VSS.n83 4.5005
R3813 VSS.n203 VSS.n83 4.5005
R3814 VSS.n184 VSS.n83 4.5005
R3815 VSS.n204 VSS.n83 4.5005
R3816 VSS.n183 VSS.n83 4.5005
R3817 VSS.n205 VSS.n83 4.5005
R3818 VSS.n182 VSS.n83 4.5005
R3819 VSS.n206 VSS.n83 4.5005
R3820 VSS.n181 VSS.n83 4.5005
R3821 VSS.n207 VSS.n83 4.5005
R3822 VSS.n180 VSS.n83 4.5005
R3823 VSS.n208 VSS.n83 4.5005
R3824 VSS.n179 VSS.n83 4.5005
R3825 VSS.n209 VSS.n83 4.5005
R3826 VSS.n178 VSS.n83 4.5005
R3827 VSS.n210 VSS.n83 4.5005
R3828 VSS.n177 VSS.n83 4.5005
R3829 VSS.n211 VSS.n83 4.5005
R3830 VSS.n176 VSS.n83 4.5005
R3831 VSS.n212 VSS.n83 4.5005
R3832 VSS.n175 VSS.n83 4.5005
R3833 VSS.n213 VSS.n83 4.5005
R3834 VSS.n174 VSS.n83 4.5005
R3835 VSS.n214 VSS.n83 4.5005
R3836 VSS.n173 VSS.n83 4.5005
R3837 VSS.n215 VSS.n83 4.5005
R3838 VSS.n172 VSS.n83 4.5005
R3839 VSS.n216 VSS.n83 4.5005
R3840 VSS.n171 VSS.n83 4.5005
R3841 VSS.n217 VSS.n83 4.5005
R3842 VSS.n170 VSS.n83 4.5005
R3843 VSS.n218 VSS.n83 4.5005
R3844 VSS.n169 VSS.n83 4.5005
R3845 VSS.n219 VSS.n83 4.5005
R3846 VSS.n168 VSS.n83 4.5005
R3847 VSS.n220 VSS.n83 4.5005
R3848 VSS.n167 VSS.n83 4.5005
R3849 VSS.n221 VSS.n83 4.5005
R3850 VSS.n166 VSS.n83 4.5005
R3851 VSS.n222 VSS.n83 4.5005
R3852 VSS.n165 VSS.n83 4.5005
R3853 VSS.n223 VSS.n83 4.5005
R3854 VSS.n164 VSS.n83 4.5005
R3855 VSS.n224 VSS.n83 4.5005
R3856 VSS.n163 VSS.n83 4.5005
R3857 VSS.n225 VSS.n83 4.5005
R3858 VSS.n162 VSS.n83 4.5005
R3859 VSS.n226 VSS.n83 4.5005
R3860 VSS.n161 VSS.n83 4.5005
R3861 VSS.n227 VSS.n83 4.5005
R3862 VSS.n160 VSS.n83 4.5005
R3863 VSS.n228 VSS.n83 4.5005
R3864 VSS.n159 VSS.n83 4.5005
R3865 VSS.n229 VSS.n83 4.5005
R3866 VSS.n158 VSS.n83 4.5005
R3867 VSS.n230 VSS.n83 4.5005
R3868 VSS.n157 VSS.n83 4.5005
R3869 VSS.n231 VSS.n83 4.5005
R3870 VSS.n156 VSS.n83 4.5005
R3871 VSS.n232 VSS.n83 4.5005
R3872 VSS.n155 VSS.n83 4.5005
R3873 VSS.n233 VSS.n83 4.5005
R3874 VSS.n154 VSS.n83 4.5005
R3875 VSS.n234 VSS.n83 4.5005
R3876 VSS.n153 VSS.n83 4.5005
R3877 VSS.n235 VSS.n83 4.5005
R3878 VSS.n4506 VSS.n83 4.5005
R3879 VSS.n236 VSS.n83 4.5005
R3880 VSS.n152 VSS.n83 4.5005
R3881 VSS.n237 VSS.n83 4.5005
R3882 VSS.n151 VSS.n83 4.5005
R3883 VSS.n238 VSS.n83 4.5005
R3884 VSS.n150 VSS.n83 4.5005
R3885 VSS.n239 VSS.n83 4.5005
R3886 VSS.n149 VSS.n83 4.5005
R3887 VSS.n240 VSS.n83 4.5005
R3888 VSS.n148 VSS.n83 4.5005
R3889 VSS.n241 VSS.n83 4.5005
R3890 VSS.n147 VSS.n83 4.5005
R3891 VSS.n242 VSS.n83 4.5005
R3892 VSS.n146 VSS.n83 4.5005
R3893 VSS.n243 VSS.n83 4.5005
R3894 VSS.n145 VSS.n83 4.5005
R3895 VSS.n244 VSS.n83 4.5005
R3896 VSS.n144 VSS.n83 4.5005
R3897 VSS.n245 VSS.n83 4.5005
R3898 VSS.n143 VSS.n83 4.5005
R3899 VSS.n246 VSS.n83 4.5005
R3900 VSS.n142 VSS.n83 4.5005
R3901 VSS.n247 VSS.n83 4.5005
R3902 VSS.n141 VSS.n83 4.5005
R3903 VSS.n248 VSS.n83 4.5005
R3904 VSS.n140 VSS.n83 4.5005
R3905 VSS.n249 VSS.n83 4.5005
R3906 VSS.n139 VSS.n83 4.5005
R3907 VSS.n250 VSS.n83 4.5005
R3908 VSS.n138 VSS.n83 4.5005
R3909 VSS.n251 VSS.n83 4.5005
R3910 VSS.n137 VSS.n83 4.5005
R3911 VSS.n252 VSS.n83 4.5005
R3912 VSS.n136 VSS.n83 4.5005
R3913 VSS.n253 VSS.n83 4.5005
R3914 VSS.n135 VSS.n83 4.5005
R3915 VSS.n254 VSS.n83 4.5005
R3916 VSS.n134 VSS.n83 4.5005
R3917 VSS.n255 VSS.n83 4.5005
R3918 VSS.n133 VSS.n83 4.5005
R3919 VSS.n256 VSS.n83 4.5005
R3920 VSS.n132 VSS.n83 4.5005
R3921 VSS.n4502 VSS.n83 4.5005
R3922 VSS.n4504 VSS.n83 4.5005
R3923 VSS.n193 VSS.n53 4.5005
R3924 VSS.n195 VSS.n53 4.5005
R3925 VSS.n192 VSS.n53 4.5005
R3926 VSS.n196 VSS.n53 4.5005
R3927 VSS.n191 VSS.n53 4.5005
R3928 VSS.n197 VSS.n53 4.5005
R3929 VSS.n190 VSS.n53 4.5005
R3930 VSS.n198 VSS.n53 4.5005
R3931 VSS.n189 VSS.n53 4.5005
R3932 VSS.n199 VSS.n53 4.5005
R3933 VSS.n188 VSS.n53 4.5005
R3934 VSS.n200 VSS.n53 4.5005
R3935 VSS.n187 VSS.n53 4.5005
R3936 VSS.n201 VSS.n53 4.5005
R3937 VSS.n186 VSS.n53 4.5005
R3938 VSS.n202 VSS.n53 4.5005
R3939 VSS.n185 VSS.n53 4.5005
R3940 VSS.n203 VSS.n53 4.5005
R3941 VSS.n184 VSS.n53 4.5005
R3942 VSS.n204 VSS.n53 4.5005
R3943 VSS.n183 VSS.n53 4.5005
R3944 VSS.n205 VSS.n53 4.5005
R3945 VSS.n182 VSS.n53 4.5005
R3946 VSS.n206 VSS.n53 4.5005
R3947 VSS.n181 VSS.n53 4.5005
R3948 VSS.n207 VSS.n53 4.5005
R3949 VSS.n180 VSS.n53 4.5005
R3950 VSS.n208 VSS.n53 4.5005
R3951 VSS.n179 VSS.n53 4.5005
R3952 VSS.n209 VSS.n53 4.5005
R3953 VSS.n178 VSS.n53 4.5005
R3954 VSS.n210 VSS.n53 4.5005
R3955 VSS.n177 VSS.n53 4.5005
R3956 VSS.n211 VSS.n53 4.5005
R3957 VSS.n176 VSS.n53 4.5005
R3958 VSS.n212 VSS.n53 4.5005
R3959 VSS.n175 VSS.n53 4.5005
R3960 VSS.n213 VSS.n53 4.5005
R3961 VSS.n174 VSS.n53 4.5005
R3962 VSS.n214 VSS.n53 4.5005
R3963 VSS.n173 VSS.n53 4.5005
R3964 VSS.n215 VSS.n53 4.5005
R3965 VSS.n172 VSS.n53 4.5005
R3966 VSS.n216 VSS.n53 4.5005
R3967 VSS.n171 VSS.n53 4.5005
R3968 VSS.n217 VSS.n53 4.5005
R3969 VSS.n170 VSS.n53 4.5005
R3970 VSS.n218 VSS.n53 4.5005
R3971 VSS.n169 VSS.n53 4.5005
R3972 VSS.n219 VSS.n53 4.5005
R3973 VSS.n168 VSS.n53 4.5005
R3974 VSS.n220 VSS.n53 4.5005
R3975 VSS.n167 VSS.n53 4.5005
R3976 VSS.n221 VSS.n53 4.5005
R3977 VSS.n166 VSS.n53 4.5005
R3978 VSS.n222 VSS.n53 4.5005
R3979 VSS.n165 VSS.n53 4.5005
R3980 VSS.n223 VSS.n53 4.5005
R3981 VSS.n164 VSS.n53 4.5005
R3982 VSS.n224 VSS.n53 4.5005
R3983 VSS.n163 VSS.n53 4.5005
R3984 VSS.n225 VSS.n53 4.5005
R3985 VSS.n162 VSS.n53 4.5005
R3986 VSS.n226 VSS.n53 4.5005
R3987 VSS.n161 VSS.n53 4.5005
R3988 VSS.n227 VSS.n53 4.5005
R3989 VSS.n160 VSS.n53 4.5005
R3990 VSS.n228 VSS.n53 4.5005
R3991 VSS.n159 VSS.n53 4.5005
R3992 VSS.n229 VSS.n53 4.5005
R3993 VSS.n158 VSS.n53 4.5005
R3994 VSS.n230 VSS.n53 4.5005
R3995 VSS.n157 VSS.n53 4.5005
R3996 VSS.n231 VSS.n53 4.5005
R3997 VSS.n156 VSS.n53 4.5005
R3998 VSS.n232 VSS.n53 4.5005
R3999 VSS.n155 VSS.n53 4.5005
R4000 VSS.n233 VSS.n53 4.5005
R4001 VSS.n154 VSS.n53 4.5005
R4002 VSS.n234 VSS.n53 4.5005
R4003 VSS.n153 VSS.n53 4.5005
R4004 VSS.n235 VSS.n53 4.5005
R4005 VSS.n4506 VSS.n53 4.5005
R4006 VSS.n236 VSS.n53 4.5005
R4007 VSS.n152 VSS.n53 4.5005
R4008 VSS.n237 VSS.n53 4.5005
R4009 VSS.n151 VSS.n53 4.5005
R4010 VSS.n238 VSS.n53 4.5005
R4011 VSS.n150 VSS.n53 4.5005
R4012 VSS.n239 VSS.n53 4.5005
R4013 VSS.n149 VSS.n53 4.5005
R4014 VSS.n240 VSS.n53 4.5005
R4015 VSS.n148 VSS.n53 4.5005
R4016 VSS.n241 VSS.n53 4.5005
R4017 VSS.n147 VSS.n53 4.5005
R4018 VSS.n242 VSS.n53 4.5005
R4019 VSS.n146 VSS.n53 4.5005
R4020 VSS.n243 VSS.n53 4.5005
R4021 VSS.n145 VSS.n53 4.5005
R4022 VSS.n244 VSS.n53 4.5005
R4023 VSS.n144 VSS.n53 4.5005
R4024 VSS.n245 VSS.n53 4.5005
R4025 VSS.n143 VSS.n53 4.5005
R4026 VSS.n246 VSS.n53 4.5005
R4027 VSS.n142 VSS.n53 4.5005
R4028 VSS.n247 VSS.n53 4.5005
R4029 VSS.n141 VSS.n53 4.5005
R4030 VSS.n248 VSS.n53 4.5005
R4031 VSS.n140 VSS.n53 4.5005
R4032 VSS.n249 VSS.n53 4.5005
R4033 VSS.n139 VSS.n53 4.5005
R4034 VSS.n250 VSS.n53 4.5005
R4035 VSS.n138 VSS.n53 4.5005
R4036 VSS.n251 VSS.n53 4.5005
R4037 VSS.n137 VSS.n53 4.5005
R4038 VSS.n252 VSS.n53 4.5005
R4039 VSS.n136 VSS.n53 4.5005
R4040 VSS.n253 VSS.n53 4.5005
R4041 VSS.n135 VSS.n53 4.5005
R4042 VSS.n254 VSS.n53 4.5005
R4043 VSS.n134 VSS.n53 4.5005
R4044 VSS.n255 VSS.n53 4.5005
R4045 VSS.n133 VSS.n53 4.5005
R4046 VSS.n256 VSS.n53 4.5005
R4047 VSS.n132 VSS.n53 4.5005
R4048 VSS.n4502 VSS.n53 4.5005
R4049 VSS.n4504 VSS.n53 4.5005
R4050 VSS.n193 VSS.n84 4.5005
R4051 VSS.n195 VSS.n84 4.5005
R4052 VSS.n192 VSS.n84 4.5005
R4053 VSS.n196 VSS.n84 4.5005
R4054 VSS.n191 VSS.n84 4.5005
R4055 VSS.n197 VSS.n84 4.5005
R4056 VSS.n190 VSS.n84 4.5005
R4057 VSS.n198 VSS.n84 4.5005
R4058 VSS.n189 VSS.n84 4.5005
R4059 VSS.n199 VSS.n84 4.5005
R4060 VSS.n188 VSS.n84 4.5005
R4061 VSS.n200 VSS.n84 4.5005
R4062 VSS.n187 VSS.n84 4.5005
R4063 VSS.n201 VSS.n84 4.5005
R4064 VSS.n186 VSS.n84 4.5005
R4065 VSS.n202 VSS.n84 4.5005
R4066 VSS.n185 VSS.n84 4.5005
R4067 VSS.n203 VSS.n84 4.5005
R4068 VSS.n184 VSS.n84 4.5005
R4069 VSS.n204 VSS.n84 4.5005
R4070 VSS.n183 VSS.n84 4.5005
R4071 VSS.n205 VSS.n84 4.5005
R4072 VSS.n182 VSS.n84 4.5005
R4073 VSS.n206 VSS.n84 4.5005
R4074 VSS.n181 VSS.n84 4.5005
R4075 VSS.n207 VSS.n84 4.5005
R4076 VSS.n180 VSS.n84 4.5005
R4077 VSS.n208 VSS.n84 4.5005
R4078 VSS.n179 VSS.n84 4.5005
R4079 VSS.n209 VSS.n84 4.5005
R4080 VSS.n178 VSS.n84 4.5005
R4081 VSS.n210 VSS.n84 4.5005
R4082 VSS.n177 VSS.n84 4.5005
R4083 VSS.n211 VSS.n84 4.5005
R4084 VSS.n176 VSS.n84 4.5005
R4085 VSS.n212 VSS.n84 4.5005
R4086 VSS.n175 VSS.n84 4.5005
R4087 VSS.n213 VSS.n84 4.5005
R4088 VSS.n174 VSS.n84 4.5005
R4089 VSS.n214 VSS.n84 4.5005
R4090 VSS.n173 VSS.n84 4.5005
R4091 VSS.n215 VSS.n84 4.5005
R4092 VSS.n172 VSS.n84 4.5005
R4093 VSS.n216 VSS.n84 4.5005
R4094 VSS.n171 VSS.n84 4.5005
R4095 VSS.n217 VSS.n84 4.5005
R4096 VSS.n170 VSS.n84 4.5005
R4097 VSS.n218 VSS.n84 4.5005
R4098 VSS.n169 VSS.n84 4.5005
R4099 VSS.n219 VSS.n84 4.5005
R4100 VSS.n168 VSS.n84 4.5005
R4101 VSS.n220 VSS.n84 4.5005
R4102 VSS.n167 VSS.n84 4.5005
R4103 VSS.n221 VSS.n84 4.5005
R4104 VSS.n166 VSS.n84 4.5005
R4105 VSS.n222 VSS.n84 4.5005
R4106 VSS.n165 VSS.n84 4.5005
R4107 VSS.n223 VSS.n84 4.5005
R4108 VSS.n164 VSS.n84 4.5005
R4109 VSS.n224 VSS.n84 4.5005
R4110 VSS.n163 VSS.n84 4.5005
R4111 VSS.n225 VSS.n84 4.5005
R4112 VSS.n162 VSS.n84 4.5005
R4113 VSS.n226 VSS.n84 4.5005
R4114 VSS.n161 VSS.n84 4.5005
R4115 VSS.n227 VSS.n84 4.5005
R4116 VSS.n160 VSS.n84 4.5005
R4117 VSS.n228 VSS.n84 4.5005
R4118 VSS.n159 VSS.n84 4.5005
R4119 VSS.n229 VSS.n84 4.5005
R4120 VSS.n158 VSS.n84 4.5005
R4121 VSS.n230 VSS.n84 4.5005
R4122 VSS.n157 VSS.n84 4.5005
R4123 VSS.n231 VSS.n84 4.5005
R4124 VSS.n156 VSS.n84 4.5005
R4125 VSS.n232 VSS.n84 4.5005
R4126 VSS.n155 VSS.n84 4.5005
R4127 VSS.n233 VSS.n84 4.5005
R4128 VSS.n154 VSS.n84 4.5005
R4129 VSS.n234 VSS.n84 4.5005
R4130 VSS.n153 VSS.n84 4.5005
R4131 VSS.n235 VSS.n84 4.5005
R4132 VSS.n4506 VSS.n84 4.5005
R4133 VSS.n236 VSS.n84 4.5005
R4134 VSS.n152 VSS.n84 4.5005
R4135 VSS.n237 VSS.n84 4.5005
R4136 VSS.n151 VSS.n84 4.5005
R4137 VSS.n238 VSS.n84 4.5005
R4138 VSS.n150 VSS.n84 4.5005
R4139 VSS.n239 VSS.n84 4.5005
R4140 VSS.n149 VSS.n84 4.5005
R4141 VSS.n240 VSS.n84 4.5005
R4142 VSS.n148 VSS.n84 4.5005
R4143 VSS.n241 VSS.n84 4.5005
R4144 VSS.n147 VSS.n84 4.5005
R4145 VSS.n242 VSS.n84 4.5005
R4146 VSS.n146 VSS.n84 4.5005
R4147 VSS.n243 VSS.n84 4.5005
R4148 VSS.n145 VSS.n84 4.5005
R4149 VSS.n244 VSS.n84 4.5005
R4150 VSS.n144 VSS.n84 4.5005
R4151 VSS.n245 VSS.n84 4.5005
R4152 VSS.n143 VSS.n84 4.5005
R4153 VSS.n246 VSS.n84 4.5005
R4154 VSS.n142 VSS.n84 4.5005
R4155 VSS.n247 VSS.n84 4.5005
R4156 VSS.n141 VSS.n84 4.5005
R4157 VSS.n248 VSS.n84 4.5005
R4158 VSS.n140 VSS.n84 4.5005
R4159 VSS.n249 VSS.n84 4.5005
R4160 VSS.n139 VSS.n84 4.5005
R4161 VSS.n250 VSS.n84 4.5005
R4162 VSS.n138 VSS.n84 4.5005
R4163 VSS.n251 VSS.n84 4.5005
R4164 VSS.n137 VSS.n84 4.5005
R4165 VSS.n252 VSS.n84 4.5005
R4166 VSS.n136 VSS.n84 4.5005
R4167 VSS.n253 VSS.n84 4.5005
R4168 VSS.n135 VSS.n84 4.5005
R4169 VSS.n254 VSS.n84 4.5005
R4170 VSS.n134 VSS.n84 4.5005
R4171 VSS.n255 VSS.n84 4.5005
R4172 VSS.n133 VSS.n84 4.5005
R4173 VSS.n256 VSS.n84 4.5005
R4174 VSS.n132 VSS.n84 4.5005
R4175 VSS.n4502 VSS.n84 4.5005
R4176 VSS.n4504 VSS.n84 4.5005
R4177 VSS.n193 VSS.n52 4.5005
R4178 VSS.n195 VSS.n52 4.5005
R4179 VSS.n192 VSS.n52 4.5005
R4180 VSS.n196 VSS.n52 4.5005
R4181 VSS.n191 VSS.n52 4.5005
R4182 VSS.n197 VSS.n52 4.5005
R4183 VSS.n190 VSS.n52 4.5005
R4184 VSS.n198 VSS.n52 4.5005
R4185 VSS.n189 VSS.n52 4.5005
R4186 VSS.n199 VSS.n52 4.5005
R4187 VSS.n188 VSS.n52 4.5005
R4188 VSS.n200 VSS.n52 4.5005
R4189 VSS.n187 VSS.n52 4.5005
R4190 VSS.n201 VSS.n52 4.5005
R4191 VSS.n186 VSS.n52 4.5005
R4192 VSS.n202 VSS.n52 4.5005
R4193 VSS.n185 VSS.n52 4.5005
R4194 VSS.n203 VSS.n52 4.5005
R4195 VSS.n184 VSS.n52 4.5005
R4196 VSS.n204 VSS.n52 4.5005
R4197 VSS.n183 VSS.n52 4.5005
R4198 VSS.n205 VSS.n52 4.5005
R4199 VSS.n182 VSS.n52 4.5005
R4200 VSS.n206 VSS.n52 4.5005
R4201 VSS.n181 VSS.n52 4.5005
R4202 VSS.n207 VSS.n52 4.5005
R4203 VSS.n180 VSS.n52 4.5005
R4204 VSS.n208 VSS.n52 4.5005
R4205 VSS.n179 VSS.n52 4.5005
R4206 VSS.n209 VSS.n52 4.5005
R4207 VSS.n178 VSS.n52 4.5005
R4208 VSS.n210 VSS.n52 4.5005
R4209 VSS.n177 VSS.n52 4.5005
R4210 VSS.n211 VSS.n52 4.5005
R4211 VSS.n176 VSS.n52 4.5005
R4212 VSS.n212 VSS.n52 4.5005
R4213 VSS.n175 VSS.n52 4.5005
R4214 VSS.n213 VSS.n52 4.5005
R4215 VSS.n174 VSS.n52 4.5005
R4216 VSS.n214 VSS.n52 4.5005
R4217 VSS.n173 VSS.n52 4.5005
R4218 VSS.n215 VSS.n52 4.5005
R4219 VSS.n172 VSS.n52 4.5005
R4220 VSS.n216 VSS.n52 4.5005
R4221 VSS.n171 VSS.n52 4.5005
R4222 VSS.n217 VSS.n52 4.5005
R4223 VSS.n170 VSS.n52 4.5005
R4224 VSS.n218 VSS.n52 4.5005
R4225 VSS.n169 VSS.n52 4.5005
R4226 VSS.n219 VSS.n52 4.5005
R4227 VSS.n168 VSS.n52 4.5005
R4228 VSS.n220 VSS.n52 4.5005
R4229 VSS.n167 VSS.n52 4.5005
R4230 VSS.n221 VSS.n52 4.5005
R4231 VSS.n166 VSS.n52 4.5005
R4232 VSS.n222 VSS.n52 4.5005
R4233 VSS.n165 VSS.n52 4.5005
R4234 VSS.n223 VSS.n52 4.5005
R4235 VSS.n164 VSS.n52 4.5005
R4236 VSS.n224 VSS.n52 4.5005
R4237 VSS.n163 VSS.n52 4.5005
R4238 VSS.n225 VSS.n52 4.5005
R4239 VSS.n162 VSS.n52 4.5005
R4240 VSS.n226 VSS.n52 4.5005
R4241 VSS.n161 VSS.n52 4.5005
R4242 VSS.n227 VSS.n52 4.5005
R4243 VSS.n160 VSS.n52 4.5005
R4244 VSS.n228 VSS.n52 4.5005
R4245 VSS.n159 VSS.n52 4.5005
R4246 VSS.n229 VSS.n52 4.5005
R4247 VSS.n158 VSS.n52 4.5005
R4248 VSS.n230 VSS.n52 4.5005
R4249 VSS.n157 VSS.n52 4.5005
R4250 VSS.n231 VSS.n52 4.5005
R4251 VSS.n156 VSS.n52 4.5005
R4252 VSS.n232 VSS.n52 4.5005
R4253 VSS.n155 VSS.n52 4.5005
R4254 VSS.n233 VSS.n52 4.5005
R4255 VSS.n154 VSS.n52 4.5005
R4256 VSS.n234 VSS.n52 4.5005
R4257 VSS.n153 VSS.n52 4.5005
R4258 VSS.n235 VSS.n52 4.5005
R4259 VSS.n4506 VSS.n52 4.5005
R4260 VSS.n236 VSS.n52 4.5005
R4261 VSS.n152 VSS.n52 4.5005
R4262 VSS.n237 VSS.n52 4.5005
R4263 VSS.n151 VSS.n52 4.5005
R4264 VSS.n238 VSS.n52 4.5005
R4265 VSS.n150 VSS.n52 4.5005
R4266 VSS.n239 VSS.n52 4.5005
R4267 VSS.n149 VSS.n52 4.5005
R4268 VSS.n240 VSS.n52 4.5005
R4269 VSS.n148 VSS.n52 4.5005
R4270 VSS.n241 VSS.n52 4.5005
R4271 VSS.n147 VSS.n52 4.5005
R4272 VSS.n242 VSS.n52 4.5005
R4273 VSS.n146 VSS.n52 4.5005
R4274 VSS.n243 VSS.n52 4.5005
R4275 VSS.n145 VSS.n52 4.5005
R4276 VSS.n244 VSS.n52 4.5005
R4277 VSS.n144 VSS.n52 4.5005
R4278 VSS.n245 VSS.n52 4.5005
R4279 VSS.n143 VSS.n52 4.5005
R4280 VSS.n246 VSS.n52 4.5005
R4281 VSS.n142 VSS.n52 4.5005
R4282 VSS.n247 VSS.n52 4.5005
R4283 VSS.n141 VSS.n52 4.5005
R4284 VSS.n248 VSS.n52 4.5005
R4285 VSS.n140 VSS.n52 4.5005
R4286 VSS.n249 VSS.n52 4.5005
R4287 VSS.n139 VSS.n52 4.5005
R4288 VSS.n250 VSS.n52 4.5005
R4289 VSS.n138 VSS.n52 4.5005
R4290 VSS.n251 VSS.n52 4.5005
R4291 VSS.n137 VSS.n52 4.5005
R4292 VSS.n252 VSS.n52 4.5005
R4293 VSS.n136 VSS.n52 4.5005
R4294 VSS.n253 VSS.n52 4.5005
R4295 VSS.n135 VSS.n52 4.5005
R4296 VSS.n254 VSS.n52 4.5005
R4297 VSS.n134 VSS.n52 4.5005
R4298 VSS.n255 VSS.n52 4.5005
R4299 VSS.n133 VSS.n52 4.5005
R4300 VSS.n256 VSS.n52 4.5005
R4301 VSS.n132 VSS.n52 4.5005
R4302 VSS.n4502 VSS.n52 4.5005
R4303 VSS.n4504 VSS.n52 4.5005
R4304 VSS.n193 VSS.n85 4.5005
R4305 VSS.n195 VSS.n85 4.5005
R4306 VSS.n192 VSS.n85 4.5005
R4307 VSS.n196 VSS.n85 4.5005
R4308 VSS.n191 VSS.n85 4.5005
R4309 VSS.n197 VSS.n85 4.5005
R4310 VSS.n190 VSS.n85 4.5005
R4311 VSS.n198 VSS.n85 4.5005
R4312 VSS.n189 VSS.n85 4.5005
R4313 VSS.n199 VSS.n85 4.5005
R4314 VSS.n188 VSS.n85 4.5005
R4315 VSS.n200 VSS.n85 4.5005
R4316 VSS.n187 VSS.n85 4.5005
R4317 VSS.n201 VSS.n85 4.5005
R4318 VSS.n186 VSS.n85 4.5005
R4319 VSS.n202 VSS.n85 4.5005
R4320 VSS.n185 VSS.n85 4.5005
R4321 VSS.n203 VSS.n85 4.5005
R4322 VSS.n184 VSS.n85 4.5005
R4323 VSS.n204 VSS.n85 4.5005
R4324 VSS.n183 VSS.n85 4.5005
R4325 VSS.n205 VSS.n85 4.5005
R4326 VSS.n182 VSS.n85 4.5005
R4327 VSS.n206 VSS.n85 4.5005
R4328 VSS.n181 VSS.n85 4.5005
R4329 VSS.n207 VSS.n85 4.5005
R4330 VSS.n180 VSS.n85 4.5005
R4331 VSS.n208 VSS.n85 4.5005
R4332 VSS.n179 VSS.n85 4.5005
R4333 VSS.n209 VSS.n85 4.5005
R4334 VSS.n178 VSS.n85 4.5005
R4335 VSS.n210 VSS.n85 4.5005
R4336 VSS.n177 VSS.n85 4.5005
R4337 VSS.n211 VSS.n85 4.5005
R4338 VSS.n176 VSS.n85 4.5005
R4339 VSS.n212 VSS.n85 4.5005
R4340 VSS.n175 VSS.n85 4.5005
R4341 VSS.n213 VSS.n85 4.5005
R4342 VSS.n174 VSS.n85 4.5005
R4343 VSS.n214 VSS.n85 4.5005
R4344 VSS.n173 VSS.n85 4.5005
R4345 VSS.n215 VSS.n85 4.5005
R4346 VSS.n172 VSS.n85 4.5005
R4347 VSS.n216 VSS.n85 4.5005
R4348 VSS.n171 VSS.n85 4.5005
R4349 VSS.n217 VSS.n85 4.5005
R4350 VSS.n170 VSS.n85 4.5005
R4351 VSS.n218 VSS.n85 4.5005
R4352 VSS.n169 VSS.n85 4.5005
R4353 VSS.n219 VSS.n85 4.5005
R4354 VSS.n168 VSS.n85 4.5005
R4355 VSS.n220 VSS.n85 4.5005
R4356 VSS.n167 VSS.n85 4.5005
R4357 VSS.n221 VSS.n85 4.5005
R4358 VSS.n166 VSS.n85 4.5005
R4359 VSS.n222 VSS.n85 4.5005
R4360 VSS.n165 VSS.n85 4.5005
R4361 VSS.n223 VSS.n85 4.5005
R4362 VSS.n164 VSS.n85 4.5005
R4363 VSS.n224 VSS.n85 4.5005
R4364 VSS.n163 VSS.n85 4.5005
R4365 VSS.n225 VSS.n85 4.5005
R4366 VSS.n162 VSS.n85 4.5005
R4367 VSS.n226 VSS.n85 4.5005
R4368 VSS.n161 VSS.n85 4.5005
R4369 VSS.n227 VSS.n85 4.5005
R4370 VSS.n160 VSS.n85 4.5005
R4371 VSS.n228 VSS.n85 4.5005
R4372 VSS.n159 VSS.n85 4.5005
R4373 VSS.n229 VSS.n85 4.5005
R4374 VSS.n158 VSS.n85 4.5005
R4375 VSS.n230 VSS.n85 4.5005
R4376 VSS.n157 VSS.n85 4.5005
R4377 VSS.n231 VSS.n85 4.5005
R4378 VSS.n156 VSS.n85 4.5005
R4379 VSS.n232 VSS.n85 4.5005
R4380 VSS.n155 VSS.n85 4.5005
R4381 VSS.n233 VSS.n85 4.5005
R4382 VSS.n154 VSS.n85 4.5005
R4383 VSS.n234 VSS.n85 4.5005
R4384 VSS.n153 VSS.n85 4.5005
R4385 VSS.n235 VSS.n85 4.5005
R4386 VSS.n4506 VSS.n85 4.5005
R4387 VSS.n236 VSS.n85 4.5005
R4388 VSS.n152 VSS.n85 4.5005
R4389 VSS.n237 VSS.n85 4.5005
R4390 VSS.n151 VSS.n85 4.5005
R4391 VSS.n238 VSS.n85 4.5005
R4392 VSS.n150 VSS.n85 4.5005
R4393 VSS.n239 VSS.n85 4.5005
R4394 VSS.n149 VSS.n85 4.5005
R4395 VSS.n240 VSS.n85 4.5005
R4396 VSS.n148 VSS.n85 4.5005
R4397 VSS.n241 VSS.n85 4.5005
R4398 VSS.n147 VSS.n85 4.5005
R4399 VSS.n242 VSS.n85 4.5005
R4400 VSS.n146 VSS.n85 4.5005
R4401 VSS.n243 VSS.n85 4.5005
R4402 VSS.n145 VSS.n85 4.5005
R4403 VSS.n244 VSS.n85 4.5005
R4404 VSS.n144 VSS.n85 4.5005
R4405 VSS.n245 VSS.n85 4.5005
R4406 VSS.n143 VSS.n85 4.5005
R4407 VSS.n246 VSS.n85 4.5005
R4408 VSS.n142 VSS.n85 4.5005
R4409 VSS.n247 VSS.n85 4.5005
R4410 VSS.n141 VSS.n85 4.5005
R4411 VSS.n248 VSS.n85 4.5005
R4412 VSS.n140 VSS.n85 4.5005
R4413 VSS.n249 VSS.n85 4.5005
R4414 VSS.n139 VSS.n85 4.5005
R4415 VSS.n250 VSS.n85 4.5005
R4416 VSS.n138 VSS.n85 4.5005
R4417 VSS.n251 VSS.n85 4.5005
R4418 VSS.n137 VSS.n85 4.5005
R4419 VSS.n252 VSS.n85 4.5005
R4420 VSS.n136 VSS.n85 4.5005
R4421 VSS.n253 VSS.n85 4.5005
R4422 VSS.n135 VSS.n85 4.5005
R4423 VSS.n254 VSS.n85 4.5005
R4424 VSS.n134 VSS.n85 4.5005
R4425 VSS.n255 VSS.n85 4.5005
R4426 VSS.n133 VSS.n85 4.5005
R4427 VSS.n256 VSS.n85 4.5005
R4428 VSS.n132 VSS.n85 4.5005
R4429 VSS.n4502 VSS.n85 4.5005
R4430 VSS.n4504 VSS.n85 4.5005
R4431 VSS.n193 VSS.n51 4.5005
R4432 VSS.n195 VSS.n51 4.5005
R4433 VSS.n192 VSS.n51 4.5005
R4434 VSS.n196 VSS.n51 4.5005
R4435 VSS.n191 VSS.n51 4.5005
R4436 VSS.n197 VSS.n51 4.5005
R4437 VSS.n190 VSS.n51 4.5005
R4438 VSS.n198 VSS.n51 4.5005
R4439 VSS.n189 VSS.n51 4.5005
R4440 VSS.n199 VSS.n51 4.5005
R4441 VSS.n188 VSS.n51 4.5005
R4442 VSS.n200 VSS.n51 4.5005
R4443 VSS.n187 VSS.n51 4.5005
R4444 VSS.n201 VSS.n51 4.5005
R4445 VSS.n186 VSS.n51 4.5005
R4446 VSS.n202 VSS.n51 4.5005
R4447 VSS.n185 VSS.n51 4.5005
R4448 VSS.n203 VSS.n51 4.5005
R4449 VSS.n184 VSS.n51 4.5005
R4450 VSS.n204 VSS.n51 4.5005
R4451 VSS.n183 VSS.n51 4.5005
R4452 VSS.n205 VSS.n51 4.5005
R4453 VSS.n182 VSS.n51 4.5005
R4454 VSS.n206 VSS.n51 4.5005
R4455 VSS.n181 VSS.n51 4.5005
R4456 VSS.n207 VSS.n51 4.5005
R4457 VSS.n180 VSS.n51 4.5005
R4458 VSS.n208 VSS.n51 4.5005
R4459 VSS.n179 VSS.n51 4.5005
R4460 VSS.n209 VSS.n51 4.5005
R4461 VSS.n178 VSS.n51 4.5005
R4462 VSS.n210 VSS.n51 4.5005
R4463 VSS.n177 VSS.n51 4.5005
R4464 VSS.n211 VSS.n51 4.5005
R4465 VSS.n176 VSS.n51 4.5005
R4466 VSS.n212 VSS.n51 4.5005
R4467 VSS.n175 VSS.n51 4.5005
R4468 VSS.n213 VSS.n51 4.5005
R4469 VSS.n174 VSS.n51 4.5005
R4470 VSS.n214 VSS.n51 4.5005
R4471 VSS.n173 VSS.n51 4.5005
R4472 VSS.n215 VSS.n51 4.5005
R4473 VSS.n172 VSS.n51 4.5005
R4474 VSS.n216 VSS.n51 4.5005
R4475 VSS.n171 VSS.n51 4.5005
R4476 VSS.n217 VSS.n51 4.5005
R4477 VSS.n170 VSS.n51 4.5005
R4478 VSS.n218 VSS.n51 4.5005
R4479 VSS.n169 VSS.n51 4.5005
R4480 VSS.n219 VSS.n51 4.5005
R4481 VSS.n168 VSS.n51 4.5005
R4482 VSS.n220 VSS.n51 4.5005
R4483 VSS.n167 VSS.n51 4.5005
R4484 VSS.n221 VSS.n51 4.5005
R4485 VSS.n166 VSS.n51 4.5005
R4486 VSS.n222 VSS.n51 4.5005
R4487 VSS.n165 VSS.n51 4.5005
R4488 VSS.n223 VSS.n51 4.5005
R4489 VSS.n164 VSS.n51 4.5005
R4490 VSS.n224 VSS.n51 4.5005
R4491 VSS.n163 VSS.n51 4.5005
R4492 VSS.n225 VSS.n51 4.5005
R4493 VSS.n162 VSS.n51 4.5005
R4494 VSS.n226 VSS.n51 4.5005
R4495 VSS.n161 VSS.n51 4.5005
R4496 VSS.n227 VSS.n51 4.5005
R4497 VSS.n160 VSS.n51 4.5005
R4498 VSS.n228 VSS.n51 4.5005
R4499 VSS.n159 VSS.n51 4.5005
R4500 VSS.n229 VSS.n51 4.5005
R4501 VSS.n158 VSS.n51 4.5005
R4502 VSS.n230 VSS.n51 4.5005
R4503 VSS.n157 VSS.n51 4.5005
R4504 VSS.n231 VSS.n51 4.5005
R4505 VSS.n156 VSS.n51 4.5005
R4506 VSS.n232 VSS.n51 4.5005
R4507 VSS.n155 VSS.n51 4.5005
R4508 VSS.n233 VSS.n51 4.5005
R4509 VSS.n154 VSS.n51 4.5005
R4510 VSS.n234 VSS.n51 4.5005
R4511 VSS.n153 VSS.n51 4.5005
R4512 VSS.n235 VSS.n51 4.5005
R4513 VSS.n4506 VSS.n51 4.5005
R4514 VSS.n236 VSS.n51 4.5005
R4515 VSS.n152 VSS.n51 4.5005
R4516 VSS.n237 VSS.n51 4.5005
R4517 VSS.n151 VSS.n51 4.5005
R4518 VSS.n238 VSS.n51 4.5005
R4519 VSS.n150 VSS.n51 4.5005
R4520 VSS.n239 VSS.n51 4.5005
R4521 VSS.n149 VSS.n51 4.5005
R4522 VSS.n240 VSS.n51 4.5005
R4523 VSS.n148 VSS.n51 4.5005
R4524 VSS.n241 VSS.n51 4.5005
R4525 VSS.n147 VSS.n51 4.5005
R4526 VSS.n242 VSS.n51 4.5005
R4527 VSS.n146 VSS.n51 4.5005
R4528 VSS.n243 VSS.n51 4.5005
R4529 VSS.n145 VSS.n51 4.5005
R4530 VSS.n244 VSS.n51 4.5005
R4531 VSS.n144 VSS.n51 4.5005
R4532 VSS.n245 VSS.n51 4.5005
R4533 VSS.n143 VSS.n51 4.5005
R4534 VSS.n246 VSS.n51 4.5005
R4535 VSS.n142 VSS.n51 4.5005
R4536 VSS.n247 VSS.n51 4.5005
R4537 VSS.n141 VSS.n51 4.5005
R4538 VSS.n248 VSS.n51 4.5005
R4539 VSS.n140 VSS.n51 4.5005
R4540 VSS.n249 VSS.n51 4.5005
R4541 VSS.n139 VSS.n51 4.5005
R4542 VSS.n250 VSS.n51 4.5005
R4543 VSS.n138 VSS.n51 4.5005
R4544 VSS.n251 VSS.n51 4.5005
R4545 VSS.n137 VSS.n51 4.5005
R4546 VSS.n252 VSS.n51 4.5005
R4547 VSS.n136 VSS.n51 4.5005
R4548 VSS.n253 VSS.n51 4.5005
R4549 VSS.n135 VSS.n51 4.5005
R4550 VSS.n254 VSS.n51 4.5005
R4551 VSS.n134 VSS.n51 4.5005
R4552 VSS.n255 VSS.n51 4.5005
R4553 VSS.n133 VSS.n51 4.5005
R4554 VSS.n256 VSS.n51 4.5005
R4555 VSS.n132 VSS.n51 4.5005
R4556 VSS.n4502 VSS.n51 4.5005
R4557 VSS.n4504 VSS.n51 4.5005
R4558 VSS.n193 VSS.n86 4.5005
R4559 VSS.n195 VSS.n86 4.5005
R4560 VSS.n192 VSS.n86 4.5005
R4561 VSS.n196 VSS.n86 4.5005
R4562 VSS.n191 VSS.n86 4.5005
R4563 VSS.n197 VSS.n86 4.5005
R4564 VSS.n190 VSS.n86 4.5005
R4565 VSS.n198 VSS.n86 4.5005
R4566 VSS.n189 VSS.n86 4.5005
R4567 VSS.n199 VSS.n86 4.5005
R4568 VSS.n188 VSS.n86 4.5005
R4569 VSS.n200 VSS.n86 4.5005
R4570 VSS.n187 VSS.n86 4.5005
R4571 VSS.n201 VSS.n86 4.5005
R4572 VSS.n186 VSS.n86 4.5005
R4573 VSS.n202 VSS.n86 4.5005
R4574 VSS.n185 VSS.n86 4.5005
R4575 VSS.n203 VSS.n86 4.5005
R4576 VSS.n184 VSS.n86 4.5005
R4577 VSS.n204 VSS.n86 4.5005
R4578 VSS.n183 VSS.n86 4.5005
R4579 VSS.n205 VSS.n86 4.5005
R4580 VSS.n182 VSS.n86 4.5005
R4581 VSS.n206 VSS.n86 4.5005
R4582 VSS.n181 VSS.n86 4.5005
R4583 VSS.n207 VSS.n86 4.5005
R4584 VSS.n180 VSS.n86 4.5005
R4585 VSS.n208 VSS.n86 4.5005
R4586 VSS.n179 VSS.n86 4.5005
R4587 VSS.n209 VSS.n86 4.5005
R4588 VSS.n178 VSS.n86 4.5005
R4589 VSS.n210 VSS.n86 4.5005
R4590 VSS.n177 VSS.n86 4.5005
R4591 VSS.n211 VSS.n86 4.5005
R4592 VSS.n176 VSS.n86 4.5005
R4593 VSS.n212 VSS.n86 4.5005
R4594 VSS.n175 VSS.n86 4.5005
R4595 VSS.n213 VSS.n86 4.5005
R4596 VSS.n174 VSS.n86 4.5005
R4597 VSS.n214 VSS.n86 4.5005
R4598 VSS.n173 VSS.n86 4.5005
R4599 VSS.n215 VSS.n86 4.5005
R4600 VSS.n172 VSS.n86 4.5005
R4601 VSS.n216 VSS.n86 4.5005
R4602 VSS.n171 VSS.n86 4.5005
R4603 VSS.n217 VSS.n86 4.5005
R4604 VSS.n170 VSS.n86 4.5005
R4605 VSS.n218 VSS.n86 4.5005
R4606 VSS.n169 VSS.n86 4.5005
R4607 VSS.n219 VSS.n86 4.5005
R4608 VSS.n168 VSS.n86 4.5005
R4609 VSS.n220 VSS.n86 4.5005
R4610 VSS.n167 VSS.n86 4.5005
R4611 VSS.n221 VSS.n86 4.5005
R4612 VSS.n166 VSS.n86 4.5005
R4613 VSS.n222 VSS.n86 4.5005
R4614 VSS.n165 VSS.n86 4.5005
R4615 VSS.n223 VSS.n86 4.5005
R4616 VSS.n164 VSS.n86 4.5005
R4617 VSS.n224 VSS.n86 4.5005
R4618 VSS.n163 VSS.n86 4.5005
R4619 VSS.n225 VSS.n86 4.5005
R4620 VSS.n162 VSS.n86 4.5005
R4621 VSS.n226 VSS.n86 4.5005
R4622 VSS.n161 VSS.n86 4.5005
R4623 VSS.n227 VSS.n86 4.5005
R4624 VSS.n160 VSS.n86 4.5005
R4625 VSS.n228 VSS.n86 4.5005
R4626 VSS.n159 VSS.n86 4.5005
R4627 VSS.n229 VSS.n86 4.5005
R4628 VSS.n158 VSS.n86 4.5005
R4629 VSS.n230 VSS.n86 4.5005
R4630 VSS.n157 VSS.n86 4.5005
R4631 VSS.n231 VSS.n86 4.5005
R4632 VSS.n156 VSS.n86 4.5005
R4633 VSS.n232 VSS.n86 4.5005
R4634 VSS.n155 VSS.n86 4.5005
R4635 VSS.n233 VSS.n86 4.5005
R4636 VSS.n154 VSS.n86 4.5005
R4637 VSS.n234 VSS.n86 4.5005
R4638 VSS.n153 VSS.n86 4.5005
R4639 VSS.n235 VSS.n86 4.5005
R4640 VSS.n4506 VSS.n86 4.5005
R4641 VSS.n236 VSS.n86 4.5005
R4642 VSS.n152 VSS.n86 4.5005
R4643 VSS.n237 VSS.n86 4.5005
R4644 VSS.n151 VSS.n86 4.5005
R4645 VSS.n238 VSS.n86 4.5005
R4646 VSS.n150 VSS.n86 4.5005
R4647 VSS.n239 VSS.n86 4.5005
R4648 VSS.n149 VSS.n86 4.5005
R4649 VSS.n240 VSS.n86 4.5005
R4650 VSS.n148 VSS.n86 4.5005
R4651 VSS.n241 VSS.n86 4.5005
R4652 VSS.n147 VSS.n86 4.5005
R4653 VSS.n242 VSS.n86 4.5005
R4654 VSS.n146 VSS.n86 4.5005
R4655 VSS.n243 VSS.n86 4.5005
R4656 VSS.n145 VSS.n86 4.5005
R4657 VSS.n244 VSS.n86 4.5005
R4658 VSS.n144 VSS.n86 4.5005
R4659 VSS.n245 VSS.n86 4.5005
R4660 VSS.n143 VSS.n86 4.5005
R4661 VSS.n246 VSS.n86 4.5005
R4662 VSS.n142 VSS.n86 4.5005
R4663 VSS.n247 VSS.n86 4.5005
R4664 VSS.n141 VSS.n86 4.5005
R4665 VSS.n248 VSS.n86 4.5005
R4666 VSS.n140 VSS.n86 4.5005
R4667 VSS.n249 VSS.n86 4.5005
R4668 VSS.n139 VSS.n86 4.5005
R4669 VSS.n250 VSS.n86 4.5005
R4670 VSS.n138 VSS.n86 4.5005
R4671 VSS.n251 VSS.n86 4.5005
R4672 VSS.n137 VSS.n86 4.5005
R4673 VSS.n252 VSS.n86 4.5005
R4674 VSS.n136 VSS.n86 4.5005
R4675 VSS.n253 VSS.n86 4.5005
R4676 VSS.n135 VSS.n86 4.5005
R4677 VSS.n254 VSS.n86 4.5005
R4678 VSS.n134 VSS.n86 4.5005
R4679 VSS.n255 VSS.n86 4.5005
R4680 VSS.n133 VSS.n86 4.5005
R4681 VSS.n256 VSS.n86 4.5005
R4682 VSS.n132 VSS.n86 4.5005
R4683 VSS.n4502 VSS.n86 4.5005
R4684 VSS.n4504 VSS.n86 4.5005
R4685 VSS.n193 VSS.n50 4.5005
R4686 VSS.n195 VSS.n50 4.5005
R4687 VSS.n192 VSS.n50 4.5005
R4688 VSS.n196 VSS.n50 4.5005
R4689 VSS.n191 VSS.n50 4.5005
R4690 VSS.n197 VSS.n50 4.5005
R4691 VSS.n190 VSS.n50 4.5005
R4692 VSS.n198 VSS.n50 4.5005
R4693 VSS.n189 VSS.n50 4.5005
R4694 VSS.n199 VSS.n50 4.5005
R4695 VSS.n188 VSS.n50 4.5005
R4696 VSS.n200 VSS.n50 4.5005
R4697 VSS.n187 VSS.n50 4.5005
R4698 VSS.n201 VSS.n50 4.5005
R4699 VSS.n186 VSS.n50 4.5005
R4700 VSS.n202 VSS.n50 4.5005
R4701 VSS.n185 VSS.n50 4.5005
R4702 VSS.n203 VSS.n50 4.5005
R4703 VSS.n184 VSS.n50 4.5005
R4704 VSS.n204 VSS.n50 4.5005
R4705 VSS.n183 VSS.n50 4.5005
R4706 VSS.n205 VSS.n50 4.5005
R4707 VSS.n182 VSS.n50 4.5005
R4708 VSS.n206 VSS.n50 4.5005
R4709 VSS.n181 VSS.n50 4.5005
R4710 VSS.n207 VSS.n50 4.5005
R4711 VSS.n180 VSS.n50 4.5005
R4712 VSS.n208 VSS.n50 4.5005
R4713 VSS.n179 VSS.n50 4.5005
R4714 VSS.n209 VSS.n50 4.5005
R4715 VSS.n178 VSS.n50 4.5005
R4716 VSS.n210 VSS.n50 4.5005
R4717 VSS.n177 VSS.n50 4.5005
R4718 VSS.n211 VSS.n50 4.5005
R4719 VSS.n176 VSS.n50 4.5005
R4720 VSS.n212 VSS.n50 4.5005
R4721 VSS.n175 VSS.n50 4.5005
R4722 VSS.n213 VSS.n50 4.5005
R4723 VSS.n174 VSS.n50 4.5005
R4724 VSS.n214 VSS.n50 4.5005
R4725 VSS.n173 VSS.n50 4.5005
R4726 VSS.n215 VSS.n50 4.5005
R4727 VSS.n172 VSS.n50 4.5005
R4728 VSS.n216 VSS.n50 4.5005
R4729 VSS.n171 VSS.n50 4.5005
R4730 VSS.n217 VSS.n50 4.5005
R4731 VSS.n170 VSS.n50 4.5005
R4732 VSS.n218 VSS.n50 4.5005
R4733 VSS.n169 VSS.n50 4.5005
R4734 VSS.n219 VSS.n50 4.5005
R4735 VSS.n168 VSS.n50 4.5005
R4736 VSS.n220 VSS.n50 4.5005
R4737 VSS.n167 VSS.n50 4.5005
R4738 VSS.n221 VSS.n50 4.5005
R4739 VSS.n166 VSS.n50 4.5005
R4740 VSS.n222 VSS.n50 4.5005
R4741 VSS.n165 VSS.n50 4.5005
R4742 VSS.n223 VSS.n50 4.5005
R4743 VSS.n164 VSS.n50 4.5005
R4744 VSS.n224 VSS.n50 4.5005
R4745 VSS.n163 VSS.n50 4.5005
R4746 VSS.n225 VSS.n50 4.5005
R4747 VSS.n162 VSS.n50 4.5005
R4748 VSS.n226 VSS.n50 4.5005
R4749 VSS.n161 VSS.n50 4.5005
R4750 VSS.n227 VSS.n50 4.5005
R4751 VSS.n160 VSS.n50 4.5005
R4752 VSS.n228 VSS.n50 4.5005
R4753 VSS.n159 VSS.n50 4.5005
R4754 VSS.n229 VSS.n50 4.5005
R4755 VSS.n158 VSS.n50 4.5005
R4756 VSS.n230 VSS.n50 4.5005
R4757 VSS.n157 VSS.n50 4.5005
R4758 VSS.n231 VSS.n50 4.5005
R4759 VSS.n156 VSS.n50 4.5005
R4760 VSS.n232 VSS.n50 4.5005
R4761 VSS.n155 VSS.n50 4.5005
R4762 VSS.n233 VSS.n50 4.5005
R4763 VSS.n154 VSS.n50 4.5005
R4764 VSS.n234 VSS.n50 4.5005
R4765 VSS.n153 VSS.n50 4.5005
R4766 VSS.n235 VSS.n50 4.5005
R4767 VSS.n4506 VSS.n50 4.5005
R4768 VSS.n236 VSS.n50 4.5005
R4769 VSS.n152 VSS.n50 4.5005
R4770 VSS.n237 VSS.n50 4.5005
R4771 VSS.n151 VSS.n50 4.5005
R4772 VSS.n238 VSS.n50 4.5005
R4773 VSS.n150 VSS.n50 4.5005
R4774 VSS.n239 VSS.n50 4.5005
R4775 VSS.n149 VSS.n50 4.5005
R4776 VSS.n240 VSS.n50 4.5005
R4777 VSS.n148 VSS.n50 4.5005
R4778 VSS.n241 VSS.n50 4.5005
R4779 VSS.n147 VSS.n50 4.5005
R4780 VSS.n242 VSS.n50 4.5005
R4781 VSS.n146 VSS.n50 4.5005
R4782 VSS.n243 VSS.n50 4.5005
R4783 VSS.n145 VSS.n50 4.5005
R4784 VSS.n244 VSS.n50 4.5005
R4785 VSS.n144 VSS.n50 4.5005
R4786 VSS.n245 VSS.n50 4.5005
R4787 VSS.n143 VSS.n50 4.5005
R4788 VSS.n246 VSS.n50 4.5005
R4789 VSS.n142 VSS.n50 4.5005
R4790 VSS.n247 VSS.n50 4.5005
R4791 VSS.n141 VSS.n50 4.5005
R4792 VSS.n248 VSS.n50 4.5005
R4793 VSS.n140 VSS.n50 4.5005
R4794 VSS.n249 VSS.n50 4.5005
R4795 VSS.n139 VSS.n50 4.5005
R4796 VSS.n250 VSS.n50 4.5005
R4797 VSS.n138 VSS.n50 4.5005
R4798 VSS.n251 VSS.n50 4.5005
R4799 VSS.n137 VSS.n50 4.5005
R4800 VSS.n252 VSS.n50 4.5005
R4801 VSS.n136 VSS.n50 4.5005
R4802 VSS.n253 VSS.n50 4.5005
R4803 VSS.n135 VSS.n50 4.5005
R4804 VSS.n254 VSS.n50 4.5005
R4805 VSS.n134 VSS.n50 4.5005
R4806 VSS.n255 VSS.n50 4.5005
R4807 VSS.n133 VSS.n50 4.5005
R4808 VSS.n256 VSS.n50 4.5005
R4809 VSS.n132 VSS.n50 4.5005
R4810 VSS.n4502 VSS.n50 4.5005
R4811 VSS.n4504 VSS.n50 4.5005
R4812 VSS.n193 VSS.n87 4.5005
R4813 VSS.n195 VSS.n87 4.5005
R4814 VSS.n192 VSS.n87 4.5005
R4815 VSS.n196 VSS.n87 4.5005
R4816 VSS.n191 VSS.n87 4.5005
R4817 VSS.n197 VSS.n87 4.5005
R4818 VSS.n190 VSS.n87 4.5005
R4819 VSS.n198 VSS.n87 4.5005
R4820 VSS.n189 VSS.n87 4.5005
R4821 VSS.n199 VSS.n87 4.5005
R4822 VSS.n188 VSS.n87 4.5005
R4823 VSS.n200 VSS.n87 4.5005
R4824 VSS.n187 VSS.n87 4.5005
R4825 VSS.n201 VSS.n87 4.5005
R4826 VSS.n186 VSS.n87 4.5005
R4827 VSS.n202 VSS.n87 4.5005
R4828 VSS.n185 VSS.n87 4.5005
R4829 VSS.n203 VSS.n87 4.5005
R4830 VSS.n184 VSS.n87 4.5005
R4831 VSS.n204 VSS.n87 4.5005
R4832 VSS.n183 VSS.n87 4.5005
R4833 VSS.n205 VSS.n87 4.5005
R4834 VSS.n182 VSS.n87 4.5005
R4835 VSS.n206 VSS.n87 4.5005
R4836 VSS.n181 VSS.n87 4.5005
R4837 VSS.n207 VSS.n87 4.5005
R4838 VSS.n180 VSS.n87 4.5005
R4839 VSS.n208 VSS.n87 4.5005
R4840 VSS.n179 VSS.n87 4.5005
R4841 VSS.n209 VSS.n87 4.5005
R4842 VSS.n178 VSS.n87 4.5005
R4843 VSS.n210 VSS.n87 4.5005
R4844 VSS.n177 VSS.n87 4.5005
R4845 VSS.n211 VSS.n87 4.5005
R4846 VSS.n176 VSS.n87 4.5005
R4847 VSS.n212 VSS.n87 4.5005
R4848 VSS.n175 VSS.n87 4.5005
R4849 VSS.n213 VSS.n87 4.5005
R4850 VSS.n174 VSS.n87 4.5005
R4851 VSS.n214 VSS.n87 4.5005
R4852 VSS.n173 VSS.n87 4.5005
R4853 VSS.n215 VSS.n87 4.5005
R4854 VSS.n172 VSS.n87 4.5005
R4855 VSS.n216 VSS.n87 4.5005
R4856 VSS.n171 VSS.n87 4.5005
R4857 VSS.n217 VSS.n87 4.5005
R4858 VSS.n170 VSS.n87 4.5005
R4859 VSS.n218 VSS.n87 4.5005
R4860 VSS.n169 VSS.n87 4.5005
R4861 VSS.n219 VSS.n87 4.5005
R4862 VSS.n168 VSS.n87 4.5005
R4863 VSS.n220 VSS.n87 4.5005
R4864 VSS.n167 VSS.n87 4.5005
R4865 VSS.n221 VSS.n87 4.5005
R4866 VSS.n166 VSS.n87 4.5005
R4867 VSS.n222 VSS.n87 4.5005
R4868 VSS.n165 VSS.n87 4.5005
R4869 VSS.n223 VSS.n87 4.5005
R4870 VSS.n164 VSS.n87 4.5005
R4871 VSS.n224 VSS.n87 4.5005
R4872 VSS.n163 VSS.n87 4.5005
R4873 VSS.n225 VSS.n87 4.5005
R4874 VSS.n162 VSS.n87 4.5005
R4875 VSS.n226 VSS.n87 4.5005
R4876 VSS.n161 VSS.n87 4.5005
R4877 VSS.n227 VSS.n87 4.5005
R4878 VSS.n160 VSS.n87 4.5005
R4879 VSS.n228 VSS.n87 4.5005
R4880 VSS.n159 VSS.n87 4.5005
R4881 VSS.n229 VSS.n87 4.5005
R4882 VSS.n158 VSS.n87 4.5005
R4883 VSS.n230 VSS.n87 4.5005
R4884 VSS.n157 VSS.n87 4.5005
R4885 VSS.n231 VSS.n87 4.5005
R4886 VSS.n156 VSS.n87 4.5005
R4887 VSS.n232 VSS.n87 4.5005
R4888 VSS.n155 VSS.n87 4.5005
R4889 VSS.n233 VSS.n87 4.5005
R4890 VSS.n154 VSS.n87 4.5005
R4891 VSS.n234 VSS.n87 4.5005
R4892 VSS.n153 VSS.n87 4.5005
R4893 VSS.n235 VSS.n87 4.5005
R4894 VSS.n4506 VSS.n87 4.5005
R4895 VSS.n236 VSS.n87 4.5005
R4896 VSS.n152 VSS.n87 4.5005
R4897 VSS.n237 VSS.n87 4.5005
R4898 VSS.n151 VSS.n87 4.5005
R4899 VSS.n238 VSS.n87 4.5005
R4900 VSS.n150 VSS.n87 4.5005
R4901 VSS.n239 VSS.n87 4.5005
R4902 VSS.n149 VSS.n87 4.5005
R4903 VSS.n240 VSS.n87 4.5005
R4904 VSS.n148 VSS.n87 4.5005
R4905 VSS.n241 VSS.n87 4.5005
R4906 VSS.n147 VSS.n87 4.5005
R4907 VSS.n242 VSS.n87 4.5005
R4908 VSS.n146 VSS.n87 4.5005
R4909 VSS.n243 VSS.n87 4.5005
R4910 VSS.n145 VSS.n87 4.5005
R4911 VSS.n244 VSS.n87 4.5005
R4912 VSS.n144 VSS.n87 4.5005
R4913 VSS.n245 VSS.n87 4.5005
R4914 VSS.n143 VSS.n87 4.5005
R4915 VSS.n246 VSS.n87 4.5005
R4916 VSS.n142 VSS.n87 4.5005
R4917 VSS.n247 VSS.n87 4.5005
R4918 VSS.n141 VSS.n87 4.5005
R4919 VSS.n248 VSS.n87 4.5005
R4920 VSS.n140 VSS.n87 4.5005
R4921 VSS.n249 VSS.n87 4.5005
R4922 VSS.n139 VSS.n87 4.5005
R4923 VSS.n250 VSS.n87 4.5005
R4924 VSS.n138 VSS.n87 4.5005
R4925 VSS.n251 VSS.n87 4.5005
R4926 VSS.n137 VSS.n87 4.5005
R4927 VSS.n252 VSS.n87 4.5005
R4928 VSS.n136 VSS.n87 4.5005
R4929 VSS.n253 VSS.n87 4.5005
R4930 VSS.n135 VSS.n87 4.5005
R4931 VSS.n254 VSS.n87 4.5005
R4932 VSS.n134 VSS.n87 4.5005
R4933 VSS.n255 VSS.n87 4.5005
R4934 VSS.n133 VSS.n87 4.5005
R4935 VSS.n256 VSS.n87 4.5005
R4936 VSS.n132 VSS.n87 4.5005
R4937 VSS.n4502 VSS.n87 4.5005
R4938 VSS.n4504 VSS.n87 4.5005
R4939 VSS.n193 VSS.n49 4.5005
R4940 VSS.n195 VSS.n49 4.5005
R4941 VSS.n192 VSS.n49 4.5005
R4942 VSS.n196 VSS.n49 4.5005
R4943 VSS.n191 VSS.n49 4.5005
R4944 VSS.n197 VSS.n49 4.5005
R4945 VSS.n190 VSS.n49 4.5005
R4946 VSS.n198 VSS.n49 4.5005
R4947 VSS.n189 VSS.n49 4.5005
R4948 VSS.n199 VSS.n49 4.5005
R4949 VSS.n188 VSS.n49 4.5005
R4950 VSS.n200 VSS.n49 4.5005
R4951 VSS.n187 VSS.n49 4.5005
R4952 VSS.n201 VSS.n49 4.5005
R4953 VSS.n186 VSS.n49 4.5005
R4954 VSS.n202 VSS.n49 4.5005
R4955 VSS.n185 VSS.n49 4.5005
R4956 VSS.n203 VSS.n49 4.5005
R4957 VSS.n184 VSS.n49 4.5005
R4958 VSS.n204 VSS.n49 4.5005
R4959 VSS.n183 VSS.n49 4.5005
R4960 VSS.n205 VSS.n49 4.5005
R4961 VSS.n182 VSS.n49 4.5005
R4962 VSS.n206 VSS.n49 4.5005
R4963 VSS.n181 VSS.n49 4.5005
R4964 VSS.n207 VSS.n49 4.5005
R4965 VSS.n180 VSS.n49 4.5005
R4966 VSS.n208 VSS.n49 4.5005
R4967 VSS.n179 VSS.n49 4.5005
R4968 VSS.n209 VSS.n49 4.5005
R4969 VSS.n178 VSS.n49 4.5005
R4970 VSS.n210 VSS.n49 4.5005
R4971 VSS.n177 VSS.n49 4.5005
R4972 VSS.n211 VSS.n49 4.5005
R4973 VSS.n176 VSS.n49 4.5005
R4974 VSS.n212 VSS.n49 4.5005
R4975 VSS.n175 VSS.n49 4.5005
R4976 VSS.n213 VSS.n49 4.5005
R4977 VSS.n174 VSS.n49 4.5005
R4978 VSS.n214 VSS.n49 4.5005
R4979 VSS.n173 VSS.n49 4.5005
R4980 VSS.n215 VSS.n49 4.5005
R4981 VSS.n172 VSS.n49 4.5005
R4982 VSS.n216 VSS.n49 4.5005
R4983 VSS.n171 VSS.n49 4.5005
R4984 VSS.n217 VSS.n49 4.5005
R4985 VSS.n170 VSS.n49 4.5005
R4986 VSS.n218 VSS.n49 4.5005
R4987 VSS.n169 VSS.n49 4.5005
R4988 VSS.n219 VSS.n49 4.5005
R4989 VSS.n168 VSS.n49 4.5005
R4990 VSS.n220 VSS.n49 4.5005
R4991 VSS.n167 VSS.n49 4.5005
R4992 VSS.n221 VSS.n49 4.5005
R4993 VSS.n166 VSS.n49 4.5005
R4994 VSS.n222 VSS.n49 4.5005
R4995 VSS.n165 VSS.n49 4.5005
R4996 VSS.n223 VSS.n49 4.5005
R4997 VSS.n164 VSS.n49 4.5005
R4998 VSS.n224 VSS.n49 4.5005
R4999 VSS.n163 VSS.n49 4.5005
R5000 VSS.n225 VSS.n49 4.5005
R5001 VSS.n162 VSS.n49 4.5005
R5002 VSS.n226 VSS.n49 4.5005
R5003 VSS.n161 VSS.n49 4.5005
R5004 VSS.n227 VSS.n49 4.5005
R5005 VSS.n160 VSS.n49 4.5005
R5006 VSS.n228 VSS.n49 4.5005
R5007 VSS.n159 VSS.n49 4.5005
R5008 VSS.n229 VSS.n49 4.5005
R5009 VSS.n158 VSS.n49 4.5005
R5010 VSS.n230 VSS.n49 4.5005
R5011 VSS.n157 VSS.n49 4.5005
R5012 VSS.n231 VSS.n49 4.5005
R5013 VSS.n156 VSS.n49 4.5005
R5014 VSS.n232 VSS.n49 4.5005
R5015 VSS.n155 VSS.n49 4.5005
R5016 VSS.n233 VSS.n49 4.5005
R5017 VSS.n154 VSS.n49 4.5005
R5018 VSS.n234 VSS.n49 4.5005
R5019 VSS.n153 VSS.n49 4.5005
R5020 VSS.n235 VSS.n49 4.5005
R5021 VSS.n4506 VSS.n49 4.5005
R5022 VSS.n236 VSS.n49 4.5005
R5023 VSS.n152 VSS.n49 4.5005
R5024 VSS.n237 VSS.n49 4.5005
R5025 VSS.n151 VSS.n49 4.5005
R5026 VSS.n238 VSS.n49 4.5005
R5027 VSS.n150 VSS.n49 4.5005
R5028 VSS.n239 VSS.n49 4.5005
R5029 VSS.n149 VSS.n49 4.5005
R5030 VSS.n240 VSS.n49 4.5005
R5031 VSS.n148 VSS.n49 4.5005
R5032 VSS.n241 VSS.n49 4.5005
R5033 VSS.n147 VSS.n49 4.5005
R5034 VSS.n242 VSS.n49 4.5005
R5035 VSS.n146 VSS.n49 4.5005
R5036 VSS.n243 VSS.n49 4.5005
R5037 VSS.n145 VSS.n49 4.5005
R5038 VSS.n244 VSS.n49 4.5005
R5039 VSS.n144 VSS.n49 4.5005
R5040 VSS.n245 VSS.n49 4.5005
R5041 VSS.n143 VSS.n49 4.5005
R5042 VSS.n246 VSS.n49 4.5005
R5043 VSS.n142 VSS.n49 4.5005
R5044 VSS.n247 VSS.n49 4.5005
R5045 VSS.n141 VSS.n49 4.5005
R5046 VSS.n248 VSS.n49 4.5005
R5047 VSS.n140 VSS.n49 4.5005
R5048 VSS.n249 VSS.n49 4.5005
R5049 VSS.n139 VSS.n49 4.5005
R5050 VSS.n250 VSS.n49 4.5005
R5051 VSS.n138 VSS.n49 4.5005
R5052 VSS.n251 VSS.n49 4.5005
R5053 VSS.n137 VSS.n49 4.5005
R5054 VSS.n252 VSS.n49 4.5005
R5055 VSS.n136 VSS.n49 4.5005
R5056 VSS.n253 VSS.n49 4.5005
R5057 VSS.n135 VSS.n49 4.5005
R5058 VSS.n254 VSS.n49 4.5005
R5059 VSS.n134 VSS.n49 4.5005
R5060 VSS.n255 VSS.n49 4.5005
R5061 VSS.n133 VSS.n49 4.5005
R5062 VSS.n256 VSS.n49 4.5005
R5063 VSS.n132 VSS.n49 4.5005
R5064 VSS.n4502 VSS.n49 4.5005
R5065 VSS.n4504 VSS.n49 4.5005
R5066 VSS.n193 VSS.n88 4.5005
R5067 VSS.n195 VSS.n88 4.5005
R5068 VSS.n192 VSS.n88 4.5005
R5069 VSS.n196 VSS.n88 4.5005
R5070 VSS.n191 VSS.n88 4.5005
R5071 VSS.n197 VSS.n88 4.5005
R5072 VSS.n190 VSS.n88 4.5005
R5073 VSS.n198 VSS.n88 4.5005
R5074 VSS.n189 VSS.n88 4.5005
R5075 VSS.n199 VSS.n88 4.5005
R5076 VSS.n188 VSS.n88 4.5005
R5077 VSS.n200 VSS.n88 4.5005
R5078 VSS.n187 VSS.n88 4.5005
R5079 VSS.n201 VSS.n88 4.5005
R5080 VSS.n186 VSS.n88 4.5005
R5081 VSS.n202 VSS.n88 4.5005
R5082 VSS.n185 VSS.n88 4.5005
R5083 VSS.n203 VSS.n88 4.5005
R5084 VSS.n184 VSS.n88 4.5005
R5085 VSS.n204 VSS.n88 4.5005
R5086 VSS.n183 VSS.n88 4.5005
R5087 VSS.n205 VSS.n88 4.5005
R5088 VSS.n182 VSS.n88 4.5005
R5089 VSS.n206 VSS.n88 4.5005
R5090 VSS.n181 VSS.n88 4.5005
R5091 VSS.n207 VSS.n88 4.5005
R5092 VSS.n180 VSS.n88 4.5005
R5093 VSS.n208 VSS.n88 4.5005
R5094 VSS.n179 VSS.n88 4.5005
R5095 VSS.n209 VSS.n88 4.5005
R5096 VSS.n178 VSS.n88 4.5005
R5097 VSS.n210 VSS.n88 4.5005
R5098 VSS.n177 VSS.n88 4.5005
R5099 VSS.n211 VSS.n88 4.5005
R5100 VSS.n176 VSS.n88 4.5005
R5101 VSS.n212 VSS.n88 4.5005
R5102 VSS.n175 VSS.n88 4.5005
R5103 VSS.n213 VSS.n88 4.5005
R5104 VSS.n174 VSS.n88 4.5005
R5105 VSS.n214 VSS.n88 4.5005
R5106 VSS.n173 VSS.n88 4.5005
R5107 VSS.n215 VSS.n88 4.5005
R5108 VSS.n172 VSS.n88 4.5005
R5109 VSS.n216 VSS.n88 4.5005
R5110 VSS.n171 VSS.n88 4.5005
R5111 VSS.n217 VSS.n88 4.5005
R5112 VSS.n170 VSS.n88 4.5005
R5113 VSS.n218 VSS.n88 4.5005
R5114 VSS.n169 VSS.n88 4.5005
R5115 VSS.n219 VSS.n88 4.5005
R5116 VSS.n168 VSS.n88 4.5005
R5117 VSS.n220 VSS.n88 4.5005
R5118 VSS.n167 VSS.n88 4.5005
R5119 VSS.n221 VSS.n88 4.5005
R5120 VSS.n166 VSS.n88 4.5005
R5121 VSS.n222 VSS.n88 4.5005
R5122 VSS.n165 VSS.n88 4.5005
R5123 VSS.n223 VSS.n88 4.5005
R5124 VSS.n164 VSS.n88 4.5005
R5125 VSS.n224 VSS.n88 4.5005
R5126 VSS.n163 VSS.n88 4.5005
R5127 VSS.n225 VSS.n88 4.5005
R5128 VSS.n162 VSS.n88 4.5005
R5129 VSS.n226 VSS.n88 4.5005
R5130 VSS.n161 VSS.n88 4.5005
R5131 VSS.n227 VSS.n88 4.5005
R5132 VSS.n160 VSS.n88 4.5005
R5133 VSS.n228 VSS.n88 4.5005
R5134 VSS.n159 VSS.n88 4.5005
R5135 VSS.n229 VSS.n88 4.5005
R5136 VSS.n158 VSS.n88 4.5005
R5137 VSS.n230 VSS.n88 4.5005
R5138 VSS.n157 VSS.n88 4.5005
R5139 VSS.n231 VSS.n88 4.5005
R5140 VSS.n156 VSS.n88 4.5005
R5141 VSS.n232 VSS.n88 4.5005
R5142 VSS.n155 VSS.n88 4.5005
R5143 VSS.n233 VSS.n88 4.5005
R5144 VSS.n154 VSS.n88 4.5005
R5145 VSS.n234 VSS.n88 4.5005
R5146 VSS.n153 VSS.n88 4.5005
R5147 VSS.n235 VSS.n88 4.5005
R5148 VSS.n4506 VSS.n88 4.5005
R5149 VSS.n236 VSS.n88 4.5005
R5150 VSS.n152 VSS.n88 4.5005
R5151 VSS.n237 VSS.n88 4.5005
R5152 VSS.n151 VSS.n88 4.5005
R5153 VSS.n238 VSS.n88 4.5005
R5154 VSS.n150 VSS.n88 4.5005
R5155 VSS.n239 VSS.n88 4.5005
R5156 VSS.n149 VSS.n88 4.5005
R5157 VSS.n240 VSS.n88 4.5005
R5158 VSS.n148 VSS.n88 4.5005
R5159 VSS.n241 VSS.n88 4.5005
R5160 VSS.n147 VSS.n88 4.5005
R5161 VSS.n242 VSS.n88 4.5005
R5162 VSS.n146 VSS.n88 4.5005
R5163 VSS.n243 VSS.n88 4.5005
R5164 VSS.n145 VSS.n88 4.5005
R5165 VSS.n244 VSS.n88 4.5005
R5166 VSS.n144 VSS.n88 4.5005
R5167 VSS.n245 VSS.n88 4.5005
R5168 VSS.n143 VSS.n88 4.5005
R5169 VSS.n246 VSS.n88 4.5005
R5170 VSS.n142 VSS.n88 4.5005
R5171 VSS.n247 VSS.n88 4.5005
R5172 VSS.n141 VSS.n88 4.5005
R5173 VSS.n248 VSS.n88 4.5005
R5174 VSS.n140 VSS.n88 4.5005
R5175 VSS.n249 VSS.n88 4.5005
R5176 VSS.n139 VSS.n88 4.5005
R5177 VSS.n250 VSS.n88 4.5005
R5178 VSS.n138 VSS.n88 4.5005
R5179 VSS.n251 VSS.n88 4.5005
R5180 VSS.n137 VSS.n88 4.5005
R5181 VSS.n252 VSS.n88 4.5005
R5182 VSS.n136 VSS.n88 4.5005
R5183 VSS.n253 VSS.n88 4.5005
R5184 VSS.n135 VSS.n88 4.5005
R5185 VSS.n254 VSS.n88 4.5005
R5186 VSS.n134 VSS.n88 4.5005
R5187 VSS.n255 VSS.n88 4.5005
R5188 VSS.n133 VSS.n88 4.5005
R5189 VSS.n256 VSS.n88 4.5005
R5190 VSS.n132 VSS.n88 4.5005
R5191 VSS.n4502 VSS.n88 4.5005
R5192 VSS.n4504 VSS.n88 4.5005
R5193 VSS.n193 VSS.n48 4.5005
R5194 VSS.n195 VSS.n48 4.5005
R5195 VSS.n192 VSS.n48 4.5005
R5196 VSS.n196 VSS.n48 4.5005
R5197 VSS.n191 VSS.n48 4.5005
R5198 VSS.n197 VSS.n48 4.5005
R5199 VSS.n190 VSS.n48 4.5005
R5200 VSS.n198 VSS.n48 4.5005
R5201 VSS.n189 VSS.n48 4.5005
R5202 VSS.n199 VSS.n48 4.5005
R5203 VSS.n188 VSS.n48 4.5005
R5204 VSS.n200 VSS.n48 4.5005
R5205 VSS.n187 VSS.n48 4.5005
R5206 VSS.n201 VSS.n48 4.5005
R5207 VSS.n186 VSS.n48 4.5005
R5208 VSS.n202 VSS.n48 4.5005
R5209 VSS.n185 VSS.n48 4.5005
R5210 VSS.n203 VSS.n48 4.5005
R5211 VSS.n184 VSS.n48 4.5005
R5212 VSS.n204 VSS.n48 4.5005
R5213 VSS.n183 VSS.n48 4.5005
R5214 VSS.n205 VSS.n48 4.5005
R5215 VSS.n182 VSS.n48 4.5005
R5216 VSS.n206 VSS.n48 4.5005
R5217 VSS.n181 VSS.n48 4.5005
R5218 VSS.n207 VSS.n48 4.5005
R5219 VSS.n180 VSS.n48 4.5005
R5220 VSS.n208 VSS.n48 4.5005
R5221 VSS.n179 VSS.n48 4.5005
R5222 VSS.n209 VSS.n48 4.5005
R5223 VSS.n178 VSS.n48 4.5005
R5224 VSS.n210 VSS.n48 4.5005
R5225 VSS.n177 VSS.n48 4.5005
R5226 VSS.n211 VSS.n48 4.5005
R5227 VSS.n176 VSS.n48 4.5005
R5228 VSS.n212 VSS.n48 4.5005
R5229 VSS.n175 VSS.n48 4.5005
R5230 VSS.n213 VSS.n48 4.5005
R5231 VSS.n174 VSS.n48 4.5005
R5232 VSS.n214 VSS.n48 4.5005
R5233 VSS.n173 VSS.n48 4.5005
R5234 VSS.n215 VSS.n48 4.5005
R5235 VSS.n172 VSS.n48 4.5005
R5236 VSS.n216 VSS.n48 4.5005
R5237 VSS.n171 VSS.n48 4.5005
R5238 VSS.n217 VSS.n48 4.5005
R5239 VSS.n170 VSS.n48 4.5005
R5240 VSS.n218 VSS.n48 4.5005
R5241 VSS.n169 VSS.n48 4.5005
R5242 VSS.n219 VSS.n48 4.5005
R5243 VSS.n168 VSS.n48 4.5005
R5244 VSS.n220 VSS.n48 4.5005
R5245 VSS.n167 VSS.n48 4.5005
R5246 VSS.n221 VSS.n48 4.5005
R5247 VSS.n166 VSS.n48 4.5005
R5248 VSS.n222 VSS.n48 4.5005
R5249 VSS.n165 VSS.n48 4.5005
R5250 VSS.n223 VSS.n48 4.5005
R5251 VSS.n164 VSS.n48 4.5005
R5252 VSS.n224 VSS.n48 4.5005
R5253 VSS.n163 VSS.n48 4.5005
R5254 VSS.n225 VSS.n48 4.5005
R5255 VSS.n162 VSS.n48 4.5005
R5256 VSS.n226 VSS.n48 4.5005
R5257 VSS.n161 VSS.n48 4.5005
R5258 VSS.n227 VSS.n48 4.5005
R5259 VSS.n160 VSS.n48 4.5005
R5260 VSS.n228 VSS.n48 4.5005
R5261 VSS.n159 VSS.n48 4.5005
R5262 VSS.n229 VSS.n48 4.5005
R5263 VSS.n158 VSS.n48 4.5005
R5264 VSS.n230 VSS.n48 4.5005
R5265 VSS.n157 VSS.n48 4.5005
R5266 VSS.n231 VSS.n48 4.5005
R5267 VSS.n156 VSS.n48 4.5005
R5268 VSS.n232 VSS.n48 4.5005
R5269 VSS.n155 VSS.n48 4.5005
R5270 VSS.n233 VSS.n48 4.5005
R5271 VSS.n154 VSS.n48 4.5005
R5272 VSS.n234 VSS.n48 4.5005
R5273 VSS.n153 VSS.n48 4.5005
R5274 VSS.n235 VSS.n48 4.5005
R5275 VSS.n4506 VSS.n48 4.5005
R5276 VSS.n236 VSS.n48 4.5005
R5277 VSS.n152 VSS.n48 4.5005
R5278 VSS.n237 VSS.n48 4.5005
R5279 VSS.n151 VSS.n48 4.5005
R5280 VSS.n238 VSS.n48 4.5005
R5281 VSS.n150 VSS.n48 4.5005
R5282 VSS.n239 VSS.n48 4.5005
R5283 VSS.n149 VSS.n48 4.5005
R5284 VSS.n240 VSS.n48 4.5005
R5285 VSS.n148 VSS.n48 4.5005
R5286 VSS.n241 VSS.n48 4.5005
R5287 VSS.n147 VSS.n48 4.5005
R5288 VSS.n242 VSS.n48 4.5005
R5289 VSS.n146 VSS.n48 4.5005
R5290 VSS.n243 VSS.n48 4.5005
R5291 VSS.n145 VSS.n48 4.5005
R5292 VSS.n244 VSS.n48 4.5005
R5293 VSS.n144 VSS.n48 4.5005
R5294 VSS.n245 VSS.n48 4.5005
R5295 VSS.n143 VSS.n48 4.5005
R5296 VSS.n246 VSS.n48 4.5005
R5297 VSS.n142 VSS.n48 4.5005
R5298 VSS.n247 VSS.n48 4.5005
R5299 VSS.n141 VSS.n48 4.5005
R5300 VSS.n248 VSS.n48 4.5005
R5301 VSS.n140 VSS.n48 4.5005
R5302 VSS.n249 VSS.n48 4.5005
R5303 VSS.n139 VSS.n48 4.5005
R5304 VSS.n250 VSS.n48 4.5005
R5305 VSS.n138 VSS.n48 4.5005
R5306 VSS.n251 VSS.n48 4.5005
R5307 VSS.n137 VSS.n48 4.5005
R5308 VSS.n252 VSS.n48 4.5005
R5309 VSS.n136 VSS.n48 4.5005
R5310 VSS.n253 VSS.n48 4.5005
R5311 VSS.n135 VSS.n48 4.5005
R5312 VSS.n254 VSS.n48 4.5005
R5313 VSS.n134 VSS.n48 4.5005
R5314 VSS.n255 VSS.n48 4.5005
R5315 VSS.n133 VSS.n48 4.5005
R5316 VSS.n256 VSS.n48 4.5005
R5317 VSS.n132 VSS.n48 4.5005
R5318 VSS.n4502 VSS.n48 4.5005
R5319 VSS.n4504 VSS.n48 4.5005
R5320 VSS.n193 VSS.n89 4.5005
R5321 VSS.n195 VSS.n89 4.5005
R5322 VSS.n192 VSS.n89 4.5005
R5323 VSS.n196 VSS.n89 4.5005
R5324 VSS.n191 VSS.n89 4.5005
R5325 VSS.n197 VSS.n89 4.5005
R5326 VSS.n190 VSS.n89 4.5005
R5327 VSS.n198 VSS.n89 4.5005
R5328 VSS.n189 VSS.n89 4.5005
R5329 VSS.n199 VSS.n89 4.5005
R5330 VSS.n188 VSS.n89 4.5005
R5331 VSS.n200 VSS.n89 4.5005
R5332 VSS.n187 VSS.n89 4.5005
R5333 VSS.n201 VSS.n89 4.5005
R5334 VSS.n186 VSS.n89 4.5005
R5335 VSS.n202 VSS.n89 4.5005
R5336 VSS.n185 VSS.n89 4.5005
R5337 VSS.n203 VSS.n89 4.5005
R5338 VSS.n184 VSS.n89 4.5005
R5339 VSS.n204 VSS.n89 4.5005
R5340 VSS.n183 VSS.n89 4.5005
R5341 VSS.n205 VSS.n89 4.5005
R5342 VSS.n182 VSS.n89 4.5005
R5343 VSS.n206 VSS.n89 4.5005
R5344 VSS.n181 VSS.n89 4.5005
R5345 VSS.n207 VSS.n89 4.5005
R5346 VSS.n180 VSS.n89 4.5005
R5347 VSS.n208 VSS.n89 4.5005
R5348 VSS.n179 VSS.n89 4.5005
R5349 VSS.n209 VSS.n89 4.5005
R5350 VSS.n178 VSS.n89 4.5005
R5351 VSS.n210 VSS.n89 4.5005
R5352 VSS.n177 VSS.n89 4.5005
R5353 VSS.n211 VSS.n89 4.5005
R5354 VSS.n176 VSS.n89 4.5005
R5355 VSS.n212 VSS.n89 4.5005
R5356 VSS.n175 VSS.n89 4.5005
R5357 VSS.n213 VSS.n89 4.5005
R5358 VSS.n174 VSS.n89 4.5005
R5359 VSS.n214 VSS.n89 4.5005
R5360 VSS.n173 VSS.n89 4.5005
R5361 VSS.n215 VSS.n89 4.5005
R5362 VSS.n172 VSS.n89 4.5005
R5363 VSS.n216 VSS.n89 4.5005
R5364 VSS.n171 VSS.n89 4.5005
R5365 VSS.n217 VSS.n89 4.5005
R5366 VSS.n170 VSS.n89 4.5005
R5367 VSS.n218 VSS.n89 4.5005
R5368 VSS.n169 VSS.n89 4.5005
R5369 VSS.n219 VSS.n89 4.5005
R5370 VSS.n168 VSS.n89 4.5005
R5371 VSS.n220 VSS.n89 4.5005
R5372 VSS.n167 VSS.n89 4.5005
R5373 VSS.n221 VSS.n89 4.5005
R5374 VSS.n166 VSS.n89 4.5005
R5375 VSS.n222 VSS.n89 4.5005
R5376 VSS.n165 VSS.n89 4.5005
R5377 VSS.n223 VSS.n89 4.5005
R5378 VSS.n164 VSS.n89 4.5005
R5379 VSS.n224 VSS.n89 4.5005
R5380 VSS.n163 VSS.n89 4.5005
R5381 VSS.n225 VSS.n89 4.5005
R5382 VSS.n162 VSS.n89 4.5005
R5383 VSS.n226 VSS.n89 4.5005
R5384 VSS.n161 VSS.n89 4.5005
R5385 VSS.n227 VSS.n89 4.5005
R5386 VSS.n160 VSS.n89 4.5005
R5387 VSS.n228 VSS.n89 4.5005
R5388 VSS.n159 VSS.n89 4.5005
R5389 VSS.n229 VSS.n89 4.5005
R5390 VSS.n158 VSS.n89 4.5005
R5391 VSS.n230 VSS.n89 4.5005
R5392 VSS.n157 VSS.n89 4.5005
R5393 VSS.n231 VSS.n89 4.5005
R5394 VSS.n156 VSS.n89 4.5005
R5395 VSS.n232 VSS.n89 4.5005
R5396 VSS.n155 VSS.n89 4.5005
R5397 VSS.n233 VSS.n89 4.5005
R5398 VSS.n154 VSS.n89 4.5005
R5399 VSS.n234 VSS.n89 4.5005
R5400 VSS.n153 VSS.n89 4.5005
R5401 VSS.n235 VSS.n89 4.5005
R5402 VSS.n4506 VSS.n89 4.5005
R5403 VSS.n236 VSS.n89 4.5005
R5404 VSS.n152 VSS.n89 4.5005
R5405 VSS.n237 VSS.n89 4.5005
R5406 VSS.n151 VSS.n89 4.5005
R5407 VSS.n238 VSS.n89 4.5005
R5408 VSS.n150 VSS.n89 4.5005
R5409 VSS.n239 VSS.n89 4.5005
R5410 VSS.n149 VSS.n89 4.5005
R5411 VSS.n240 VSS.n89 4.5005
R5412 VSS.n148 VSS.n89 4.5005
R5413 VSS.n241 VSS.n89 4.5005
R5414 VSS.n147 VSS.n89 4.5005
R5415 VSS.n242 VSS.n89 4.5005
R5416 VSS.n146 VSS.n89 4.5005
R5417 VSS.n243 VSS.n89 4.5005
R5418 VSS.n145 VSS.n89 4.5005
R5419 VSS.n244 VSS.n89 4.5005
R5420 VSS.n144 VSS.n89 4.5005
R5421 VSS.n245 VSS.n89 4.5005
R5422 VSS.n143 VSS.n89 4.5005
R5423 VSS.n246 VSS.n89 4.5005
R5424 VSS.n142 VSS.n89 4.5005
R5425 VSS.n247 VSS.n89 4.5005
R5426 VSS.n141 VSS.n89 4.5005
R5427 VSS.n248 VSS.n89 4.5005
R5428 VSS.n140 VSS.n89 4.5005
R5429 VSS.n249 VSS.n89 4.5005
R5430 VSS.n139 VSS.n89 4.5005
R5431 VSS.n250 VSS.n89 4.5005
R5432 VSS.n138 VSS.n89 4.5005
R5433 VSS.n251 VSS.n89 4.5005
R5434 VSS.n137 VSS.n89 4.5005
R5435 VSS.n252 VSS.n89 4.5005
R5436 VSS.n136 VSS.n89 4.5005
R5437 VSS.n253 VSS.n89 4.5005
R5438 VSS.n135 VSS.n89 4.5005
R5439 VSS.n254 VSS.n89 4.5005
R5440 VSS.n134 VSS.n89 4.5005
R5441 VSS.n255 VSS.n89 4.5005
R5442 VSS.n133 VSS.n89 4.5005
R5443 VSS.n256 VSS.n89 4.5005
R5444 VSS.n132 VSS.n89 4.5005
R5445 VSS.n4502 VSS.n89 4.5005
R5446 VSS.n4504 VSS.n89 4.5005
R5447 VSS.n193 VSS.n47 4.5005
R5448 VSS.n195 VSS.n47 4.5005
R5449 VSS.n192 VSS.n47 4.5005
R5450 VSS.n196 VSS.n47 4.5005
R5451 VSS.n191 VSS.n47 4.5005
R5452 VSS.n197 VSS.n47 4.5005
R5453 VSS.n190 VSS.n47 4.5005
R5454 VSS.n198 VSS.n47 4.5005
R5455 VSS.n189 VSS.n47 4.5005
R5456 VSS.n199 VSS.n47 4.5005
R5457 VSS.n188 VSS.n47 4.5005
R5458 VSS.n200 VSS.n47 4.5005
R5459 VSS.n187 VSS.n47 4.5005
R5460 VSS.n201 VSS.n47 4.5005
R5461 VSS.n186 VSS.n47 4.5005
R5462 VSS.n202 VSS.n47 4.5005
R5463 VSS.n185 VSS.n47 4.5005
R5464 VSS.n203 VSS.n47 4.5005
R5465 VSS.n184 VSS.n47 4.5005
R5466 VSS.n204 VSS.n47 4.5005
R5467 VSS.n183 VSS.n47 4.5005
R5468 VSS.n205 VSS.n47 4.5005
R5469 VSS.n182 VSS.n47 4.5005
R5470 VSS.n206 VSS.n47 4.5005
R5471 VSS.n181 VSS.n47 4.5005
R5472 VSS.n207 VSS.n47 4.5005
R5473 VSS.n180 VSS.n47 4.5005
R5474 VSS.n208 VSS.n47 4.5005
R5475 VSS.n179 VSS.n47 4.5005
R5476 VSS.n209 VSS.n47 4.5005
R5477 VSS.n178 VSS.n47 4.5005
R5478 VSS.n210 VSS.n47 4.5005
R5479 VSS.n177 VSS.n47 4.5005
R5480 VSS.n211 VSS.n47 4.5005
R5481 VSS.n176 VSS.n47 4.5005
R5482 VSS.n212 VSS.n47 4.5005
R5483 VSS.n175 VSS.n47 4.5005
R5484 VSS.n213 VSS.n47 4.5005
R5485 VSS.n174 VSS.n47 4.5005
R5486 VSS.n214 VSS.n47 4.5005
R5487 VSS.n173 VSS.n47 4.5005
R5488 VSS.n215 VSS.n47 4.5005
R5489 VSS.n172 VSS.n47 4.5005
R5490 VSS.n216 VSS.n47 4.5005
R5491 VSS.n171 VSS.n47 4.5005
R5492 VSS.n217 VSS.n47 4.5005
R5493 VSS.n170 VSS.n47 4.5005
R5494 VSS.n218 VSS.n47 4.5005
R5495 VSS.n169 VSS.n47 4.5005
R5496 VSS.n219 VSS.n47 4.5005
R5497 VSS.n168 VSS.n47 4.5005
R5498 VSS.n220 VSS.n47 4.5005
R5499 VSS.n167 VSS.n47 4.5005
R5500 VSS.n221 VSS.n47 4.5005
R5501 VSS.n166 VSS.n47 4.5005
R5502 VSS.n222 VSS.n47 4.5005
R5503 VSS.n165 VSS.n47 4.5005
R5504 VSS.n223 VSS.n47 4.5005
R5505 VSS.n164 VSS.n47 4.5005
R5506 VSS.n224 VSS.n47 4.5005
R5507 VSS.n163 VSS.n47 4.5005
R5508 VSS.n225 VSS.n47 4.5005
R5509 VSS.n162 VSS.n47 4.5005
R5510 VSS.n226 VSS.n47 4.5005
R5511 VSS.n161 VSS.n47 4.5005
R5512 VSS.n227 VSS.n47 4.5005
R5513 VSS.n160 VSS.n47 4.5005
R5514 VSS.n228 VSS.n47 4.5005
R5515 VSS.n159 VSS.n47 4.5005
R5516 VSS.n229 VSS.n47 4.5005
R5517 VSS.n158 VSS.n47 4.5005
R5518 VSS.n230 VSS.n47 4.5005
R5519 VSS.n157 VSS.n47 4.5005
R5520 VSS.n231 VSS.n47 4.5005
R5521 VSS.n156 VSS.n47 4.5005
R5522 VSS.n232 VSS.n47 4.5005
R5523 VSS.n155 VSS.n47 4.5005
R5524 VSS.n233 VSS.n47 4.5005
R5525 VSS.n154 VSS.n47 4.5005
R5526 VSS.n234 VSS.n47 4.5005
R5527 VSS.n153 VSS.n47 4.5005
R5528 VSS.n235 VSS.n47 4.5005
R5529 VSS.n4506 VSS.n47 4.5005
R5530 VSS.n236 VSS.n47 4.5005
R5531 VSS.n152 VSS.n47 4.5005
R5532 VSS.n237 VSS.n47 4.5005
R5533 VSS.n151 VSS.n47 4.5005
R5534 VSS.n238 VSS.n47 4.5005
R5535 VSS.n150 VSS.n47 4.5005
R5536 VSS.n239 VSS.n47 4.5005
R5537 VSS.n149 VSS.n47 4.5005
R5538 VSS.n240 VSS.n47 4.5005
R5539 VSS.n148 VSS.n47 4.5005
R5540 VSS.n241 VSS.n47 4.5005
R5541 VSS.n147 VSS.n47 4.5005
R5542 VSS.n242 VSS.n47 4.5005
R5543 VSS.n146 VSS.n47 4.5005
R5544 VSS.n243 VSS.n47 4.5005
R5545 VSS.n145 VSS.n47 4.5005
R5546 VSS.n244 VSS.n47 4.5005
R5547 VSS.n144 VSS.n47 4.5005
R5548 VSS.n245 VSS.n47 4.5005
R5549 VSS.n143 VSS.n47 4.5005
R5550 VSS.n246 VSS.n47 4.5005
R5551 VSS.n142 VSS.n47 4.5005
R5552 VSS.n247 VSS.n47 4.5005
R5553 VSS.n141 VSS.n47 4.5005
R5554 VSS.n248 VSS.n47 4.5005
R5555 VSS.n140 VSS.n47 4.5005
R5556 VSS.n249 VSS.n47 4.5005
R5557 VSS.n139 VSS.n47 4.5005
R5558 VSS.n250 VSS.n47 4.5005
R5559 VSS.n138 VSS.n47 4.5005
R5560 VSS.n251 VSS.n47 4.5005
R5561 VSS.n137 VSS.n47 4.5005
R5562 VSS.n252 VSS.n47 4.5005
R5563 VSS.n136 VSS.n47 4.5005
R5564 VSS.n253 VSS.n47 4.5005
R5565 VSS.n135 VSS.n47 4.5005
R5566 VSS.n254 VSS.n47 4.5005
R5567 VSS.n134 VSS.n47 4.5005
R5568 VSS.n255 VSS.n47 4.5005
R5569 VSS.n133 VSS.n47 4.5005
R5570 VSS.n256 VSS.n47 4.5005
R5571 VSS.n132 VSS.n47 4.5005
R5572 VSS.n4502 VSS.n47 4.5005
R5573 VSS.n4504 VSS.n47 4.5005
R5574 VSS.n193 VSS.n90 4.5005
R5575 VSS.n195 VSS.n90 4.5005
R5576 VSS.n192 VSS.n90 4.5005
R5577 VSS.n196 VSS.n90 4.5005
R5578 VSS.n191 VSS.n90 4.5005
R5579 VSS.n197 VSS.n90 4.5005
R5580 VSS.n190 VSS.n90 4.5005
R5581 VSS.n198 VSS.n90 4.5005
R5582 VSS.n189 VSS.n90 4.5005
R5583 VSS.n199 VSS.n90 4.5005
R5584 VSS.n188 VSS.n90 4.5005
R5585 VSS.n200 VSS.n90 4.5005
R5586 VSS.n187 VSS.n90 4.5005
R5587 VSS.n201 VSS.n90 4.5005
R5588 VSS.n186 VSS.n90 4.5005
R5589 VSS.n202 VSS.n90 4.5005
R5590 VSS.n185 VSS.n90 4.5005
R5591 VSS.n203 VSS.n90 4.5005
R5592 VSS.n184 VSS.n90 4.5005
R5593 VSS.n204 VSS.n90 4.5005
R5594 VSS.n183 VSS.n90 4.5005
R5595 VSS.n205 VSS.n90 4.5005
R5596 VSS.n182 VSS.n90 4.5005
R5597 VSS.n206 VSS.n90 4.5005
R5598 VSS.n181 VSS.n90 4.5005
R5599 VSS.n207 VSS.n90 4.5005
R5600 VSS.n180 VSS.n90 4.5005
R5601 VSS.n208 VSS.n90 4.5005
R5602 VSS.n179 VSS.n90 4.5005
R5603 VSS.n209 VSS.n90 4.5005
R5604 VSS.n178 VSS.n90 4.5005
R5605 VSS.n210 VSS.n90 4.5005
R5606 VSS.n177 VSS.n90 4.5005
R5607 VSS.n211 VSS.n90 4.5005
R5608 VSS.n176 VSS.n90 4.5005
R5609 VSS.n212 VSS.n90 4.5005
R5610 VSS.n175 VSS.n90 4.5005
R5611 VSS.n213 VSS.n90 4.5005
R5612 VSS.n174 VSS.n90 4.5005
R5613 VSS.n214 VSS.n90 4.5005
R5614 VSS.n173 VSS.n90 4.5005
R5615 VSS.n215 VSS.n90 4.5005
R5616 VSS.n172 VSS.n90 4.5005
R5617 VSS.n216 VSS.n90 4.5005
R5618 VSS.n171 VSS.n90 4.5005
R5619 VSS.n217 VSS.n90 4.5005
R5620 VSS.n170 VSS.n90 4.5005
R5621 VSS.n218 VSS.n90 4.5005
R5622 VSS.n169 VSS.n90 4.5005
R5623 VSS.n219 VSS.n90 4.5005
R5624 VSS.n168 VSS.n90 4.5005
R5625 VSS.n220 VSS.n90 4.5005
R5626 VSS.n167 VSS.n90 4.5005
R5627 VSS.n221 VSS.n90 4.5005
R5628 VSS.n166 VSS.n90 4.5005
R5629 VSS.n222 VSS.n90 4.5005
R5630 VSS.n165 VSS.n90 4.5005
R5631 VSS.n223 VSS.n90 4.5005
R5632 VSS.n164 VSS.n90 4.5005
R5633 VSS.n224 VSS.n90 4.5005
R5634 VSS.n163 VSS.n90 4.5005
R5635 VSS.n225 VSS.n90 4.5005
R5636 VSS.n162 VSS.n90 4.5005
R5637 VSS.n226 VSS.n90 4.5005
R5638 VSS.n161 VSS.n90 4.5005
R5639 VSS.n227 VSS.n90 4.5005
R5640 VSS.n160 VSS.n90 4.5005
R5641 VSS.n228 VSS.n90 4.5005
R5642 VSS.n159 VSS.n90 4.5005
R5643 VSS.n229 VSS.n90 4.5005
R5644 VSS.n158 VSS.n90 4.5005
R5645 VSS.n230 VSS.n90 4.5005
R5646 VSS.n157 VSS.n90 4.5005
R5647 VSS.n231 VSS.n90 4.5005
R5648 VSS.n156 VSS.n90 4.5005
R5649 VSS.n232 VSS.n90 4.5005
R5650 VSS.n155 VSS.n90 4.5005
R5651 VSS.n233 VSS.n90 4.5005
R5652 VSS.n154 VSS.n90 4.5005
R5653 VSS.n234 VSS.n90 4.5005
R5654 VSS.n153 VSS.n90 4.5005
R5655 VSS.n235 VSS.n90 4.5005
R5656 VSS.n4506 VSS.n90 4.5005
R5657 VSS.n236 VSS.n90 4.5005
R5658 VSS.n152 VSS.n90 4.5005
R5659 VSS.n237 VSS.n90 4.5005
R5660 VSS.n151 VSS.n90 4.5005
R5661 VSS.n238 VSS.n90 4.5005
R5662 VSS.n150 VSS.n90 4.5005
R5663 VSS.n239 VSS.n90 4.5005
R5664 VSS.n149 VSS.n90 4.5005
R5665 VSS.n240 VSS.n90 4.5005
R5666 VSS.n148 VSS.n90 4.5005
R5667 VSS.n241 VSS.n90 4.5005
R5668 VSS.n147 VSS.n90 4.5005
R5669 VSS.n242 VSS.n90 4.5005
R5670 VSS.n146 VSS.n90 4.5005
R5671 VSS.n243 VSS.n90 4.5005
R5672 VSS.n145 VSS.n90 4.5005
R5673 VSS.n244 VSS.n90 4.5005
R5674 VSS.n144 VSS.n90 4.5005
R5675 VSS.n245 VSS.n90 4.5005
R5676 VSS.n143 VSS.n90 4.5005
R5677 VSS.n246 VSS.n90 4.5005
R5678 VSS.n142 VSS.n90 4.5005
R5679 VSS.n247 VSS.n90 4.5005
R5680 VSS.n141 VSS.n90 4.5005
R5681 VSS.n248 VSS.n90 4.5005
R5682 VSS.n140 VSS.n90 4.5005
R5683 VSS.n249 VSS.n90 4.5005
R5684 VSS.n139 VSS.n90 4.5005
R5685 VSS.n250 VSS.n90 4.5005
R5686 VSS.n138 VSS.n90 4.5005
R5687 VSS.n251 VSS.n90 4.5005
R5688 VSS.n137 VSS.n90 4.5005
R5689 VSS.n252 VSS.n90 4.5005
R5690 VSS.n136 VSS.n90 4.5005
R5691 VSS.n253 VSS.n90 4.5005
R5692 VSS.n135 VSS.n90 4.5005
R5693 VSS.n254 VSS.n90 4.5005
R5694 VSS.n134 VSS.n90 4.5005
R5695 VSS.n255 VSS.n90 4.5005
R5696 VSS.n133 VSS.n90 4.5005
R5697 VSS.n256 VSS.n90 4.5005
R5698 VSS.n132 VSS.n90 4.5005
R5699 VSS.n4502 VSS.n90 4.5005
R5700 VSS.n4504 VSS.n90 4.5005
R5701 VSS.n193 VSS.n46 4.5005
R5702 VSS.n195 VSS.n46 4.5005
R5703 VSS.n192 VSS.n46 4.5005
R5704 VSS.n196 VSS.n46 4.5005
R5705 VSS.n191 VSS.n46 4.5005
R5706 VSS.n197 VSS.n46 4.5005
R5707 VSS.n190 VSS.n46 4.5005
R5708 VSS.n198 VSS.n46 4.5005
R5709 VSS.n189 VSS.n46 4.5005
R5710 VSS.n199 VSS.n46 4.5005
R5711 VSS.n188 VSS.n46 4.5005
R5712 VSS.n200 VSS.n46 4.5005
R5713 VSS.n187 VSS.n46 4.5005
R5714 VSS.n201 VSS.n46 4.5005
R5715 VSS.n186 VSS.n46 4.5005
R5716 VSS.n202 VSS.n46 4.5005
R5717 VSS.n185 VSS.n46 4.5005
R5718 VSS.n203 VSS.n46 4.5005
R5719 VSS.n184 VSS.n46 4.5005
R5720 VSS.n204 VSS.n46 4.5005
R5721 VSS.n183 VSS.n46 4.5005
R5722 VSS.n205 VSS.n46 4.5005
R5723 VSS.n182 VSS.n46 4.5005
R5724 VSS.n206 VSS.n46 4.5005
R5725 VSS.n181 VSS.n46 4.5005
R5726 VSS.n207 VSS.n46 4.5005
R5727 VSS.n180 VSS.n46 4.5005
R5728 VSS.n208 VSS.n46 4.5005
R5729 VSS.n179 VSS.n46 4.5005
R5730 VSS.n209 VSS.n46 4.5005
R5731 VSS.n178 VSS.n46 4.5005
R5732 VSS.n210 VSS.n46 4.5005
R5733 VSS.n177 VSS.n46 4.5005
R5734 VSS.n211 VSS.n46 4.5005
R5735 VSS.n176 VSS.n46 4.5005
R5736 VSS.n212 VSS.n46 4.5005
R5737 VSS.n175 VSS.n46 4.5005
R5738 VSS.n213 VSS.n46 4.5005
R5739 VSS.n174 VSS.n46 4.5005
R5740 VSS.n214 VSS.n46 4.5005
R5741 VSS.n173 VSS.n46 4.5005
R5742 VSS.n215 VSS.n46 4.5005
R5743 VSS.n172 VSS.n46 4.5005
R5744 VSS.n216 VSS.n46 4.5005
R5745 VSS.n171 VSS.n46 4.5005
R5746 VSS.n217 VSS.n46 4.5005
R5747 VSS.n170 VSS.n46 4.5005
R5748 VSS.n218 VSS.n46 4.5005
R5749 VSS.n169 VSS.n46 4.5005
R5750 VSS.n219 VSS.n46 4.5005
R5751 VSS.n168 VSS.n46 4.5005
R5752 VSS.n220 VSS.n46 4.5005
R5753 VSS.n167 VSS.n46 4.5005
R5754 VSS.n221 VSS.n46 4.5005
R5755 VSS.n166 VSS.n46 4.5005
R5756 VSS.n222 VSS.n46 4.5005
R5757 VSS.n165 VSS.n46 4.5005
R5758 VSS.n223 VSS.n46 4.5005
R5759 VSS.n164 VSS.n46 4.5005
R5760 VSS.n224 VSS.n46 4.5005
R5761 VSS.n163 VSS.n46 4.5005
R5762 VSS.n225 VSS.n46 4.5005
R5763 VSS.n162 VSS.n46 4.5005
R5764 VSS.n226 VSS.n46 4.5005
R5765 VSS.n161 VSS.n46 4.5005
R5766 VSS.n227 VSS.n46 4.5005
R5767 VSS.n160 VSS.n46 4.5005
R5768 VSS.n228 VSS.n46 4.5005
R5769 VSS.n159 VSS.n46 4.5005
R5770 VSS.n229 VSS.n46 4.5005
R5771 VSS.n158 VSS.n46 4.5005
R5772 VSS.n230 VSS.n46 4.5005
R5773 VSS.n157 VSS.n46 4.5005
R5774 VSS.n231 VSS.n46 4.5005
R5775 VSS.n156 VSS.n46 4.5005
R5776 VSS.n232 VSS.n46 4.5005
R5777 VSS.n155 VSS.n46 4.5005
R5778 VSS.n233 VSS.n46 4.5005
R5779 VSS.n154 VSS.n46 4.5005
R5780 VSS.n234 VSS.n46 4.5005
R5781 VSS.n153 VSS.n46 4.5005
R5782 VSS.n235 VSS.n46 4.5005
R5783 VSS.n4506 VSS.n46 4.5005
R5784 VSS.n236 VSS.n46 4.5005
R5785 VSS.n152 VSS.n46 4.5005
R5786 VSS.n237 VSS.n46 4.5005
R5787 VSS.n151 VSS.n46 4.5005
R5788 VSS.n238 VSS.n46 4.5005
R5789 VSS.n150 VSS.n46 4.5005
R5790 VSS.n239 VSS.n46 4.5005
R5791 VSS.n149 VSS.n46 4.5005
R5792 VSS.n240 VSS.n46 4.5005
R5793 VSS.n148 VSS.n46 4.5005
R5794 VSS.n241 VSS.n46 4.5005
R5795 VSS.n147 VSS.n46 4.5005
R5796 VSS.n242 VSS.n46 4.5005
R5797 VSS.n146 VSS.n46 4.5005
R5798 VSS.n243 VSS.n46 4.5005
R5799 VSS.n145 VSS.n46 4.5005
R5800 VSS.n244 VSS.n46 4.5005
R5801 VSS.n144 VSS.n46 4.5005
R5802 VSS.n245 VSS.n46 4.5005
R5803 VSS.n143 VSS.n46 4.5005
R5804 VSS.n246 VSS.n46 4.5005
R5805 VSS.n142 VSS.n46 4.5005
R5806 VSS.n247 VSS.n46 4.5005
R5807 VSS.n141 VSS.n46 4.5005
R5808 VSS.n248 VSS.n46 4.5005
R5809 VSS.n140 VSS.n46 4.5005
R5810 VSS.n249 VSS.n46 4.5005
R5811 VSS.n139 VSS.n46 4.5005
R5812 VSS.n250 VSS.n46 4.5005
R5813 VSS.n138 VSS.n46 4.5005
R5814 VSS.n251 VSS.n46 4.5005
R5815 VSS.n137 VSS.n46 4.5005
R5816 VSS.n252 VSS.n46 4.5005
R5817 VSS.n136 VSS.n46 4.5005
R5818 VSS.n253 VSS.n46 4.5005
R5819 VSS.n135 VSS.n46 4.5005
R5820 VSS.n254 VSS.n46 4.5005
R5821 VSS.n134 VSS.n46 4.5005
R5822 VSS.n255 VSS.n46 4.5005
R5823 VSS.n133 VSS.n46 4.5005
R5824 VSS.n256 VSS.n46 4.5005
R5825 VSS.n132 VSS.n46 4.5005
R5826 VSS.n4502 VSS.n46 4.5005
R5827 VSS.n4504 VSS.n46 4.5005
R5828 VSS.n193 VSS.n91 4.5005
R5829 VSS.n195 VSS.n91 4.5005
R5830 VSS.n192 VSS.n91 4.5005
R5831 VSS.n196 VSS.n91 4.5005
R5832 VSS.n191 VSS.n91 4.5005
R5833 VSS.n197 VSS.n91 4.5005
R5834 VSS.n190 VSS.n91 4.5005
R5835 VSS.n198 VSS.n91 4.5005
R5836 VSS.n189 VSS.n91 4.5005
R5837 VSS.n199 VSS.n91 4.5005
R5838 VSS.n188 VSS.n91 4.5005
R5839 VSS.n200 VSS.n91 4.5005
R5840 VSS.n187 VSS.n91 4.5005
R5841 VSS.n201 VSS.n91 4.5005
R5842 VSS.n186 VSS.n91 4.5005
R5843 VSS.n202 VSS.n91 4.5005
R5844 VSS.n185 VSS.n91 4.5005
R5845 VSS.n203 VSS.n91 4.5005
R5846 VSS.n184 VSS.n91 4.5005
R5847 VSS.n204 VSS.n91 4.5005
R5848 VSS.n183 VSS.n91 4.5005
R5849 VSS.n205 VSS.n91 4.5005
R5850 VSS.n182 VSS.n91 4.5005
R5851 VSS.n206 VSS.n91 4.5005
R5852 VSS.n181 VSS.n91 4.5005
R5853 VSS.n207 VSS.n91 4.5005
R5854 VSS.n180 VSS.n91 4.5005
R5855 VSS.n208 VSS.n91 4.5005
R5856 VSS.n179 VSS.n91 4.5005
R5857 VSS.n209 VSS.n91 4.5005
R5858 VSS.n178 VSS.n91 4.5005
R5859 VSS.n210 VSS.n91 4.5005
R5860 VSS.n177 VSS.n91 4.5005
R5861 VSS.n211 VSS.n91 4.5005
R5862 VSS.n176 VSS.n91 4.5005
R5863 VSS.n212 VSS.n91 4.5005
R5864 VSS.n175 VSS.n91 4.5005
R5865 VSS.n213 VSS.n91 4.5005
R5866 VSS.n174 VSS.n91 4.5005
R5867 VSS.n214 VSS.n91 4.5005
R5868 VSS.n173 VSS.n91 4.5005
R5869 VSS.n215 VSS.n91 4.5005
R5870 VSS.n172 VSS.n91 4.5005
R5871 VSS.n216 VSS.n91 4.5005
R5872 VSS.n171 VSS.n91 4.5005
R5873 VSS.n217 VSS.n91 4.5005
R5874 VSS.n170 VSS.n91 4.5005
R5875 VSS.n218 VSS.n91 4.5005
R5876 VSS.n169 VSS.n91 4.5005
R5877 VSS.n219 VSS.n91 4.5005
R5878 VSS.n168 VSS.n91 4.5005
R5879 VSS.n220 VSS.n91 4.5005
R5880 VSS.n167 VSS.n91 4.5005
R5881 VSS.n221 VSS.n91 4.5005
R5882 VSS.n166 VSS.n91 4.5005
R5883 VSS.n222 VSS.n91 4.5005
R5884 VSS.n165 VSS.n91 4.5005
R5885 VSS.n223 VSS.n91 4.5005
R5886 VSS.n164 VSS.n91 4.5005
R5887 VSS.n224 VSS.n91 4.5005
R5888 VSS.n163 VSS.n91 4.5005
R5889 VSS.n225 VSS.n91 4.5005
R5890 VSS.n162 VSS.n91 4.5005
R5891 VSS.n226 VSS.n91 4.5005
R5892 VSS.n161 VSS.n91 4.5005
R5893 VSS.n227 VSS.n91 4.5005
R5894 VSS.n160 VSS.n91 4.5005
R5895 VSS.n228 VSS.n91 4.5005
R5896 VSS.n159 VSS.n91 4.5005
R5897 VSS.n229 VSS.n91 4.5005
R5898 VSS.n158 VSS.n91 4.5005
R5899 VSS.n230 VSS.n91 4.5005
R5900 VSS.n157 VSS.n91 4.5005
R5901 VSS.n231 VSS.n91 4.5005
R5902 VSS.n156 VSS.n91 4.5005
R5903 VSS.n232 VSS.n91 4.5005
R5904 VSS.n155 VSS.n91 4.5005
R5905 VSS.n233 VSS.n91 4.5005
R5906 VSS.n154 VSS.n91 4.5005
R5907 VSS.n234 VSS.n91 4.5005
R5908 VSS.n153 VSS.n91 4.5005
R5909 VSS.n235 VSS.n91 4.5005
R5910 VSS.n4506 VSS.n91 4.5005
R5911 VSS.n236 VSS.n91 4.5005
R5912 VSS.n152 VSS.n91 4.5005
R5913 VSS.n237 VSS.n91 4.5005
R5914 VSS.n151 VSS.n91 4.5005
R5915 VSS.n238 VSS.n91 4.5005
R5916 VSS.n150 VSS.n91 4.5005
R5917 VSS.n239 VSS.n91 4.5005
R5918 VSS.n149 VSS.n91 4.5005
R5919 VSS.n240 VSS.n91 4.5005
R5920 VSS.n148 VSS.n91 4.5005
R5921 VSS.n241 VSS.n91 4.5005
R5922 VSS.n147 VSS.n91 4.5005
R5923 VSS.n242 VSS.n91 4.5005
R5924 VSS.n146 VSS.n91 4.5005
R5925 VSS.n243 VSS.n91 4.5005
R5926 VSS.n145 VSS.n91 4.5005
R5927 VSS.n244 VSS.n91 4.5005
R5928 VSS.n144 VSS.n91 4.5005
R5929 VSS.n245 VSS.n91 4.5005
R5930 VSS.n143 VSS.n91 4.5005
R5931 VSS.n246 VSS.n91 4.5005
R5932 VSS.n142 VSS.n91 4.5005
R5933 VSS.n247 VSS.n91 4.5005
R5934 VSS.n141 VSS.n91 4.5005
R5935 VSS.n248 VSS.n91 4.5005
R5936 VSS.n140 VSS.n91 4.5005
R5937 VSS.n249 VSS.n91 4.5005
R5938 VSS.n139 VSS.n91 4.5005
R5939 VSS.n250 VSS.n91 4.5005
R5940 VSS.n138 VSS.n91 4.5005
R5941 VSS.n251 VSS.n91 4.5005
R5942 VSS.n137 VSS.n91 4.5005
R5943 VSS.n252 VSS.n91 4.5005
R5944 VSS.n136 VSS.n91 4.5005
R5945 VSS.n253 VSS.n91 4.5005
R5946 VSS.n135 VSS.n91 4.5005
R5947 VSS.n254 VSS.n91 4.5005
R5948 VSS.n134 VSS.n91 4.5005
R5949 VSS.n255 VSS.n91 4.5005
R5950 VSS.n133 VSS.n91 4.5005
R5951 VSS.n256 VSS.n91 4.5005
R5952 VSS.n132 VSS.n91 4.5005
R5953 VSS.n4502 VSS.n91 4.5005
R5954 VSS.n4504 VSS.n91 4.5005
R5955 VSS.n193 VSS.n45 4.5005
R5956 VSS.n195 VSS.n45 4.5005
R5957 VSS.n192 VSS.n45 4.5005
R5958 VSS.n196 VSS.n45 4.5005
R5959 VSS.n191 VSS.n45 4.5005
R5960 VSS.n197 VSS.n45 4.5005
R5961 VSS.n190 VSS.n45 4.5005
R5962 VSS.n198 VSS.n45 4.5005
R5963 VSS.n189 VSS.n45 4.5005
R5964 VSS.n199 VSS.n45 4.5005
R5965 VSS.n188 VSS.n45 4.5005
R5966 VSS.n200 VSS.n45 4.5005
R5967 VSS.n187 VSS.n45 4.5005
R5968 VSS.n201 VSS.n45 4.5005
R5969 VSS.n186 VSS.n45 4.5005
R5970 VSS.n202 VSS.n45 4.5005
R5971 VSS.n185 VSS.n45 4.5005
R5972 VSS.n203 VSS.n45 4.5005
R5973 VSS.n184 VSS.n45 4.5005
R5974 VSS.n204 VSS.n45 4.5005
R5975 VSS.n183 VSS.n45 4.5005
R5976 VSS.n205 VSS.n45 4.5005
R5977 VSS.n182 VSS.n45 4.5005
R5978 VSS.n206 VSS.n45 4.5005
R5979 VSS.n181 VSS.n45 4.5005
R5980 VSS.n207 VSS.n45 4.5005
R5981 VSS.n180 VSS.n45 4.5005
R5982 VSS.n208 VSS.n45 4.5005
R5983 VSS.n179 VSS.n45 4.5005
R5984 VSS.n209 VSS.n45 4.5005
R5985 VSS.n178 VSS.n45 4.5005
R5986 VSS.n210 VSS.n45 4.5005
R5987 VSS.n177 VSS.n45 4.5005
R5988 VSS.n211 VSS.n45 4.5005
R5989 VSS.n176 VSS.n45 4.5005
R5990 VSS.n212 VSS.n45 4.5005
R5991 VSS.n175 VSS.n45 4.5005
R5992 VSS.n213 VSS.n45 4.5005
R5993 VSS.n174 VSS.n45 4.5005
R5994 VSS.n214 VSS.n45 4.5005
R5995 VSS.n173 VSS.n45 4.5005
R5996 VSS.n215 VSS.n45 4.5005
R5997 VSS.n172 VSS.n45 4.5005
R5998 VSS.n216 VSS.n45 4.5005
R5999 VSS.n171 VSS.n45 4.5005
R6000 VSS.n217 VSS.n45 4.5005
R6001 VSS.n170 VSS.n45 4.5005
R6002 VSS.n218 VSS.n45 4.5005
R6003 VSS.n169 VSS.n45 4.5005
R6004 VSS.n219 VSS.n45 4.5005
R6005 VSS.n168 VSS.n45 4.5005
R6006 VSS.n220 VSS.n45 4.5005
R6007 VSS.n167 VSS.n45 4.5005
R6008 VSS.n221 VSS.n45 4.5005
R6009 VSS.n166 VSS.n45 4.5005
R6010 VSS.n222 VSS.n45 4.5005
R6011 VSS.n165 VSS.n45 4.5005
R6012 VSS.n223 VSS.n45 4.5005
R6013 VSS.n164 VSS.n45 4.5005
R6014 VSS.n224 VSS.n45 4.5005
R6015 VSS.n163 VSS.n45 4.5005
R6016 VSS.n225 VSS.n45 4.5005
R6017 VSS.n162 VSS.n45 4.5005
R6018 VSS.n226 VSS.n45 4.5005
R6019 VSS.n161 VSS.n45 4.5005
R6020 VSS.n227 VSS.n45 4.5005
R6021 VSS.n160 VSS.n45 4.5005
R6022 VSS.n228 VSS.n45 4.5005
R6023 VSS.n159 VSS.n45 4.5005
R6024 VSS.n229 VSS.n45 4.5005
R6025 VSS.n158 VSS.n45 4.5005
R6026 VSS.n230 VSS.n45 4.5005
R6027 VSS.n157 VSS.n45 4.5005
R6028 VSS.n231 VSS.n45 4.5005
R6029 VSS.n156 VSS.n45 4.5005
R6030 VSS.n232 VSS.n45 4.5005
R6031 VSS.n155 VSS.n45 4.5005
R6032 VSS.n233 VSS.n45 4.5005
R6033 VSS.n154 VSS.n45 4.5005
R6034 VSS.n234 VSS.n45 4.5005
R6035 VSS.n153 VSS.n45 4.5005
R6036 VSS.n235 VSS.n45 4.5005
R6037 VSS.n4506 VSS.n45 4.5005
R6038 VSS.n236 VSS.n45 4.5005
R6039 VSS.n152 VSS.n45 4.5005
R6040 VSS.n237 VSS.n45 4.5005
R6041 VSS.n151 VSS.n45 4.5005
R6042 VSS.n238 VSS.n45 4.5005
R6043 VSS.n150 VSS.n45 4.5005
R6044 VSS.n239 VSS.n45 4.5005
R6045 VSS.n149 VSS.n45 4.5005
R6046 VSS.n240 VSS.n45 4.5005
R6047 VSS.n148 VSS.n45 4.5005
R6048 VSS.n241 VSS.n45 4.5005
R6049 VSS.n147 VSS.n45 4.5005
R6050 VSS.n242 VSS.n45 4.5005
R6051 VSS.n146 VSS.n45 4.5005
R6052 VSS.n243 VSS.n45 4.5005
R6053 VSS.n145 VSS.n45 4.5005
R6054 VSS.n244 VSS.n45 4.5005
R6055 VSS.n144 VSS.n45 4.5005
R6056 VSS.n245 VSS.n45 4.5005
R6057 VSS.n143 VSS.n45 4.5005
R6058 VSS.n246 VSS.n45 4.5005
R6059 VSS.n142 VSS.n45 4.5005
R6060 VSS.n247 VSS.n45 4.5005
R6061 VSS.n141 VSS.n45 4.5005
R6062 VSS.n248 VSS.n45 4.5005
R6063 VSS.n140 VSS.n45 4.5005
R6064 VSS.n249 VSS.n45 4.5005
R6065 VSS.n139 VSS.n45 4.5005
R6066 VSS.n250 VSS.n45 4.5005
R6067 VSS.n138 VSS.n45 4.5005
R6068 VSS.n251 VSS.n45 4.5005
R6069 VSS.n137 VSS.n45 4.5005
R6070 VSS.n252 VSS.n45 4.5005
R6071 VSS.n136 VSS.n45 4.5005
R6072 VSS.n253 VSS.n45 4.5005
R6073 VSS.n135 VSS.n45 4.5005
R6074 VSS.n254 VSS.n45 4.5005
R6075 VSS.n134 VSS.n45 4.5005
R6076 VSS.n255 VSS.n45 4.5005
R6077 VSS.n133 VSS.n45 4.5005
R6078 VSS.n256 VSS.n45 4.5005
R6079 VSS.n132 VSS.n45 4.5005
R6080 VSS.n4502 VSS.n45 4.5005
R6081 VSS.n4504 VSS.n45 4.5005
R6082 VSS.n193 VSS.n92 4.5005
R6083 VSS.n195 VSS.n92 4.5005
R6084 VSS.n192 VSS.n92 4.5005
R6085 VSS.n196 VSS.n92 4.5005
R6086 VSS.n191 VSS.n92 4.5005
R6087 VSS.n197 VSS.n92 4.5005
R6088 VSS.n190 VSS.n92 4.5005
R6089 VSS.n198 VSS.n92 4.5005
R6090 VSS.n189 VSS.n92 4.5005
R6091 VSS.n199 VSS.n92 4.5005
R6092 VSS.n188 VSS.n92 4.5005
R6093 VSS.n200 VSS.n92 4.5005
R6094 VSS.n187 VSS.n92 4.5005
R6095 VSS.n201 VSS.n92 4.5005
R6096 VSS.n186 VSS.n92 4.5005
R6097 VSS.n202 VSS.n92 4.5005
R6098 VSS.n185 VSS.n92 4.5005
R6099 VSS.n203 VSS.n92 4.5005
R6100 VSS.n184 VSS.n92 4.5005
R6101 VSS.n204 VSS.n92 4.5005
R6102 VSS.n183 VSS.n92 4.5005
R6103 VSS.n205 VSS.n92 4.5005
R6104 VSS.n182 VSS.n92 4.5005
R6105 VSS.n206 VSS.n92 4.5005
R6106 VSS.n181 VSS.n92 4.5005
R6107 VSS.n207 VSS.n92 4.5005
R6108 VSS.n180 VSS.n92 4.5005
R6109 VSS.n208 VSS.n92 4.5005
R6110 VSS.n179 VSS.n92 4.5005
R6111 VSS.n209 VSS.n92 4.5005
R6112 VSS.n178 VSS.n92 4.5005
R6113 VSS.n210 VSS.n92 4.5005
R6114 VSS.n177 VSS.n92 4.5005
R6115 VSS.n211 VSS.n92 4.5005
R6116 VSS.n176 VSS.n92 4.5005
R6117 VSS.n212 VSS.n92 4.5005
R6118 VSS.n175 VSS.n92 4.5005
R6119 VSS.n213 VSS.n92 4.5005
R6120 VSS.n174 VSS.n92 4.5005
R6121 VSS.n214 VSS.n92 4.5005
R6122 VSS.n173 VSS.n92 4.5005
R6123 VSS.n215 VSS.n92 4.5005
R6124 VSS.n172 VSS.n92 4.5005
R6125 VSS.n216 VSS.n92 4.5005
R6126 VSS.n171 VSS.n92 4.5005
R6127 VSS.n217 VSS.n92 4.5005
R6128 VSS.n170 VSS.n92 4.5005
R6129 VSS.n218 VSS.n92 4.5005
R6130 VSS.n169 VSS.n92 4.5005
R6131 VSS.n219 VSS.n92 4.5005
R6132 VSS.n168 VSS.n92 4.5005
R6133 VSS.n220 VSS.n92 4.5005
R6134 VSS.n167 VSS.n92 4.5005
R6135 VSS.n221 VSS.n92 4.5005
R6136 VSS.n166 VSS.n92 4.5005
R6137 VSS.n222 VSS.n92 4.5005
R6138 VSS.n165 VSS.n92 4.5005
R6139 VSS.n223 VSS.n92 4.5005
R6140 VSS.n164 VSS.n92 4.5005
R6141 VSS.n224 VSS.n92 4.5005
R6142 VSS.n163 VSS.n92 4.5005
R6143 VSS.n225 VSS.n92 4.5005
R6144 VSS.n162 VSS.n92 4.5005
R6145 VSS.n226 VSS.n92 4.5005
R6146 VSS.n161 VSS.n92 4.5005
R6147 VSS.n227 VSS.n92 4.5005
R6148 VSS.n160 VSS.n92 4.5005
R6149 VSS.n228 VSS.n92 4.5005
R6150 VSS.n159 VSS.n92 4.5005
R6151 VSS.n229 VSS.n92 4.5005
R6152 VSS.n158 VSS.n92 4.5005
R6153 VSS.n230 VSS.n92 4.5005
R6154 VSS.n157 VSS.n92 4.5005
R6155 VSS.n231 VSS.n92 4.5005
R6156 VSS.n156 VSS.n92 4.5005
R6157 VSS.n232 VSS.n92 4.5005
R6158 VSS.n155 VSS.n92 4.5005
R6159 VSS.n233 VSS.n92 4.5005
R6160 VSS.n154 VSS.n92 4.5005
R6161 VSS.n234 VSS.n92 4.5005
R6162 VSS.n153 VSS.n92 4.5005
R6163 VSS.n235 VSS.n92 4.5005
R6164 VSS.n4506 VSS.n92 4.5005
R6165 VSS.n236 VSS.n92 4.5005
R6166 VSS.n152 VSS.n92 4.5005
R6167 VSS.n237 VSS.n92 4.5005
R6168 VSS.n151 VSS.n92 4.5005
R6169 VSS.n238 VSS.n92 4.5005
R6170 VSS.n150 VSS.n92 4.5005
R6171 VSS.n239 VSS.n92 4.5005
R6172 VSS.n149 VSS.n92 4.5005
R6173 VSS.n240 VSS.n92 4.5005
R6174 VSS.n148 VSS.n92 4.5005
R6175 VSS.n241 VSS.n92 4.5005
R6176 VSS.n147 VSS.n92 4.5005
R6177 VSS.n242 VSS.n92 4.5005
R6178 VSS.n146 VSS.n92 4.5005
R6179 VSS.n243 VSS.n92 4.5005
R6180 VSS.n145 VSS.n92 4.5005
R6181 VSS.n244 VSS.n92 4.5005
R6182 VSS.n144 VSS.n92 4.5005
R6183 VSS.n245 VSS.n92 4.5005
R6184 VSS.n143 VSS.n92 4.5005
R6185 VSS.n246 VSS.n92 4.5005
R6186 VSS.n142 VSS.n92 4.5005
R6187 VSS.n247 VSS.n92 4.5005
R6188 VSS.n141 VSS.n92 4.5005
R6189 VSS.n248 VSS.n92 4.5005
R6190 VSS.n140 VSS.n92 4.5005
R6191 VSS.n249 VSS.n92 4.5005
R6192 VSS.n139 VSS.n92 4.5005
R6193 VSS.n250 VSS.n92 4.5005
R6194 VSS.n138 VSS.n92 4.5005
R6195 VSS.n251 VSS.n92 4.5005
R6196 VSS.n137 VSS.n92 4.5005
R6197 VSS.n252 VSS.n92 4.5005
R6198 VSS.n136 VSS.n92 4.5005
R6199 VSS.n253 VSS.n92 4.5005
R6200 VSS.n135 VSS.n92 4.5005
R6201 VSS.n254 VSS.n92 4.5005
R6202 VSS.n134 VSS.n92 4.5005
R6203 VSS.n255 VSS.n92 4.5005
R6204 VSS.n133 VSS.n92 4.5005
R6205 VSS.n256 VSS.n92 4.5005
R6206 VSS.n132 VSS.n92 4.5005
R6207 VSS.n4502 VSS.n92 4.5005
R6208 VSS.n4504 VSS.n92 4.5005
R6209 VSS.n193 VSS.n44 4.5005
R6210 VSS.n195 VSS.n44 4.5005
R6211 VSS.n192 VSS.n44 4.5005
R6212 VSS.n196 VSS.n44 4.5005
R6213 VSS.n191 VSS.n44 4.5005
R6214 VSS.n197 VSS.n44 4.5005
R6215 VSS.n190 VSS.n44 4.5005
R6216 VSS.n198 VSS.n44 4.5005
R6217 VSS.n189 VSS.n44 4.5005
R6218 VSS.n199 VSS.n44 4.5005
R6219 VSS.n188 VSS.n44 4.5005
R6220 VSS.n200 VSS.n44 4.5005
R6221 VSS.n187 VSS.n44 4.5005
R6222 VSS.n201 VSS.n44 4.5005
R6223 VSS.n186 VSS.n44 4.5005
R6224 VSS.n202 VSS.n44 4.5005
R6225 VSS.n185 VSS.n44 4.5005
R6226 VSS.n203 VSS.n44 4.5005
R6227 VSS.n184 VSS.n44 4.5005
R6228 VSS.n204 VSS.n44 4.5005
R6229 VSS.n183 VSS.n44 4.5005
R6230 VSS.n205 VSS.n44 4.5005
R6231 VSS.n182 VSS.n44 4.5005
R6232 VSS.n206 VSS.n44 4.5005
R6233 VSS.n181 VSS.n44 4.5005
R6234 VSS.n207 VSS.n44 4.5005
R6235 VSS.n180 VSS.n44 4.5005
R6236 VSS.n208 VSS.n44 4.5005
R6237 VSS.n179 VSS.n44 4.5005
R6238 VSS.n209 VSS.n44 4.5005
R6239 VSS.n178 VSS.n44 4.5005
R6240 VSS.n210 VSS.n44 4.5005
R6241 VSS.n177 VSS.n44 4.5005
R6242 VSS.n211 VSS.n44 4.5005
R6243 VSS.n176 VSS.n44 4.5005
R6244 VSS.n212 VSS.n44 4.5005
R6245 VSS.n175 VSS.n44 4.5005
R6246 VSS.n213 VSS.n44 4.5005
R6247 VSS.n174 VSS.n44 4.5005
R6248 VSS.n214 VSS.n44 4.5005
R6249 VSS.n173 VSS.n44 4.5005
R6250 VSS.n215 VSS.n44 4.5005
R6251 VSS.n172 VSS.n44 4.5005
R6252 VSS.n216 VSS.n44 4.5005
R6253 VSS.n171 VSS.n44 4.5005
R6254 VSS.n217 VSS.n44 4.5005
R6255 VSS.n170 VSS.n44 4.5005
R6256 VSS.n218 VSS.n44 4.5005
R6257 VSS.n169 VSS.n44 4.5005
R6258 VSS.n219 VSS.n44 4.5005
R6259 VSS.n168 VSS.n44 4.5005
R6260 VSS.n220 VSS.n44 4.5005
R6261 VSS.n167 VSS.n44 4.5005
R6262 VSS.n221 VSS.n44 4.5005
R6263 VSS.n166 VSS.n44 4.5005
R6264 VSS.n222 VSS.n44 4.5005
R6265 VSS.n165 VSS.n44 4.5005
R6266 VSS.n223 VSS.n44 4.5005
R6267 VSS.n164 VSS.n44 4.5005
R6268 VSS.n224 VSS.n44 4.5005
R6269 VSS.n163 VSS.n44 4.5005
R6270 VSS.n225 VSS.n44 4.5005
R6271 VSS.n162 VSS.n44 4.5005
R6272 VSS.n226 VSS.n44 4.5005
R6273 VSS.n161 VSS.n44 4.5005
R6274 VSS.n227 VSS.n44 4.5005
R6275 VSS.n160 VSS.n44 4.5005
R6276 VSS.n228 VSS.n44 4.5005
R6277 VSS.n159 VSS.n44 4.5005
R6278 VSS.n229 VSS.n44 4.5005
R6279 VSS.n158 VSS.n44 4.5005
R6280 VSS.n230 VSS.n44 4.5005
R6281 VSS.n157 VSS.n44 4.5005
R6282 VSS.n231 VSS.n44 4.5005
R6283 VSS.n156 VSS.n44 4.5005
R6284 VSS.n232 VSS.n44 4.5005
R6285 VSS.n155 VSS.n44 4.5005
R6286 VSS.n233 VSS.n44 4.5005
R6287 VSS.n154 VSS.n44 4.5005
R6288 VSS.n234 VSS.n44 4.5005
R6289 VSS.n153 VSS.n44 4.5005
R6290 VSS.n235 VSS.n44 4.5005
R6291 VSS.n4506 VSS.n44 4.5005
R6292 VSS.n236 VSS.n44 4.5005
R6293 VSS.n152 VSS.n44 4.5005
R6294 VSS.n237 VSS.n44 4.5005
R6295 VSS.n151 VSS.n44 4.5005
R6296 VSS.n238 VSS.n44 4.5005
R6297 VSS.n150 VSS.n44 4.5005
R6298 VSS.n239 VSS.n44 4.5005
R6299 VSS.n149 VSS.n44 4.5005
R6300 VSS.n240 VSS.n44 4.5005
R6301 VSS.n148 VSS.n44 4.5005
R6302 VSS.n241 VSS.n44 4.5005
R6303 VSS.n147 VSS.n44 4.5005
R6304 VSS.n242 VSS.n44 4.5005
R6305 VSS.n146 VSS.n44 4.5005
R6306 VSS.n243 VSS.n44 4.5005
R6307 VSS.n145 VSS.n44 4.5005
R6308 VSS.n244 VSS.n44 4.5005
R6309 VSS.n144 VSS.n44 4.5005
R6310 VSS.n245 VSS.n44 4.5005
R6311 VSS.n143 VSS.n44 4.5005
R6312 VSS.n246 VSS.n44 4.5005
R6313 VSS.n142 VSS.n44 4.5005
R6314 VSS.n247 VSS.n44 4.5005
R6315 VSS.n141 VSS.n44 4.5005
R6316 VSS.n248 VSS.n44 4.5005
R6317 VSS.n140 VSS.n44 4.5005
R6318 VSS.n249 VSS.n44 4.5005
R6319 VSS.n139 VSS.n44 4.5005
R6320 VSS.n250 VSS.n44 4.5005
R6321 VSS.n138 VSS.n44 4.5005
R6322 VSS.n251 VSS.n44 4.5005
R6323 VSS.n137 VSS.n44 4.5005
R6324 VSS.n252 VSS.n44 4.5005
R6325 VSS.n136 VSS.n44 4.5005
R6326 VSS.n253 VSS.n44 4.5005
R6327 VSS.n135 VSS.n44 4.5005
R6328 VSS.n254 VSS.n44 4.5005
R6329 VSS.n134 VSS.n44 4.5005
R6330 VSS.n255 VSS.n44 4.5005
R6331 VSS.n133 VSS.n44 4.5005
R6332 VSS.n256 VSS.n44 4.5005
R6333 VSS.n132 VSS.n44 4.5005
R6334 VSS.n4502 VSS.n44 4.5005
R6335 VSS.n4504 VSS.n44 4.5005
R6336 VSS.n193 VSS.n93 4.5005
R6337 VSS.n195 VSS.n93 4.5005
R6338 VSS.n192 VSS.n93 4.5005
R6339 VSS.n196 VSS.n93 4.5005
R6340 VSS.n191 VSS.n93 4.5005
R6341 VSS.n197 VSS.n93 4.5005
R6342 VSS.n190 VSS.n93 4.5005
R6343 VSS.n198 VSS.n93 4.5005
R6344 VSS.n189 VSS.n93 4.5005
R6345 VSS.n199 VSS.n93 4.5005
R6346 VSS.n188 VSS.n93 4.5005
R6347 VSS.n200 VSS.n93 4.5005
R6348 VSS.n187 VSS.n93 4.5005
R6349 VSS.n201 VSS.n93 4.5005
R6350 VSS.n186 VSS.n93 4.5005
R6351 VSS.n202 VSS.n93 4.5005
R6352 VSS.n185 VSS.n93 4.5005
R6353 VSS.n203 VSS.n93 4.5005
R6354 VSS.n184 VSS.n93 4.5005
R6355 VSS.n204 VSS.n93 4.5005
R6356 VSS.n183 VSS.n93 4.5005
R6357 VSS.n205 VSS.n93 4.5005
R6358 VSS.n182 VSS.n93 4.5005
R6359 VSS.n206 VSS.n93 4.5005
R6360 VSS.n181 VSS.n93 4.5005
R6361 VSS.n207 VSS.n93 4.5005
R6362 VSS.n180 VSS.n93 4.5005
R6363 VSS.n208 VSS.n93 4.5005
R6364 VSS.n179 VSS.n93 4.5005
R6365 VSS.n209 VSS.n93 4.5005
R6366 VSS.n178 VSS.n93 4.5005
R6367 VSS.n210 VSS.n93 4.5005
R6368 VSS.n177 VSS.n93 4.5005
R6369 VSS.n211 VSS.n93 4.5005
R6370 VSS.n176 VSS.n93 4.5005
R6371 VSS.n212 VSS.n93 4.5005
R6372 VSS.n175 VSS.n93 4.5005
R6373 VSS.n213 VSS.n93 4.5005
R6374 VSS.n174 VSS.n93 4.5005
R6375 VSS.n214 VSS.n93 4.5005
R6376 VSS.n173 VSS.n93 4.5005
R6377 VSS.n215 VSS.n93 4.5005
R6378 VSS.n172 VSS.n93 4.5005
R6379 VSS.n216 VSS.n93 4.5005
R6380 VSS.n171 VSS.n93 4.5005
R6381 VSS.n217 VSS.n93 4.5005
R6382 VSS.n170 VSS.n93 4.5005
R6383 VSS.n218 VSS.n93 4.5005
R6384 VSS.n169 VSS.n93 4.5005
R6385 VSS.n219 VSS.n93 4.5005
R6386 VSS.n168 VSS.n93 4.5005
R6387 VSS.n220 VSS.n93 4.5005
R6388 VSS.n167 VSS.n93 4.5005
R6389 VSS.n221 VSS.n93 4.5005
R6390 VSS.n166 VSS.n93 4.5005
R6391 VSS.n222 VSS.n93 4.5005
R6392 VSS.n165 VSS.n93 4.5005
R6393 VSS.n223 VSS.n93 4.5005
R6394 VSS.n164 VSS.n93 4.5005
R6395 VSS.n224 VSS.n93 4.5005
R6396 VSS.n163 VSS.n93 4.5005
R6397 VSS.n225 VSS.n93 4.5005
R6398 VSS.n162 VSS.n93 4.5005
R6399 VSS.n226 VSS.n93 4.5005
R6400 VSS.n161 VSS.n93 4.5005
R6401 VSS.n227 VSS.n93 4.5005
R6402 VSS.n160 VSS.n93 4.5005
R6403 VSS.n228 VSS.n93 4.5005
R6404 VSS.n159 VSS.n93 4.5005
R6405 VSS.n229 VSS.n93 4.5005
R6406 VSS.n158 VSS.n93 4.5005
R6407 VSS.n230 VSS.n93 4.5005
R6408 VSS.n157 VSS.n93 4.5005
R6409 VSS.n231 VSS.n93 4.5005
R6410 VSS.n156 VSS.n93 4.5005
R6411 VSS.n232 VSS.n93 4.5005
R6412 VSS.n155 VSS.n93 4.5005
R6413 VSS.n233 VSS.n93 4.5005
R6414 VSS.n154 VSS.n93 4.5005
R6415 VSS.n234 VSS.n93 4.5005
R6416 VSS.n153 VSS.n93 4.5005
R6417 VSS.n235 VSS.n93 4.5005
R6418 VSS.n4506 VSS.n93 4.5005
R6419 VSS.n236 VSS.n93 4.5005
R6420 VSS.n152 VSS.n93 4.5005
R6421 VSS.n237 VSS.n93 4.5005
R6422 VSS.n151 VSS.n93 4.5005
R6423 VSS.n238 VSS.n93 4.5005
R6424 VSS.n150 VSS.n93 4.5005
R6425 VSS.n239 VSS.n93 4.5005
R6426 VSS.n149 VSS.n93 4.5005
R6427 VSS.n240 VSS.n93 4.5005
R6428 VSS.n148 VSS.n93 4.5005
R6429 VSS.n241 VSS.n93 4.5005
R6430 VSS.n147 VSS.n93 4.5005
R6431 VSS.n242 VSS.n93 4.5005
R6432 VSS.n146 VSS.n93 4.5005
R6433 VSS.n243 VSS.n93 4.5005
R6434 VSS.n145 VSS.n93 4.5005
R6435 VSS.n244 VSS.n93 4.5005
R6436 VSS.n144 VSS.n93 4.5005
R6437 VSS.n245 VSS.n93 4.5005
R6438 VSS.n143 VSS.n93 4.5005
R6439 VSS.n246 VSS.n93 4.5005
R6440 VSS.n142 VSS.n93 4.5005
R6441 VSS.n247 VSS.n93 4.5005
R6442 VSS.n141 VSS.n93 4.5005
R6443 VSS.n248 VSS.n93 4.5005
R6444 VSS.n140 VSS.n93 4.5005
R6445 VSS.n249 VSS.n93 4.5005
R6446 VSS.n139 VSS.n93 4.5005
R6447 VSS.n250 VSS.n93 4.5005
R6448 VSS.n138 VSS.n93 4.5005
R6449 VSS.n251 VSS.n93 4.5005
R6450 VSS.n137 VSS.n93 4.5005
R6451 VSS.n252 VSS.n93 4.5005
R6452 VSS.n136 VSS.n93 4.5005
R6453 VSS.n253 VSS.n93 4.5005
R6454 VSS.n135 VSS.n93 4.5005
R6455 VSS.n254 VSS.n93 4.5005
R6456 VSS.n134 VSS.n93 4.5005
R6457 VSS.n255 VSS.n93 4.5005
R6458 VSS.n133 VSS.n93 4.5005
R6459 VSS.n256 VSS.n93 4.5005
R6460 VSS.n132 VSS.n93 4.5005
R6461 VSS.n4502 VSS.n93 4.5005
R6462 VSS.n4504 VSS.n93 4.5005
R6463 VSS.n193 VSS.n43 4.5005
R6464 VSS.n195 VSS.n43 4.5005
R6465 VSS.n192 VSS.n43 4.5005
R6466 VSS.n196 VSS.n43 4.5005
R6467 VSS.n191 VSS.n43 4.5005
R6468 VSS.n197 VSS.n43 4.5005
R6469 VSS.n190 VSS.n43 4.5005
R6470 VSS.n198 VSS.n43 4.5005
R6471 VSS.n189 VSS.n43 4.5005
R6472 VSS.n199 VSS.n43 4.5005
R6473 VSS.n188 VSS.n43 4.5005
R6474 VSS.n200 VSS.n43 4.5005
R6475 VSS.n187 VSS.n43 4.5005
R6476 VSS.n201 VSS.n43 4.5005
R6477 VSS.n186 VSS.n43 4.5005
R6478 VSS.n202 VSS.n43 4.5005
R6479 VSS.n185 VSS.n43 4.5005
R6480 VSS.n203 VSS.n43 4.5005
R6481 VSS.n184 VSS.n43 4.5005
R6482 VSS.n204 VSS.n43 4.5005
R6483 VSS.n183 VSS.n43 4.5005
R6484 VSS.n205 VSS.n43 4.5005
R6485 VSS.n182 VSS.n43 4.5005
R6486 VSS.n206 VSS.n43 4.5005
R6487 VSS.n181 VSS.n43 4.5005
R6488 VSS.n207 VSS.n43 4.5005
R6489 VSS.n180 VSS.n43 4.5005
R6490 VSS.n208 VSS.n43 4.5005
R6491 VSS.n179 VSS.n43 4.5005
R6492 VSS.n209 VSS.n43 4.5005
R6493 VSS.n178 VSS.n43 4.5005
R6494 VSS.n210 VSS.n43 4.5005
R6495 VSS.n177 VSS.n43 4.5005
R6496 VSS.n211 VSS.n43 4.5005
R6497 VSS.n176 VSS.n43 4.5005
R6498 VSS.n212 VSS.n43 4.5005
R6499 VSS.n175 VSS.n43 4.5005
R6500 VSS.n213 VSS.n43 4.5005
R6501 VSS.n174 VSS.n43 4.5005
R6502 VSS.n214 VSS.n43 4.5005
R6503 VSS.n173 VSS.n43 4.5005
R6504 VSS.n215 VSS.n43 4.5005
R6505 VSS.n172 VSS.n43 4.5005
R6506 VSS.n216 VSS.n43 4.5005
R6507 VSS.n171 VSS.n43 4.5005
R6508 VSS.n217 VSS.n43 4.5005
R6509 VSS.n170 VSS.n43 4.5005
R6510 VSS.n218 VSS.n43 4.5005
R6511 VSS.n169 VSS.n43 4.5005
R6512 VSS.n219 VSS.n43 4.5005
R6513 VSS.n168 VSS.n43 4.5005
R6514 VSS.n220 VSS.n43 4.5005
R6515 VSS.n167 VSS.n43 4.5005
R6516 VSS.n221 VSS.n43 4.5005
R6517 VSS.n166 VSS.n43 4.5005
R6518 VSS.n222 VSS.n43 4.5005
R6519 VSS.n165 VSS.n43 4.5005
R6520 VSS.n223 VSS.n43 4.5005
R6521 VSS.n164 VSS.n43 4.5005
R6522 VSS.n224 VSS.n43 4.5005
R6523 VSS.n163 VSS.n43 4.5005
R6524 VSS.n225 VSS.n43 4.5005
R6525 VSS.n162 VSS.n43 4.5005
R6526 VSS.n226 VSS.n43 4.5005
R6527 VSS.n161 VSS.n43 4.5005
R6528 VSS.n227 VSS.n43 4.5005
R6529 VSS.n160 VSS.n43 4.5005
R6530 VSS.n228 VSS.n43 4.5005
R6531 VSS.n159 VSS.n43 4.5005
R6532 VSS.n229 VSS.n43 4.5005
R6533 VSS.n158 VSS.n43 4.5005
R6534 VSS.n230 VSS.n43 4.5005
R6535 VSS.n157 VSS.n43 4.5005
R6536 VSS.n231 VSS.n43 4.5005
R6537 VSS.n156 VSS.n43 4.5005
R6538 VSS.n232 VSS.n43 4.5005
R6539 VSS.n155 VSS.n43 4.5005
R6540 VSS.n233 VSS.n43 4.5005
R6541 VSS.n154 VSS.n43 4.5005
R6542 VSS.n234 VSS.n43 4.5005
R6543 VSS.n153 VSS.n43 4.5005
R6544 VSS.n235 VSS.n43 4.5005
R6545 VSS.n4506 VSS.n43 4.5005
R6546 VSS.n236 VSS.n43 4.5005
R6547 VSS.n152 VSS.n43 4.5005
R6548 VSS.n237 VSS.n43 4.5005
R6549 VSS.n151 VSS.n43 4.5005
R6550 VSS.n238 VSS.n43 4.5005
R6551 VSS.n150 VSS.n43 4.5005
R6552 VSS.n239 VSS.n43 4.5005
R6553 VSS.n149 VSS.n43 4.5005
R6554 VSS.n240 VSS.n43 4.5005
R6555 VSS.n148 VSS.n43 4.5005
R6556 VSS.n241 VSS.n43 4.5005
R6557 VSS.n147 VSS.n43 4.5005
R6558 VSS.n242 VSS.n43 4.5005
R6559 VSS.n146 VSS.n43 4.5005
R6560 VSS.n243 VSS.n43 4.5005
R6561 VSS.n145 VSS.n43 4.5005
R6562 VSS.n244 VSS.n43 4.5005
R6563 VSS.n144 VSS.n43 4.5005
R6564 VSS.n245 VSS.n43 4.5005
R6565 VSS.n143 VSS.n43 4.5005
R6566 VSS.n246 VSS.n43 4.5005
R6567 VSS.n142 VSS.n43 4.5005
R6568 VSS.n247 VSS.n43 4.5005
R6569 VSS.n141 VSS.n43 4.5005
R6570 VSS.n248 VSS.n43 4.5005
R6571 VSS.n140 VSS.n43 4.5005
R6572 VSS.n249 VSS.n43 4.5005
R6573 VSS.n139 VSS.n43 4.5005
R6574 VSS.n250 VSS.n43 4.5005
R6575 VSS.n138 VSS.n43 4.5005
R6576 VSS.n251 VSS.n43 4.5005
R6577 VSS.n137 VSS.n43 4.5005
R6578 VSS.n252 VSS.n43 4.5005
R6579 VSS.n136 VSS.n43 4.5005
R6580 VSS.n253 VSS.n43 4.5005
R6581 VSS.n135 VSS.n43 4.5005
R6582 VSS.n254 VSS.n43 4.5005
R6583 VSS.n134 VSS.n43 4.5005
R6584 VSS.n255 VSS.n43 4.5005
R6585 VSS.n133 VSS.n43 4.5005
R6586 VSS.n256 VSS.n43 4.5005
R6587 VSS.n132 VSS.n43 4.5005
R6588 VSS.n4502 VSS.n43 4.5005
R6589 VSS.n4504 VSS.n43 4.5005
R6590 VSS.n193 VSS.n94 4.5005
R6591 VSS.n195 VSS.n94 4.5005
R6592 VSS.n192 VSS.n94 4.5005
R6593 VSS.n196 VSS.n94 4.5005
R6594 VSS.n191 VSS.n94 4.5005
R6595 VSS.n197 VSS.n94 4.5005
R6596 VSS.n190 VSS.n94 4.5005
R6597 VSS.n198 VSS.n94 4.5005
R6598 VSS.n189 VSS.n94 4.5005
R6599 VSS.n199 VSS.n94 4.5005
R6600 VSS.n188 VSS.n94 4.5005
R6601 VSS.n200 VSS.n94 4.5005
R6602 VSS.n187 VSS.n94 4.5005
R6603 VSS.n201 VSS.n94 4.5005
R6604 VSS.n186 VSS.n94 4.5005
R6605 VSS.n202 VSS.n94 4.5005
R6606 VSS.n185 VSS.n94 4.5005
R6607 VSS.n203 VSS.n94 4.5005
R6608 VSS.n184 VSS.n94 4.5005
R6609 VSS.n204 VSS.n94 4.5005
R6610 VSS.n183 VSS.n94 4.5005
R6611 VSS.n205 VSS.n94 4.5005
R6612 VSS.n182 VSS.n94 4.5005
R6613 VSS.n206 VSS.n94 4.5005
R6614 VSS.n181 VSS.n94 4.5005
R6615 VSS.n207 VSS.n94 4.5005
R6616 VSS.n180 VSS.n94 4.5005
R6617 VSS.n208 VSS.n94 4.5005
R6618 VSS.n179 VSS.n94 4.5005
R6619 VSS.n209 VSS.n94 4.5005
R6620 VSS.n178 VSS.n94 4.5005
R6621 VSS.n210 VSS.n94 4.5005
R6622 VSS.n177 VSS.n94 4.5005
R6623 VSS.n211 VSS.n94 4.5005
R6624 VSS.n176 VSS.n94 4.5005
R6625 VSS.n212 VSS.n94 4.5005
R6626 VSS.n175 VSS.n94 4.5005
R6627 VSS.n213 VSS.n94 4.5005
R6628 VSS.n174 VSS.n94 4.5005
R6629 VSS.n214 VSS.n94 4.5005
R6630 VSS.n173 VSS.n94 4.5005
R6631 VSS.n215 VSS.n94 4.5005
R6632 VSS.n172 VSS.n94 4.5005
R6633 VSS.n216 VSS.n94 4.5005
R6634 VSS.n171 VSS.n94 4.5005
R6635 VSS.n217 VSS.n94 4.5005
R6636 VSS.n170 VSS.n94 4.5005
R6637 VSS.n218 VSS.n94 4.5005
R6638 VSS.n169 VSS.n94 4.5005
R6639 VSS.n219 VSS.n94 4.5005
R6640 VSS.n168 VSS.n94 4.5005
R6641 VSS.n220 VSS.n94 4.5005
R6642 VSS.n167 VSS.n94 4.5005
R6643 VSS.n221 VSS.n94 4.5005
R6644 VSS.n166 VSS.n94 4.5005
R6645 VSS.n222 VSS.n94 4.5005
R6646 VSS.n165 VSS.n94 4.5005
R6647 VSS.n223 VSS.n94 4.5005
R6648 VSS.n164 VSS.n94 4.5005
R6649 VSS.n224 VSS.n94 4.5005
R6650 VSS.n163 VSS.n94 4.5005
R6651 VSS.n225 VSS.n94 4.5005
R6652 VSS.n162 VSS.n94 4.5005
R6653 VSS.n226 VSS.n94 4.5005
R6654 VSS.n161 VSS.n94 4.5005
R6655 VSS.n227 VSS.n94 4.5005
R6656 VSS.n160 VSS.n94 4.5005
R6657 VSS.n228 VSS.n94 4.5005
R6658 VSS.n159 VSS.n94 4.5005
R6659 VSS.n229 VSS.n94 4.5005
R6660 VSS.n158 VSS.n94 4.5005
R6661 VSS.n230 VSS.n94 4.5005
R6662 VSS.n157 VSS.n94 4.5005
R6663 VSS.n231 VSS.n94 4.5005
R6664 VSS.n156 VSS.n94 4.5005
R6665 VSS.n232 VSS.n94 4.5005
R6666 VSS.n155 VSS.n94 4.5005
R6667 VSS.n233 VSS.n94 4.5005
R6668 VSS.n154 VSS.n94 4.5005
R6669 VSS.n234 VSS.n94 4.5005
R6670 VSS.n153 VSS.n94 4.5005
R6671 VSS.n235 VSS.n94 4.5005
R6672 VSS.n4506 VSS.n94 4.5005
R6673 VSS.n236 VSS.n94 4.5005
R6674 VSS.n152 VSS.n94 4.5005
R6675 VSS.n237 VSS.n94 4.5005
R6676 VSS.n151 VSS.n94 4.5005
R6677 VSS.n238 VSS.n94 4.5005
R6678 VSS.n150 VSS.n94 4.5005
R6679 VSS.n239 VSS.n94 4.5005
R6680 VSS.n149 VSS.n94 4.5005
R6681 VSS.n240 VSS.n94 4.5005
R6682 VSS.n148 VSS.n94 4.5005
R6683 VSS.n241 VSS.n94 4.5005
R6684 VSS.n147 VSS.n94 4.5005
R6685 VSS.n242 VSS.n94 4.5005
R6686 VSS.n146 VSS.n94 4.5005
R6687 VSS.n243 VSS.n94 4.5005
R6688 VSS.n145 VSS.n94 4.5005
R6689 VSS.n244 VSS.n94 4.5005
R6690 VSS.n144 VSS.n94 4.5005
R6691 VSS.n245 VSS.n94 4.5005
R6692 VSS.n143 VSS.n94 4.5005
R6693 VSS.n246 VSS.n94 4.5005
R6694 VSS.n142 VSS.n94 4.5005
R6695 VSS.n247 VSS.n94 4.5005
R6696 VSS.n141 VSS.n94 4.5005
R6697 VSS.n248 VSS.n94 4.5005
R6698 VSS.n140 VSS.n94 4.5005
R6699 VSS.n249 VSS.n94 4.5005
R6700 VSS.n139 VSS.n94 4.5005
R6701 VSS.n250 VSS.n94 4.5005
R6702 VSS.n138 VSS.n94 4.5005
R6703 VSS.n251 VSS.n94 4.5005
R6704 VSS.n137 VSS.n94 4.5005
R6705 VSS.n252 VSS.n94 4.5005
R6706 VSS.n136 VSS.n94 4.5005
R6707 VSS.n253 VSS.n94 4.5005
R6708 VSS.n135 VSS.n94 4.5005
R6709 VSS.n254 VSS.n94 4.5005
R6710 VSS.n134 VSS.n94 4.5005
R6711 VSS.n255 VSS.n94 4.5005
R6712 VSS.n133 VSS.n94 4.5005
R6713 VSS.n256 VSS.n94 4.5005
R6714 VSS.n132 VSS.n94 4.5005
R6715 VSS.n4502 VSS.n94 4.5005
R6716 VSS.n4504 VSS.n94 4.5005
R6717 VSS.n193 VSS.n42 4.5005
R6718 VSS.n195 VSS.n42 4.5005
R6719 VSS.n192 VSS.n42 4.5005
R6720 VSS.n196 VSS.n42 4.5005
R6721 VSS.n191 VSS.n42 4.5005
R6722 VSS.n197 VSS.n42 4.5005
R6723 VSS.n190 VSS.n42 4.5005
R6724 VSS.n198 VSS.n42 4.5005
R6725 VSS.n189 VSS.n42 4.5005
R6726 VSS.n199 VSS.n42 4.5005
R6727 VSS.n188 VSS.n42 4.5005
R6728 VSS.n200 VSS.n42 4.5005
R6729 VSS.n187 VSS.n42 4.5005
R6730 VSS.n201 VSS.n42 4.5005
R6731 VSS.n186 VSS.n42 4.5005
R6732 VSS.n202 VSS.n42 4.5005
R6733 VSS.n185 VSS.n42 4.5005
R6734 VSS.n203 VSS.n42 4.5005
R6735 VSS.n184 VSS.n42 4.5005
R6736 VSS.n204 VSS.n42 4.5005
R6737 VSS.n183 VSS.n42 4.5005
R6738 VSS.n205 VSS.n42 4.5005
R6739 VSS.n182 VSS.n42 4.5005
R6740 VSS.n206 VSS.n42 4.5005
R6741 VSS.n181 VSS.n42 4.5005
R6742 VSS.n207 VSS.n42 4.5005
R6743 VSS.n180 VSS.n42 4.5005
R6744 VSS.n208 VSS.n42 4.5005
R6745 VSS.n179 VSS.n42 4.5005
R6746 VSS.n209 VSS.n42 4.5005
R6747 VSS.n178 VSS.n42 4.5005
R6748 VSS.n210 VSS.n42 4.5005
R6749 VSS.n177 VSS.n42 4.5005
R6750 VSS.n211 VSS.n42 4.5005
R6751 VSS.n176 VSS.n42 4.5005
R6752 VSS.n212 VSS.n42 4.5005
R6753 VSS.n175 VSS.n42 4.5005
R6754 VSS.n213 VSS.n42 4.5005
R6755 VSS.n174 VSS.n42 4.5005
R6756 VSS.n214 VSS.n42 4.5005
R6757 VSS.n173 VSS.n42 4.5005
R6758 VSS.n215 VSS.n42 4.5005
R6759 VSS.n172 VSS.n42 4.5005
R6760 VSS.n216 VSS.n42 4.5005
R6761 VSS.n171 VSS.n42 4.5005
R6762 VSS.n217 VSS.n42 4.5005
R6763 VSS.n170 VSS.n42 4.5005
R6764 VSS.n218 VSS.n42 4.5005
R6765 VSS.n169 VSS.n42 4.5005
R6766 VSS.n219 VSS.n42 4.5005
R6767 VSS.n168 VSS.n42 4.5005
R6768 VSS.n220 VSS.n42 4.5005
R6769 VSS.n167 VSS.n42 4.5005
R6770 VSS.n221 VSS.n42 4.5005
R6771 VSS.n166 VSS.n42 4.5005
R6772 VSS.n222 VSS.n42 4.5005
R6773 VSS.n165 VSS.n42 4.5005
R6774 VSS.n223 VSS.n42 4.5005
R6775 VSS.n164 VSS.n42 4.5005
R6776 VSS.n224 VSS.n42 4.5005
R6777 VSS.n163 VSS.n42 4.5005
R6778 VSS.n225 VSS.n42 4.5005
R6779 VSS.n162 VSS.n42 4.5005
R6780 VSS.n226 VSS.n42 4.5005
R6781 VSS.n161 VSS.n42 4.5005
R6782 VSS.n227 VSS.n42 4.5005
R6783 VSS.n160 VSS.n42 4.5005
R6784 VSS.n228 VSS.n42 4.5005
R6785 VSS.n159 VSS.n42 4.5005
R6786 VSS.n229 VSS.n42 4.5005
R6787 VSS.n158 VSS.n42 4.5005
R6788 VSS.n230 VSS.n42 4.5005
R6789 VSS.n157 VSS.n42 4.5005
R6790 VSS.n231 VSS.n42 4.5005
R6791 VSS.n156 VSS.n42 4.5005
R6792 VSS.n232 VSS.n42 4.5005
R6793 VSS.n155 VSS.n42 4.5005
R6794 VSS.n233 VSS.n42 4.5005
R6795 VSS.n154 VSS.n42 4.5005
R6796 VSS.n234 VSS.n42 4.5005
R6797 VSS.n153 VSS.n42 4.5005
R6798 VSS.n235 VSS.n42 4.5005
R6799 VSS.n4506 VSS.n42 4.5005
R6800 VSS.n236 VSS.n42 4.5005
R6801 VSS.n152 VSS.n42 4.5005
R6802 VSS.n237 VSS.n42 4.5005
R6803 VSS.n151 VSS.n42 4.5005
R6804 VSS.n238 VSS.n42 4.5005
R6805 VSS.n150 VSS.n42 4.5005
R6806 VSS.n239 VSS.n42 4.5005
R6807 VSS.n149 VSS.n42 4.5005
R6808 VSS.n240 VSS.n42 4.5005
R6809 VSS.n148 VSS.n42 4.5005
R6810 VSS.n241 VSS.n42 4.5005
R6811 VSS.n147 VSS.n42 4.5005
R6812 VSS.n242 VSS.n42 4.5005
R6813 VSS.n146 VSS.n42 4.5005
R6814 VSS.n243 VSS.n42 4.5005
R6815 VSS.n145 VSS.n42 4.5005
R6816 VSS.n244 VSS.n42 4.5005
R6817 VSS.n144 VSS.n42 4.5005
R6818 VSS.n245 VSS.n42 4.5005
R6819 VSS.n143 VSS.n42 4.5005
R6820 VSS.n246 VSS.n42 4.5005
R6821 VSS.n142 VSS.n42 4.5005
R6822 VSS.n247 VSS.n42 4.5005
R6823 VSS.n141 VSS.n42 4.5005
R6824 VSS.n248 VSS.n42 4.5005
R6825 VSS.n140 VSS.n42 4.5005
R6826 VSS.n249 VSS.n42 4.5005
R6827 VSS.n139 VSS.n42 4.5005
R6828 VSS.n250 VSS.n42 4.5005
R6829 VSS.n138 VSS.n42 4.5005
R6830 VSS.n251 VSS.n42 4.5005
R6831 VSS.n137 VSS.n42 4.5005
R6832 VSS.n252 VSS.n42 4.5005
R6833 VSS.n136 VSS.n42 4.5005
R6834 VSS.n253 VSS.n42 4.5005
R6835 VSS.n135 VSS.n42 4.5005
R6836 VSS.n254 VSS.n42 4.5005
R6837 VSS.n134 VSS.n42 4.5005
R6838 VSS.n255 VSS.n42 4.5005
R6839 VSS.n133 VSS.n42 4.5005
R6840 VSS.n256 VSS.n42 4.5005
R6841 VSS.n132 VSS.n42 4.5005
R6842 VSS.n4502 VSS.n42 4.5005
R6843 VSS.n4504 VSS.n42 4.5005
R6844 VSS.n193 VSS.n95 4.5005
R6845 VSS.n195 VSS.n95 4.5005
R6846 VSS.n192 VSS.n95 4.5005
R6847 VSS.n196 VSS.n95 4.5005
R6848 VSS.n191 VSS.n95 4.5005
R6849 VSS.n197 VSS.n95 4.5005
R6850 VSS.n190 VSS.n95 4.5005
R6851 VSS.n198 VSS.n95 4.5005
R6852 VSS.n189 VSS.n95 4.5005
R6853 VSS.n199 VSS.n95 4.5005
R6854 VSS.n188 VSS.n95 4.5005
R6855 VSS.n200 VSS.n95 4.5005
R6856 VSS.n187 VSS.n95 4.5005
R6857 VSS.n201 VSS.n95 4.5005
R6858 VSS.n186 VSS.n95 4.5005
R6859 VSS.n202 VSS.n95 4.5005
R6860 VSS.n185 VSS.n95 4.5005
R6861 VSS.n203 VSS.n95 4.5005
R6862 VSS.n184 VSS.n95 4.5005
R6863 VSS.n204 VSS.n95 4.5005
R6864 VSS.n183 VSS.n95 4.5005
R6865 VSS.n205 VSS.n95 4.5005
R6866 VSS.n182 VSS.n95 4.5005
R6867 VSS.n206 VSS.n95 4.5005
R6868 VSS.n181 VSS.n95 4.5005
R6869 VSS.n207 VSS.n95 4.5005
R6870 VSS.n180 VSS.n95 4.5005
R6871 VSS.n208 VSS.n95 4.5005
R6872 VSS.n179 VSS.n95 4.5005
R6873 VSS.n209 VSS.n95 4.5005
R6874 VSS.n178 VSS.n95 4.5005
R6875 VSS.n210 VSS.n95 4.5005
R6876 VSS.n177 VSS.n95 4.5005
R6877 VSS.n211 VSS.n95 4.5005
R6878 VSS.n176 VSS.n95 4.5005
R6879 VSS.n212 VSS.n95 4.5005
R6880 VSS.n175 VSS.n95 4.5005
R6881 VSS.n213 VSS.n95 4.5005
R6882 VSS.n174 VSS.n95 4.5005
R6883 VSS.n214 VSS.n95 4.5005
R6884 VSS.n173 VSS.n95 4.5005
R6885 VSS.n215 VSS.n95 4.5005
R6886 VSS.n172 VSS.n95 4.5005
R6887 VSS.n216 VSS.n95 4.5005
R6888 VSS.n171 VSS.n95 4.5005
R6889 VSS.n217 VSS.n95 4.5005
R6890 VSS.n170 VSS.n95 4.5005
R6891 VSS.n218 VSS.n95 4.5005
R6892 VSS.n169 VSS.n95 4.5005
R6893 VSS.n219 VSS.n95 4.5005
R6894 VSS.n168 VSS.n95 4.5005
R6895 VSS.n220 VSS.n95 4.5005
R6896 VSS.n167 VSS.n95 4.5005
R6897 VSS.n221 VSS.n95 4.5005
R6898 VSS.n166 VSS.n95 4.5005
R6899 VSS.n222 VSS.n95 4.5005
R6900 VSS.n165 VSS.n95 4.5005
R6901 VSS.n223 VSS.n95 4.5005
R6902 VSS.n164 VSS.n95 4.5005
R6903 VSS.n224 VSS.n95 4.5005
R6904 VSS.n163 VSS.n95 4.5005
R6905 VSS.n225 VSS.n95 4.5005
R6906 VSS.n162 VSS.n95 4.5005
R6907 VSS.n226 VSS.n95 4.5005
R6908 VSS.n161 VSS.n95 4.5005
R6909 VSS.n227 VSS.n95 4.5005
R6910 VSS.n160 VSS.n95 4.5005
R6911 VSS.n228 VSS.n95 4.5005
R6912 VSS.n159 VSS.n95 4.5005
R6913 VSS.n229 VSS.n95 4.5005
R6914 VSS.n158 VSS.n95 4.5005
R6915 VSS.n230 VSS.n95 4.5005
R6916 VSS.n157 VSS.n95 4.5005
R6917 VSS.n231 VSS.n95 4.5005
R6918 VSS.n156 VSS.n95 4.5005
R6919 VSS.n232 VSS.n95 4.5005
R6920 VSS.n155 VSS.n95 4.5005
R6921 VSS.n233 VSS.n95 4.5005
R6922 VSS.n154 VSS.n95 4.5005
R6923 VSS.n234 VSS.n95 4.5005
R6924 VSS.n153 VSS.n95 4.5005
R6925 VSS.n235 VSS.n95 4.5005
R6926 VSS.n4506 VSS.n95 4.5005
R6927 VSS.n236 VSS.n95 4.5005
R6928 VSS.n152 VSS.n95 4.5005
R6929 VSS.n237 VSS.n95 4.5005
R6930 VSS.n151 VSS.n95 4.5005
R6931 VSS.n238 VSS.n95 4.5005
R6932 VSS.n150 VSS.n95 4.5005
R6933 VSS.n239 VSS.n95 4.5005
R6934 VSS.n149 VSS.n95 4.5005
R6935 VSS.n240 VSS.n95 4.5005
R6936 VSS.n148 VSS.n95 4.5005
R6937 VSS.n241 VSS.n95 4.5005
R6938 VSS.n147 VSS.n95 4.5005
R6939 VSS.n242 VSS.n95 4.5005
R6940 VSS.n146 VSS.n95 4.5005
R6941 VSS.n243 VSS.n95 4.5005
R6942 VSS.n145 VSS.n95 4.5005
R6943 VSS.n244 VSS.n95 4.5005
R6944 VSS.n144 VSS.n95 4.5005
R6945 VSS.n245 VSS.n95 4.5005
R6946 VSS.n143 VSS.n95 4.5005
R6947 VSS.n246 VSS.n95 4.5005
R6948 VSS.n142 VSS.n95 4.5005
R6949 VSS.n247 VSS.n95 4.5005
R6950 VSS.n141 VSS.n95 4.5005
R6951 VSS.n248 VSS.n95 4.5005
R6952 VSS.n140 VSS.n95 4.5005
R6953 VSS.n249 VSS.n95 4.5005
R6954 VSS.n139 VSS.n95 4.5005
R6955 VSS.n250 VSS.n95 4.5005
R6956 VSS.n138 VSS.n95 4.5005
R6957 VSS.n251 VSS.n95 4.5005
R6958 VSS.n137 VSS.n95 4.5005
R6959 VSS.n252 VSS.n95 4.5005
R6960 VSS.n136 VSS.n95 4.5005
R6961 VSS.n253 VSS.n95 4.5005
R6962 VSS.n135 VSS.n95 4.5005
R6963 VSS.n254 VSS.n95 4.5005
R6964 VSS.n134 VSS.n95 4.5005
R6965 VSS.n255 VSS.n95 4.5005
R6966 VSS.n133 VSS.n95 4.5005
R6967 VSS.n256 VSS.n95 4.5005
R6968 VSS.n132 VSS.n95 4.5005
R6969 VSS.n4502 VSS.n95 4.5005
R6970 VSS.n4504 VSS.n95 4.5005
R6971 VSS.n193 VSS.n41 4.5005
R6972 VSS.n195 VSS.n41 4.5005
R6973 VSS.n192 VSS.n41 4.5005
R6974 VSS.n196 VSS.n41 4.5005
R6975 VSS.n191 VSS.n41 4.5005
R6976 VSS.n197 VSS.n41 4.5005
R6977 VSS.n190 VSS.n41 4.5005
R6978 VSS.n198 VSS.n41 4.5005
R6979 VSS.n189 VSS.n41 4.5005
R6980 VSS.n199 VSS.n41 4.5005
R6981 VSS.n188 VSS.n41 4.5005
R6982 VSS.n200 VSS.n41 4.5005
R6983 VSS.n187 VSS.n41 4.5005
R6984 VSS.n201 VSS.n41 4.5005
R6985 VSS.n186 VSS.n41 4.5005
R6986 VSS.n202 VSS.n41 4.5005
R6987 VSS.n185 VSS.n41 4.5005
R6988 VSS.n203 VSS.n41 4.5005
R6989 VSS.n184 VSS.n41 4.5005
R6990 VSS.n204 VSS.n41 4.5005
R6991 VSS.n183 VSS.n41 4.5005
R6992 VSS.n205 VSS.n41 4.5005
R6993 VSS.n182 VSS.n41 4.5005
R6994 VSS.n206 VSS.n41 4.5005
R6995 VSS.n181 VSS.n41 4.5005
R6996 VSS.n207 VSS.n41 4.5005
R6997 VSS.n180 VSS.n41 4.5005
R6998 VSS.n208 VSS.n41 4.5005
R6999 VSS.n179 VSS.n41 4.5005
R7000 VSS.n209 VSS.n41 4.5005
R7001 VSS.n178 VSS.n41 4.5005
R7002 VSS.n210 VSS.n41 4.5005
R7003 VSS.n177 VSS.n41 4.5005
R7004 VSS.n211 VSS.n41 4.5005
R7005 VSS.n176 VSS.n41 4.5005
R7006 VSS.n212 VSS.n41 4.5005
R7007 VSS.n175 VSS.n41 4.5005
R7008 VSS.n213 VSS.n41 4.5005
R7009 VSS.n174 VSS.n41 4.5005
R7010 VSS.n214 VSS.n41 4.5005
R7011 VSS.n173 VSS.n41 4.5005
R7012 VSS.n215 VSS.n41 4.5005
R7013 VSS.n172 VSS.n41 4.5005
R7014 VSS.n216 VSS.n41 4.5005
R7015 VSS.n171 VSS.n41 4.5005
R7016 VSS.n217 VSS.n41 4.5005
R7017 VSS.n170 VSS.n41 4.5005
R7018 VSS.n218 VSS.n41 4.5005
R7019 VSS.n169 VSS.n41 4.5005
R7020 VSS.n219 VSS.n41 4.5005
R7021 VSS.n168 VSS.n41 4.5005
R7022 VSS.n220 VSS.n41 4.5005
R7023 VSS.n167 VSS.n41 4.5005
R7024 VSS.n221 VSS.n41 4.5005
R7025 VSS.n166 VSS.n41 4.5005
R7026 VSS.n222 VSS.n41 4.5005
R7027 VSS.n165 VSS.n41 4.5005
R7028 VSS.n223 VSS.n41 4.5005
R7029 VSS.n164 VSS.n41 4.5005
R7030 VSS.n224 VSS.n41 4.5005
R7031 VSS.n163 VSS.n41 4.5005
R7032 VSS.n225 VSS.n41 4.5005
R7033 VSS.n162 VSS.n41 4.5005
R7034 VSS.n226 VSS.n41 4.5005
R7035 VSS.n161 VSS.n41 4.5005
R7036 VSS.n227 VSS.n41 4.5005
R7037 VSS.n160 VSS.n41 4.5005
R7038 VSS.n228 VSS.n41 4.5005
R7039 VSS.n159 VSS.n41 4.5005
R7040 VSS.n229 VSS.n41 4.5005
R7041 VSS.n158 VSS.n41 4.5005
R7042 VSS.n230 VSS.n41 4.5005
R7043 VSS.n157 VSS.n41 4.5005
R7044 VSS.n231 VSS.n41 4.5005
R7045 VSS.n156 VSS.n41 4.5005
R7046 VSS.n232 VSS.n41 4.5005
R7047 VSS.n155 VSS.n41 4.5005
R7048 VSS.n233 VSS.n41 4.5005
R7049 VSS.n154 VSS.n41 4.5005
R7050 VSS.n234 VSS.n41 4.5005
R7051 VSS.n153 VSS.n41 4.5005
R7052 VSS.n235 VSS.n41 4.5005
R7053 VSS.n4506 VSS.n41 4.5005
R7054 VSS.n236 VSS.n41 4.5005
R7055 VSS.n152 VSS.n41 4.5005
R7056 VSS.n237 VSS.n41 4.5005
R7057 VSS.n151 VSS.n41 4.5005
R7058 VSS.n238 VSS.n41 4.5005
R7059 VSS.n150 VSS.n41 4.5005
R7060 VSS.n239 VSS.n41 4.5005
R7061 VSS.n149 VSS.n41 4.5005
R7062 VSS.n240 VSS.n41 4.5005
R7063 VSS.n148 VSS.n41 4.5005
R7064 VSS.n241 VSS.n41 4.5005
R7065 VSS.n147 VSS.n41 4.5005
R7066 VSS.n242 VSS.n41 4.5005
R7067 VSS.n146 VSS.n41 4.5005
R7068 VSS.n243 VSS.n41 4.5005
R7069 VSS.n145 VSS.n41 4.5005
R7070 VSS.n244 VSS.n41 4.5005
R7071 VSS.n144 VSS.n41 4.5005
R7072 VSS.n245 VSS.n41 4.5005
R7073 VSS.n143 VSS.n41 4.5005
R7074 VSS.n246 VSS.n41 4.5005
R7075 VSS.n142 VSS.n41 4.5005
R7076 VSS.n247 VSS.n41 4.5005
R7077 VSS.n141 VSS.n41 4.5005
R7078 VSS.n248 VSS.n41 4.5005
R7079 VSS.n140 VSS.n41 4.5005
R7080 VSS.n249 VSS.n41 4.5005
R7081 VSS.n139 VSS.n41 4.5005
R7082 VSS.n250 VSS.n41 4.5005
R7083 VSS.n138 VSS.n41 4.5005
R7084 VSS.n251 VSS.n41 4.5005
R7085 VSS.n137 VSS.n41 4.5005
R7086 VSS.n252 VSS.n41 4.5005
R7087 VSS.n136 VSS.n41 4.5005
R7088 VSS.n253 VSS.n41 4.5005
R7089 VSS.n135 VSS.n41 4.5005
R7090 VSS.n254 VSS.n41 4.5005
R7091 VSS.n134 VSS.n41 4.5005
R7092 VSS.n255 VSS.n41 4.5005
R7093 VSS.n133 VSS.n41 4.5005
R7094 VSS.n256 VSS.n41 4.5005
R7095 VSS.n132 VSS.n41 4.5005
R7096 VSS.n4502 VSS.n41 4.5005
R7097 VSS.n4504 VSS.n41 4.5005
R7098 VSS.n193 VSS.n96 4.5005
R7099 VSS.n195 VSS.n96 4.5005
R7100 VSS.n192 VSS.n96 4.5005
R7101 VSS.n196 VSS.n96 4.5005
R7102 VSS.n191 VSS.n96 4.5005
R7103 VSS.n197 VSS.n96 4.5005
R7104 VSS.n190 VSS.n96 4.5005
R7105 VSS.n198 VSS.n96 4.5005
R7106 VSS.n189 VSS.n96 4.5005
R7107 VSS.n199 VSS.n96 4.5005
R7108 VSS.n188 VSS.n96 4.5005
R7109 VSS.n200 VSS.n96 4.5005
R7110 VSS.n187 VSS.n96 4.5005
R7111 VSS.n201 VSS.n96 4.5005
R7112 VSS.n186 VSS.n96 4.5005
R7113 VSS.n202 VSS.n96 4.5005
R7114 VSS.n185 VSS.n96 4.5005
R7115 VSS.n203 VSS.n96 4.5005
R7116 VSS.n184 VSS.n96 4.5005
R7117 VSS.n204 VSS.n96 4.5005
R7118 VSS.n183 VSS.n96 4.5005
R7119 VSS.n205 VSS.n96 4.5005
R7120 VSS.n182 VSS.n96 4.5005
R7121 VSS.n206 VSS.n96 4.5005
R7122 VSS.n181 VSS.n96 4.5005
R7123 VSS.n207 VSS.n96 4.5005
R7124 VSS.n180 VSS.n96 4.5005
R7125 VSS.n208 VSS.n96 4.5005
R7126 VSS.n179 VSS.n96 4.5005
R7127 VSS.n209 VSS.n96 4.5005
R7128 VSS.n178 VSS.n96 4.5005
R7129 VSS.n210 VSS.n96 4.5005
R7130 VSS.n177 VSS.n96 4.5005
R7131 VSS.n211 VSS.n96 4.5005
R7132 VSS.n176 VSS.n96 4.5005
R7133 VSS.n212 VSS.n96 4.5005
R7134 VSS.n175 VSS.n96 4.5005
R7135 VSS.n213 VSS.n96 4.5005
R7136 VSS.n174 VSS.n96 4.5005
R7137 VSS.n214 VSS.n96 4.5005
R7138 VSS.n173 VSS.n96 4.5005
R7139 VSS.n215 VSS.n96 4.5005
R7140 VSS.n172 VSS.n96 4.5005
R7141 VSS.n216 VSS.n96 4.5005
R7142 VSS.n171 VSS.n96 4.5005
R7143 VSS.n217 VSS.n96 4.5005
R7144 VSS.n170 VSS.n96 4.5005
R7145 VSS.n218 VSS.n96 4.5005
R7146 VSS.n169 VSS.n96 4.5005
R7147 VSS.n219 VSS.n96 4.5005
R7148 VSS.n168 VSS.n96 4.5005
R7149 VSS.n220 VSS.n96 4.5005
R7150 VSS.n167 VSS.n96 4.5005
R7151 VSS.n221 VSS.n96 4.5005
R7152 VSS.n166 VSS.n96 4.5005
R7153 VSS.n222 VSS.n96 4.5005
R7154 VSS.n165 VSS.n96 4.5005
R7155 VSS.n223 VSS.n96 4.5005
R7156 VSS.n164 VSS.n96 4.5005
R7157 VSS.n224 VSS.n96 4.5005
R7158 VSS.n163 VSS.n96 4.5005
R7159 VSS.n225 VSS.n96 4.5005
R7160 VSS.n162 VSS.n96 4.5005
R7161 VSS.n226 VSS.n96 4.5005
R7162 VSS.n161 VSS.n96 4.5005
R7163 VSS.n227 VSS.n96 4.5005
R7164 VSS.n160 VSS.n96 4.5005
R7165 VSS.n228 VSS.n96 4.5005
R7166 VSS.n159 VSS.n96 4.5005
R7167 VSS.n229 VSS.n96 4.5005
R7168 VSS.n158 VSS.n96 4.5005
R7169 VSS.n230 VSS.n96 4.5005
R7170 VSS.n157 VSS.n96 4.5005
R7171 VSS.n231 VSS.n96 4.5005
R7172 VSS.n156 VSS.n96 4.5005
R7173 VSS.n232 VSS.n96 4.5005
R7174 VSS.n155 VSS.n96 4.5005
R7175 VSS.n233 VSS.n96 4.5005
R7176 VSS.n154 VSS.n96 4.5005
R7177 VSS.n234 VSS.n96 4.5005
R7178 VSS.n153 VSS.n96 4.5005
R7179 VSS.n235 VSS.n96 4.5005
R7180 VSS.n4506 VSS.n96 4.5005
R7181 VSS.n236 VSS.n96 4.5005
R7182 VSS.n152 VSS.n96 4.5005
R7183 VSS.n237 VSS.n96 4.5005
R7184 VSS.n151 VSS.n96 4.5005
R7185 VSS.n238 VSS.n96 4.5005
R7186 VSS.n150 VSS.n96 4.5005
R7187 VSS.n239 VSS.n96 4.5005
R7188 VSS.n149 VSS.n96 4.5005
R7189 VSS.n240 VSS.n96 4.5005
R7190 VSS.n148 VSS.n96 4.5005
R7191 VSS.n241 VSS.n96 4.5005
R7192 VSS.n147 VSS.n96 4.5005
R7193 VSS.n242 VSS.n96 4.5005
R7194 VSS.n146 VSS.n96 4.5005
R7195 VSS.n243 VSS.n96 4.5005
R7196 VSS.n145 VSS.n96 4.5005
R7197 VSS.n244 VSS.n96 4.5005
R7198 VSS.n144 VSS.n96 4.5005
R7199 VSS.n245 VSS.n96 4.5005
R7200 VSS.n143 VSS.n96 4.5005
R7201 VSS.n246 VSS.n96 4.5005
R7202 VSS.n142 VSS.n96 4.5005
R7203 VSS.n247 VSS.n96 4.5005
R7204 VSS.n141 VSS.n96 4.5005
R7205 VSS.n248 VSS.n96 4.5005
R7206 VSS.n140 VSS.n96 4.5005
R7207 VSS.n249 VSS.n96 4.5005
R7208 VSS.n139 VSS.n96 4.5005
R7209 VSS.n250 VSS.n96 4.5005
R7210 VSS.n138 VSS.n96 4.5005
R7211 VSS.n251 VSS.n96 4.5005
R7212 VSS.n137 VSS.n96 4.5005
R7213 VSS.n252 VSS.n96 4.5005
R7214 VSS.n136 VSS.n96 4.5005
R7215 VSS.n253 VSS.n96 4.5005
R7216 VSS.n135 VSS.n96 4.5005
R7217 VSS.n254 VSS.n96 4.5005
R7218 VSS.n134 VSS.n96 4.5005
R7219 VSS.n255 VSS.n96 4.5005
R7220 VSS.n133 VSS.n96 4.5005
R7221 VSS.n256 VSS.n96 4.5005
R7222 VSS.n132 VSS.n96 4.5005
R7223 VSS.n4502 VSS.n96 4.5005
R7224 VSS.n4504 VSS.n96 4.5005
R7225 VSS.n193 VSS.n40 4.5005
R7226 VSS.n195 VSS.n40 4.5005
R7227 VSS.n192 VSS.n40 4.5005
R7228 VSS.n196 VSS.n40 4.5005
R7229 VSS.n191 VSS.n40 4.5005
R7230 VSS.n197 VSS.n40 4.5005
R7231 VSS.n190 VSS.n40 4.5005
R7232 VSS.n198 VSS.n40 4.5005
R7233 VSS.n189 VSS.n40 4.5005
R7234 VSS.n199 VSS.n40 4.5005
R7235 VSS.n188 VSS.n40 4.5005
R7236 VSS.n200 VSS.n40 4.5005
R7237 VSS.n187 VSS.n40 4.5005
R7238 VSS.n201 VSS.n40 4.5005
R7239 VSS.n186 VSS.n40 4.5005
R7240 VSS.n202 VSS.n40 4.5005
R7241 VSS.n185 VSS.n40 4.5005
R7242 VSS.n203 VSS.n40 4.5005
R7243 VSS.n184 VSS.n40 4.5005
R7244 VSS.n204 VSS.n40 4.5005
R7245 VSS.n183 VSS.n40 4.5005
R7246 VSS.n205 VSS.n40 4.5005
R7247 VSS.n182 VSS.n40 4.5005
R7248 VSS.n206 VSS.n40 4.5005
R7249 VSS.n181 VSS.n40 4.5005
R7250 VSS.n207 VSS.n40 4.5005
R7251 VSS.n180 VSS.n40 4.5005
R7252 VSS.n208 VSS.n40 4.5005
R7253 VSS.n179 VSS.n40 4.5005
R7254 VSS.n209 VSS.n40 4.5005
R7255 VSS.n178 VSS.n40 4.5005
R7256 VSS.n210 VSS.n40 4.5005
R7257 VSS.n177 VSS.n40 4.5005
R7258 VSS.n211 VSS.n40 4.5005
R7259 VSS.n176 VSS.n40 4.5005
R7260 VSS.n212 VSS.n40 4.5005
R7261 VSS.n175 VSS.n40 4.5005
R7262 VSS.n213 VSS.n40 4.5005
R7263 VSS.n174 VSS.n40 4.5005
R7264 VSS.n214 VSS.n40 4.5005
R7265 VSS.n173 VSS.n40 4.5005
R7266 VSS.n215 VSS.n40 4.5005
R7267 VSS.n172 VSS.n40 4.5005
R7268 VSS.n216 VSS.n40 4.5005
R7269 VSS.n171 VSS.n40 4.5005
R7270 VSS.n217 VSS.n40 4.5005
R7271 VSS.n170 VSS.n40 4.5005
R7272 VSS.n218 VSS.n40 4.5005
R7273 VSS.n169 VSS.n40 4.5005
R7274 VSS.n219 VSS.n40 4.5005
R7275 VSS.n168 VSS.n40 4.5005
R7276 VSS.n220 VSS.n40 4.5005
R7277 VSS.n167 VSS.n40 4.5005
R7278 VSS.n221 VSS.n40 4.5005
R7279 VSS.n166 VSS.n40 4.5005
R7280 VSS.n222 VSS.n40 4.5005
R7281 VSS.n165 VSS.n40 4.5005
R7282 VSS.n223 VSS.n40 4.5005
R7283 VSS.n164 VSS.n40 4.5005
R7284 VSS.n224 VSS.n40 4.5005
R7285 VSS.n163 VSS.n40 4.5005
R7286 VSS.n225 VSS.n40 4.5005
R7287 VSS.n162 VSS.n40 4.5005
R7288 VSS.n226 VSS.n40 4.5005
R7289 VSS.n161 VSS.n40 4.5005
R7290 VSS.n227 VSS.n40 4.5005
R7291 VSS.n160 VSS.n40 4.5005
R7292 VSS.n228 VSS.n40 4.5005
R7293 VSS.n159 VSS.n40 4.5005
R7294 VSS.n229 VSS.n40 4.5005
R7295 VSS.n158 VSS.n40 4.5005
R7296 VSS.n230 VSS.n40 4.5005
R7297 VSS.n157 VSS.n40 4.5005
R7298 VSS.n231 VSS.n40 4.5005
R7299 VSS.n156 VSS.n40 4.5005
R7300 VSS.n232 VSS.n40 4.5005
R7301 VSS.n155 VSS.n40 4.5005
R7302 VSS.n233 VSS.n40 4.5005
R7303 VSS.n154 VSS.n40 4.5005
R7304 VSS.n234 VSS.n40 4.5005
R7305 VSS.n153 VSS.n40 4.5005
R7306 VSS.n235 VSS.n40 4.5005
R7307 VSS.n4506 VSS.n40 4.5005
R7308 VSS.n236 VSS.n40 4.5005
R7309 VSS.n152 VSS.n40 4.5005
R7310 VSS.n237 VSS.n40 4.5005
R7311 VSS.n151 VSS.n40 4.5005
R7312 VSS.n238 VSS.n40 4.5005
R7313 VSS.n150 VSS.n40 4.5005
R7314 VSS.n239 VSS.n40 4.5005
R7315 VSS.n149 VSS.n40 4.5005
R7316 VSS.n240 VSS.n40 4.5005
R7317 VSS.n148 VSS.n40 4.5005
R7318 VSS.n241 VSS.n40 4.5005
R7319 VSS.n147 VSS.n40 4.5005
R7320 VSS.n242 VSS.n40 4.5005
R7321 VSS.n146 VSS.n40 4.5005
R7322 VSS.n243 VSS.n40 4.5005
R7323 VSS.n145 VSS.n40 4.5005
R7324 VSS.n244 VSS.n40 4.5005
R7325 VSS.n144 VSS.n40 4.5005
R7326 VSS.n245 VSS.n40 4.5005
R7327 VSS.n143 VSS.n40 4.5005
R7328 VSS.n246 VSS.n40 4.5005
R7329 VSS.n142 VSS.n40 4.5005
R7330 VSS.n247 VSS.n40 4.5005
R7331 VSS.n141 VSS.n40 4.5005
R7332 VSS.n248 VSS.n40 4.5005
R7333 VSS.n140 VSS.n40 4.5005
R7334 VSS.n249 VSS.n40 4.5005
R7335 VSS.n139 VSS.n40 4.5005
R7336 VSS.n250 VSS.n40 4.5005
R7337 VSS.n138 VSS.n40 4.5005
R7338 VSS.n251 VSS.n40 4.5005
R7339 VSS.n137 VSS.n40 4.5005
R7340 VSS.n252 VSS.n40 4.5005
R7341 VSS.n136 VSS.n40 4.5005
R7342 VSS.n253 VSS.n40 4.5005
R7343 VSS.n135 VSS.n40 4.5005
R7344 VSS.n254 VSS.n40 4.5005
R7345 VSS.n134 VSS.n40 4.5005
R7346 VSS.n255 VSS.n40 4.5005
R7347 VSS.n133 VSS.n40 4.5005
R7348 VSS.n256 VSS.n40 4.5005
R7349 VSS.n132 VSS.n40 4.5005
R7350 VSS.n4502 VSS.n40 4.5005
R7351 VSS.n4504 VSS.n40 4.5005
R7352 VSS.n193 VSS.n97 4.5005
R7353 VSS.n195 VSS.n97 4.5005
R7354 VSS.n192 VSS.n97 4.5005
R7355 VSS.n196 VSS.n97 4.5005
R7356 VSS.n191 VSS.n97 4.5005
R7357 VSS.n197 VSS.n97 4.5005
R7358 VSS.n190 VSS.n97 4.5005
R7359 VSS.n198 VSS.n97 4.5005
R7360 VSS.n189 VSS.n97 4.5005
R7361 VSS.n199 VSS.n97 4.5005
R7362 VSS.n188 VSS.n97 4.5005
R7363 VSS.n200 VSS.n97 4.5005
R7364 VSS.n187 VSS.n97 4.5005
R7365 VSS.n201 VSS.n97 4.5005
R7366 VSS.n186 VSS.n97 4.5005
R7367 VSS.n202 VSS.n97 4.5005
R7368 VSS.n185 VSS.n97 4.5005
R7369 VSS.n203 VSS.n97 4.5005
R7370 VSS.n184 VSS.n97 4.5005
R7371 VSS.n204 VSS.n97 4.5005
R7372 VSS.n183 VSS.n97 4.5005
R7373 VSS.n205 VSS.n97 4.5005
R7374 VSS.n182 VSS.n97 4.5005
R7375 VSS.n206 VSS.n97 4.5005
R7376 VSS.n181 VSS.n97 4.5005
R7377 VSS.n207 VSS.n97 4.5005
R7378 VSS.n180 VSS.n97 4.5005
R7379 VSS.n208 VSS.n97 4.5005
R7380 VSS.n179 VSS.n97 4.5005
R7381 VSS.n209 VSS.n97 4.5005
R7382 VSS.n178 VSS.n97 4.5005
R7383 VSS.n210 VSS.n97 4.5005
R7384 VSS.n177 VSS.n97 4.5005
R7385 VSS.n211 VSS.n97 4.5005
R7386 VSS.n176 VSS.n97 4.5005
R7387 VSS.n212 VSS.n97 4.5005
R7388 VSS.n175 VSS.n97 4.5005
R7389 VSS.n213 VSS.n97 4.5005
R7390 VSS.n174 VSS.n97 4.5005
R7391 VSS.n214 VSS.n97 4.5005
R7392 VSS.n173 VSS.n97 4.5005
R7393 VSS.n215 VSS.n97 4.5005
R7394 VSS.n172 VSS.n97 4.5005
R7395 VSS.n216 VSS.n97 4.5005
R7396 VSS.n171 VSS.n97 4.5005
R7397 VSS.n217 VSS.n97 4.5005
R7398 VSS.n170 VSS.n97 4.5005
R7399 VSS.n218 VSS.n97 4.5005
R7400 VSS.n169 VSS.n97 4.5005
R7401 VSS.n219 VSS.n97 4.5005
R7402 VSS.n168 VSS.n97 4.5005
R7403 VSS.n220 VSS.n97 4.5005
R7404 VSS.n167 VSS.n97 4.5005
R7405 VSS.n221 VSS.n97 4.5005
R7406 VSS.n166 VSS.n97 4.5005
R7407 VSS.n222 VSS.n97 4.5005
R7408 VSS.n165 VSS.n97 4.5005
R7409 VSS.n223 VSS.n97 4.5005
R7410 VSS.n164 VSS.n97 4.5005
R7411 VSS.n224 VSS.n97 4.5005
R7412 VSS.n163 VSS.n97 4.5005
R7413 VSS.n225 VSS.n97 4.5005
R7414 VSS.n162 VSS.n97 4.5005
R7415 VSS.n226 VSS.n97 4.5005
R7416 VSS.n161 VSS.n97 4.5005
R7417 VSS.n227 VSS.n97 4.5005
R7418 VSS.n160 VSS.n97 4.5005
R7419 VSS.n228 VSS.n97 4.5005
R7420 VSS.n159 VSS.n97 4.5005
R7421 VSS.n229 VSS.n97 4.5005
R7422 VSS.n158 VSS.n97 4.5005
R7423 VSS.n230 VSS.n97 4.5005
R7424 VSS.n157 VSS.n97 4.5005
R7425 VSS.n231 VSS.n97 4.5005
R7426 VSS.n156 VSS.n97 4.5005
R7427 VSS.n232 VSS.n97 4.5005
R7428 VSS.n155 VSS.n97 4.5005
R7429 VSS.n233 VSS.n97 4.5005
R7430 VSS.n154 VSS.n97 4.5005
R7431 VSS.n234 VSS.n97 4.5005
R7432 VSS.n153 VSS.n97 4.5005
R7433 VSS.n235 VSS.n97 4.5005
R7434 VSS.n4506 VSS.n97 4.5005
R7435 VSS.n236 VSS.n97 4.5005
R7436 VSS.n152 VSS.n97 4.5005
R7437 VSS.n237 VSS.n97 4.5005
R7438 VSS.n151 VSS.n97 4.5005
R7439 VSS.n238 VSS.n97 4.5005
R7440 VSS.n150 VSS.n97 4.5005
R7441 VSS.n239 VSS.n97 4.5005
R7442 VSS.n149 VSS.n97 4.5005
R7443 VSS.n240 VSS.n97 4.5005
R7444 VSS.n148 VSS.n97 4.5005
R7445 VSS.n241 VSS.n97 4.5005
R7446 VSS.n147 VSS.n97 4.5005
R7447 VSS.n242 VSS.n97 4.5005
R7448 VSS.n146 VSS.n97 4.5005
R7449 VSS.n243 VSS.n97 4.5005
R7450 VSS.n145 VSS.n97 4.5005
R7451 VSS.n244 VSS.n97 4.5005
R7452 VSS.n144 VSS.n97 4.5005
R7453 VSS.n245 VSS.n97 4.5005
R7454 VSS.n143 VSS.n97 4.5005
R7455 VSS.n246 VSS.n97 4.5005
R7456 VSS.n142 VSS.n97 4.5005
R7457 VSS.n247 VSS.n97 4.5005
R7458 VSS.n141 VSS.n97 4.5005
R7459 VSS.n248 VSS.n97 4.5005
R7460 VSS.n140 VSS.n97 4.5005
R7461 VSS.n249 VSS.n97 4.5005
R7462 VSS.n139 VSS.n97 4.5005
R7463 VSS.n250 VSS.n97 4.5005
R7464 VSS.n138 VSS.n97 4.5005
R7465 VSS.n251 VSS.n97 4.5005
R7466 VSS.n137 VSS.n97 4.5005
R7467 VSS.n252 VSS.n97 4.5005
R7468 VSS.n136 VSS.n97 4.5005
R7469 VSS.n253 VSS.n97 4.5005
R7470 VSS.n135 VSS.n97 4.5005
R7471 VSS.n254 VSS.n97 4.5005
R7472 VSS.n134 VSS.n97 4.5005
R7473 VSS.n255 VSS.n97 4.5005
R7474 VSS.n133 VSS.n97 4.5005
R7475 VSS.n256 VSS.n97 4.5005
R7476 VSS.n132 VSS.n97 4.5005
R7477 VSS.n4502 VSS.n97 4.5005
R7478 VSS.n4504 VSS.n97 4.5005
R7479 VSS.n193 VSS.n39 4.5005
R7480 VSS.n195 VSS.n39 4.5005
R7481 VSS.n192 VSS.n39 4.5005
R7482 VSS.n196 VSS.n39 4.5005
R7483 VSS.n191 VSS.n39 4.5005
R7484 VSS.n197 VSS.n39 4.5005
R7485 VSS.n190 VSS.n39 4.5005
R7486 VSS.n198 VSS.n39 4.5005
R7487 VSS.n189 VSS.n39 4.5005
R7488 VSS.n199 VSS.n39 4.5005
R7489 VSS.n188 VSS.n39 4.5005
R7490 VSS.n200 VSS.n39 4.5005
R7491 VSS.n187 VSS.n39 4.5005
R7492 VSS.n201 VSS.n39 4.5005
R7493 VSS.n186 VSS.n39 4.5005
R7494 VSS.n202 VSS.n39 4.5005
R7495 VSS.n185 VSS.n39 4.5005
R7496 VSS.n203 VSS.n39 4.5005
R7497 VSS.n184 VSS.n39 4.5005
R7498 VSS.n204 VSS.n39 4.5005
R7499 VSS.n183 VSS.n39 4.5005
R7500 VSS.n205 VSS.n39 4.5005
R7501 VSS.n182 VSS.n39 4.5005
R7502 VSS.n206 VSS.n39 4.5005
R7503 VSS.n181 VSS.n39 4.5005
R7504 VSS.n207 VSS.n39 4.5005
R7505 VSS.n180 VSS.n39 4.5005
R7506 VSS.n208 VSS.n39 4.5005
R7507 VSS.n179 VSS.n39 4.5005
R7508 VSS.n209 VSS.n39 4.5005
R7509 VSS.n178 VSS.n39 4.5005
R7510 VSS.n210 VSS.n39 4.5005
R7511 VSS.n177 VSS.n39 4.5005
R7512 VSS.n211 VSS.n39 4.5005
R7513 VSS.n176 VSS.n39 4.5005
R7514 VSS.n212 VSS.n39 4.5005
R7515 VSS.n175 VSS.n39 4.5005
R7516 VSS.n213 VSS.n39 4.5005
R7517 VSS.n174 VSS.n39 4.5005
R7518 VSS.n214 VSS.n39 4.5005
R7519 VSS.n173 VSS.n39 4.5005
R7520 VSS.n215 VSS.n39 4.5005
R7521 VSS.n172 VSS.n39 4.5005
R7522 VSS.n216 VSS.n39 4.5005
R7523 VSS.n171 VSS.n39 4.5005
R7524 VSS.n217 VSS.n39 4.5005
R7525 VSS.n170 VSS.n39 4.5005
R7526 VSS.n218 VSS.n39 4.5005
R7527 VSS.n169 VSS.n39 4.5005
R7528 VSS.n219 VSS.n39 4.5005
R7529 VSS.n168 VSS.n39 4.5005
R7530 VSS.n220 VSS.n39 4.5005
R7531 VSS.n167 VSS.n39 4.5005
R7532 VSS.n221 VSS.n39 4.5005
R7533 VSS.n166 VSS.n39 4.5005
R7534 VSS.n222 VSS.n39 4.5005
R7535 VSS.n165 VSS.n39 4.5005
R7536 VSS.n223 VSS.n39 4.5005
R7537 VSS.n164 VSS.n39 4.5005
R7538 VSS.n224 VSS.n39 4.5005
R7539 VSS.n163 VSS.n39 4.5005
R7540 VSS.n225 VSS.n39 4.5005
R7541 VSS.n162 VSS.n39 4.5005
R7542 VSS.n226 VSS.n39 4.5005
R7543 VSS.n161 VSS.n39 4.5005
R7544 VSS.n227 VSS.n39 4.5005
R7545 VSS.n160 VSS.n39 4.5005
R7546 VSS.n228 VSS.n39 4.5005
R7547 VSS.n159 VSS.n39 4.5005
R7548 VSS.n229 VSS.n39 4.5005
R7549 VSS.n158 VSS.n39 4.5005
R7550 VSS.n230 VSS.n39 4.5005
R7551 VSS.n157 VSS.n39 4.5005
R7552 VSS.n231 VSS.n39 4.5005
R7553 VSS.n156 VSS.n39 4.5005
R7554 VSS.n232 VSS.n39 4.5005
R7555 VSS.n155 VSS.n39 4.5005
R7556 VSS.n233 VSS.n39 4.5005
R7557 VSS.n154 VSS.n39 4.5005
R7558 VSS.n234 VSS.n39 4.5005
R7559 VSS.n153 VSS.n39 4.5005
R7560 VSS.n235 VSS.n39 4.5005
R7561 VSS.n4506 VSS.n39 4.5005
R7562 VSS.n236 VSS.n39 4.5005
R7563 VSS.n152 VSS.n39 4.5005
R7564 VSS.n237 VSS.n39 4.5005
R7565 VSS.n151 VSS.n39 4.5005
R7566 VSS.n238 VSS.n39 4.5005
R7567 VSS.n150 VSS.n39 4.5005
R7568 VSS.n239 VSS.n39 4.5005
R7569 VSS.n149 VSS.n39 4.5005
R7570 VSS.n240 VSS.n39 4.5005
R7571 VSS.n148 VSS.n39 4.5005
R7572 VSS.n241 VSS.n39 4.5005
R7573 VSS.n147 VSS.n39 4.5005
R7574 VSS.n242 VSS.n39 4.5005
R7575 VSS.n146 VSS.n39 4.5005
R7576 VSS.n243 VSS.n39 4.5005
R7577 VSS.n145 VSS.n39 4.5005
R7578 VSS.n244 VSS.n39 4.5005
R7579 VSS.n144 VSS.n39 4.5005
R7580 VSS.n245 VSS.n39 4.5005
R7581 VSS.n143 VSS.n39 4.5005
R7582 VSS.n246 VSS.n39 4.5005
R7583 VSS.n142 VSS.n39 4.5005
R7584 VSS.n247 VSS.n39 4.5005
R7585 VSS.n141 VSS.n39 4.5005
R7586 VSS.n248 VSS.n39 4.5005
R7587 VSS.n140 VSS.n39 4.5005
R7588 VSS.n249 VSS.n39 4.5005
R7589 VSS.n139 VSS.n39 4.5005
R7590 VSS.n250 VSS.n39 4.5005
R7591 VSS.n138 VSS.n39 4.5005
R7592 VSS.n251 VSS.n39 4.5005
R7593 VSS.n137 VSS.n39 4.5005
R7594 VSS.n252 VSS.n39 4.5005
R7595 VSS.n136 VSS.n39 4.5005
R7596 VSS.n253 VSS.n39 4.5005
R7597 VSS.n135 VSS.n39 4.5005
R7598 VSS.n254 VSS.n39 4.5005
R7599 VSS.n134 VSS.n39 4.5005
R7600 VSS.n255 VSS.n39 4.5005
R7601 VSS.n133 VSS.n39 4.5005
R7602 VSS.n256 VSS.n39 4.5005
R7603 VSS.n132 VSS.n39 4.5005
R7604 VSS.n4502 VSS.n39 4.5005
R7605 VSS.n4504 VSS.n39 4.5005
R7606 VSS.n193 VSS.n98 4.5005
R7607 VSS.n195 VSS.n98 4.5005
R7608 VSS.n192 VSS.n98 4.5005
R7609 VSS.n196 VSS.n98 4.5005
R7610 VSS.n191 VSS.n98 4.5005
R7611 VSS.n197 VSS.n98 4.5005
R7612 VSS.n190 VSS.n98 4.5005
R7613 VSS.n198 VSS.n98 4.5005
R7614 VSS.n189 VSS.n98 4.5005
R7615 VSS.n199 VSS.n98 4.5005
R7616 VSS.n188 VSS.n98 4.5005
R7617 VSS.n200 VSS.n98 4.5005
R7618 VSS.n187 VSS.n98 4.5005
R7619 VSS.n201 VSS.n98 4.5005
R7620 VSS.n186 VSS.n98 4.5005
R7621 VSS.n202 VSS.n98 4.5005
R7622 VSS.n185 VSS.n98 4.5005
R7623 VSS.n203 VSS.n98 4.5005
R7624 VSS.n184 VSS.n98 4.5005
R7625 VSS.n204 VSS.n98 4.5005
R7626 VSS.n183 VSS.n98 4.5005
R7627 VSS.n205 VSS.n98 4.5005
R7628 VSS.n182 VSS.n98 4.5005
R7629 VSS.n206 VSS.n98 4.5005
R7630 VSS.n181 VSS.n98 4.5005
R7631 VSS.n207 VSS.n98 4.5005
R7632 VSS.n180 VSS.n98 4.5005
R7633 VSS.n208 VSS.n98 4.5005
R7634 VSS.n179 VSS.n98 4.5005
R7635 VSS.n209 VSS.n98 4.5005
R7636 VSS.n178 VSS.n98 4.5005
R7637 VSS.n210 VSS.n98 4.5005
R7638 VSS.n177 VSS.n98 4.5005
R7639 VSS.n211 VSS.n98 4.5005
R7640 VSS.n176 VSS.n98 4.5005
R7641 VSS.n212 VSS.n98 4.5005
R7642 VSS.n175 VSS.n98 4.5005
R7643 VSS.n213 VSS.n98 4.5005
R7644 VSS.n174 VSS.n98 4.5005
R7645 VSS.n214 VSS.n98 4.5005
R7646 VSS.n173 VSS.n98 4.5005
R7647 VSS.n215 VSS.n98 4.5005
R7648 VSS.n172 VSS.n98 4.5005
R7649 VSS.n216 VSS.n98 4.5005
R7650 VSS.n171 VSS.n98 4.5005
R7651 VSS.n217 VSS.n98 4.5005
R7652 VSS.n170 VSS.n98 4.5005
R7653 VSS.n218 VSS.n98 4.5005
R7654 VSS.n169 VSS.n98 4.5005
R7655 VSS.n219 VSS.n98 4.5005
R7656 VSS.n168 VSS.n98 4.5005
R7657 VSS.n220 VSS.n98 4.5005
R7658 VSS.n167 VSS.n98 4.5005
R7659 VSS.n221 VSS.n98 4.5005
R7660 VSS.n166 VSS.n98 4.5005
R7661 VSS.n222 VSS.n98 4.5005
R7662 VSS.n165 VSS.n98 4.5005
R7663 VSS.n223 VSS.n98 4.5005
R7664 VSS.n164 VSS.n98 4.5005
R7665 VSS.n224 VSS.n98 4.5005
R7666 VSS.n163 VSS.n98 4.5005
R7667 VSS.n225 VSS.n98 4.5005
R7668 VSS.n162 VSS.n98 4.5005
R7669 VSS.n226 VSS.n98 4.5005
R7670 VSS.n161 VSS.n98 4.5005
R7671 VSS.n227 VSS.n98 4.5005
R7672 VSS.n160 VSS.n98 4.5005
R7673 VSS.n228 VSS.n98 4.5005
R7674 VSS.n159 VSS.n98 4.5005
R7675 VSS.n229 VSS.n98 4.5005
R7676 VSS.n158 VSS.n98 4.5005
R7677 VSS.n230 VSS.n98 4.5005
R7678 VSS.n157 VSS.n98 4.5005
R7679 VSS.n231 VSS.n98 4.5005
R7680 VSS.n156 VSS.n98 4.5005
R7681 VSS.n232 VSS.n98 4.5005
R7682 VSS.n155 VSS.n98 4.5005
R7683 VSS.n233 VSS.n98 4.5005
R7684 VSS.n154 VSS.n98 4.5005
R7685 VSS.n234 VSS.n98 4.5005
R7686 VSS.n153 VSS.n98 4.5005
R7687 VSS.n235 VSS.n98 4.5005
R7688 VSS.n4506 VSS.n98 4.5005
R7689 VSS.n236 VSS.n98 4.5005
R7690 VSS.n152 VSS.n98 4.5005
R7691 VSS.n237 VSS.n98 4.5005
R7692 VSS.n151 VSS.n98 4.5005
R7693 VSS.n238 VSS.n98 4.5005
R7694 VSS.n150 VSS.n98 4.5005
R7695 VSS.n239 VSS.n98 4.5005
R7696 VSS.n149 VSS.n98 4.5005
R7697 VSS.n240 VSS.n98 4.5005
R7698 VSS.n148 VSS.n98 4.5005
R7699 VSS.n241 VSS.n98 4.5005
R7700 VSS.n147 VSS.n98 4.5005
R7701 VSS.n242 VSS.n98 4.5005
R7702 VSS.n146 VSS.n98 4.5005
R7703 VSS.n243 VSS.n98 4.5005
R7704 VSS.n145 VSS.n98 4.5005
R7705 VSS.n244 VSS.n98 4.5005
R7706 VSS.n144 VSS.n98 4.5005
R7707 VSS.n245 VSS.n98 4.5005
R7708 VSS.n143 VSS.n98 4.5005
R7709 VSS.n246 VSS.n98 4.5005
R7710 VSS.n142 VSS.n98 4.5005
R7711 VSS.n247 VSS.n98 4.5005
R7712 VSS.n141 VSS.n98 4.5005
R7713 VSS.n248 VSS.n98 4.5005
R7714 VSS.n140 VSS.n98 4.5005
R7715 VSS.n249 VSS.n98 4.5005
R7716 VSS.n139 VSS.n98 4.5005
R7717 VSS.n250 VSS.n98 4.5005
R7718 VSS.n138 VSS.n98 4.5005
R7719 VSS.n251 VSS.n98 4.5005
R7720 VSS.n137 VSS.n98 4.5005
R7721 VSS.n252 VSS.n98 4.5005
R7722 VSS.n136 VSS.n98 4.5005
R7723 VSS.n253 VSS.n98 4.5005
R7724 VSS.n135 VSS.n98 4.5005
R7725 VSS.n254 VSS.n98 4.5005
R7726 VSS.n134 VSS.n98 4.5005
R7727 VSS.n255 VSS.n98 4.5005
R7728 VSS.n133 VSS.n98 4.5005
R7729 VSS.n256 VSS.n98 4.5005
R7730 VSS.n132 VSS.n98 4.5005
R7731 VSS.n4502 VSS.n98 4.5005
R7732 VSS.n4504 VSS.n98 4.5005
R7733 VSS.n193 VSS.n38 4.5005
R7734 VSS.n195 VSS.n38 4.5005
R7735 VSS.n192 VSS.n38 4.5005
R7736 VSS.n196 VSS.n38 4.5005
R7737 VSS.n191 VSS.n38 4.5005
R7738 VSS.n197 VSS.n38 4.5005
R7739 VSS.n190 VSS.n38 4.5005
R7740 VSS.n198 VSS.n38 4.5005
R7741 VSS.n189 VSS.n38 4.5005
R7742 VSS.n199 VSS.n38 4.5005
R7743 VSS.n188 VSS.n38 4.5005
R7744 VSS.n200 VSS.n38 4.5005
R7745 VSS.n187 VSS.n38 4.5005
R7746 VSS.n201 VSS.n38 4.5005
R7747 VSS.n186 VSS.n38 4.5005
R7748 VSS.n202 VSS.n38 4.5005
R7749 VSS.n185 VSS.n38 4.5005
R7750 VSS.n203 VSS.n38 4.5005
R7751 VSS.n184 VSS.n38 4.5005
R7752 VSS.n204 VSS.n38 4.5005
R7753 VSS.n183 VSS.n38 4.5005
R7754 VSS.n205 VSS.n38 4.5005
R7755 VSS.n182 VSS.n38 4.5005
R7756 VSS.n206 VSS.n38 4.5005
R7757 VSS.n181 VSS.n38 4.5005
R7758 VSS.n207 VSS.n38 4.5005
R7759 VSS.n180 VSS.n38 4.5005
R7760 VSS.n208 VSS.n38 4.5005
R7761 VSS.n179 VSS.n38 4.5005
R7762 VSS.n209 VSS.n38 4.5005
R7763 VSS.n178 VSS.n38 4.5005
R7764 VSS.n210 VSS.n38 4.5005
R7765 VSS.n177 VSS.n38 4.5005
R7766 VSS.n211 VSS.n38 4.5005
R7767 VSS.n176 VSS.n38 4.5005
R7768 VSS.n212 VSS.n38 4.5005
R7769 VSS.n175 VSS.n38 4.5005
R7770 VSS.n213 VSS.n38 4.5005
R7771 VSS.n174 VSS.n38 4.5005
R7772 VSS.n214 VSS.n38 4.5005
R7773 VSS.n173 VSS.n38 4.5005
R7774 VSS.n215 VSS.n38 4.5005
R7775 VSS.n172 VSS.n38 4.5005
R7776 VSS.n216 VSS.n38 4.5005
R7777 VSS.n171 VSS.n38 4.5005
R7778 VSS.n217 VSS.n38 4.5005
R7779 VSS.n170 VSS.n38 4.5005
R7780 VSS.n218 VSS.n38 4.5005
R7781 VSS.n169 VSS.n38 4.5005
R7782 VSS.n219 VSS.n38 4.5005
R7783 VSS.n168 VSS.n38 4.5005
R7784 VSS.n220 VSS.n38 4.5005
R7785 VSS.n167 VSS.n38 4.5005
R7786 VSS.n221 VSS.n38 4.5005
R7787 VSS.n166 VSS.n38 4.5005
R7788 VSS.n222 VSS.n38 4.5005
R7789 VSS.n165 VSS.n38 4.5005
R7790 VSS.n223 VSS.n38 4.5005
R7791 VSS.n164 VSS.n38 4.5005
R7792 VSS.n224 VSS.n38 4.5005
R7793 VSS.n163 VSS.n38 4.5005
R7794 VSS.n225 VSS.n38 4.5005
R7795 VSS.n162 VSS.n38 4.5005
R7796 VSS.n226 VSS.n38 4.5005
R7797 VSS.n161 VSS.n38 4.5005
R7798 VSS.n227 VSS.n38 4.5005
R7799 VSS.n160 VSS.n38 4.5005
R7800 VSS.n228 VSS.n38 4.5005
R7801 VSS.n159 VSS.n38 4.5005
R7802 VSS.n229 VSS.n38 4.5005
R7803 VSS.n158 VSS.n38 4.5005
R7804 VSS.n230 VSS.n38 4.5005
R7805 VSS.n157 VSS.n38 4.5005
R7806 VSS.n231 VSS.n38 4.5005
R7807 VSS.n156 VSS.n38 4.5005
R7808 VSS.n232 VSS.n38 4.5005
R7809 VSS.n155 VSS.n38 4.5005
R7810 VSS.n233 VSS.n38 4.5005
R7811 VSS.n154 VSS.n38 4.5005
R7812 VSS.n234 VSS.n38 4.5005
R7813 VSS.n153 VSS.n38 4.5005
R7814 VSS.n235 VSS.n38 4.5005
R7815 VSS.n4506 VSS.n38 4.5005
R7816 VSS.n236 VSS.n38 4.5005
R7817 VSS.n152 VSS.n38 4.5005
R7818 VSS.n237 VSS.n38 4.5005
R7819 VSS.n151 VSS.n38 4.5005
R7820 VSS.n238 VSS.n38 4.5005
R7821 VSS.n150 VSS.n38 4.5005
R7822 VSS.n239 VSS.n38 4.5005
R7823 VSS.n149 VSS.n38 4.5005
R7824 VSS.n240 VSS.n38 4.5005
R7825 VSS.n148 VSS.n38 4.5005
R7826 VSS.n241 VSS.n38 4.5005
R7827 VSS.n147 VSS.n38 4.5005
R7828 VSS.n242 VSS.n38 4.5005
R7829 VSS.n146 VSS.n38 4.5005
R7830 VSS.n243 VSS.n38 4.5005
R7831 VSS.n145 VSS.n38 4.5005
R7832 VSS.n244 VSS.n38 4.5005
R7833 VSS.n144 VSS.n38 4.5005
R7834 VSS.n245 VSS.n38 4.5005
R7835 VSS.n143 VSS.n38 4.5005
R7836 VSS.n246 VSS.n38 4.5005
R7837 VSS.n142 VSS.n38 4.5005
R7838 VSS.n247 VSS.n38 4.5005
R7839 VSS.n141 VSS.n38 4.5005
R7840 VSS.n248 VSS.n38 4.5005
R7841 VSS.n140 VSS.n38 4.5005
R7842 VSS.n249 VSS.n38 4.5005
R7843 VSS.n139 VSS.n38 4.5005
R7844 VSS.n250 VSS.n38 4.5005
R7845 VSS.n138 VSS.n38 4.5005
R7846 VSS.n251 VSS.n38 4.5005
R7847 VSS.n137 VSS.n38 4.5005
R7848 VSS.n252 VSS.n38 4.5005
R7849 VSS.n136 VSS.n38 4.5005
R7850 VSS.n253 VSS.n38 4.5005
R7851 VSS.n135 VSS.n38 4.5005
R7852 VSS.n254 VSS.n38 4.5005
R7853 VSS.n134 VSS.n38 4.5005
R7854 VSS.n255 VSS.n38 4.5005
R7855 VSS.n133 VSS.n38 4.5005
R7856 VSS.n256 VSS.n38 4.5005
R7857 VSS.n132 VSS.n38 4.5005
R7858 VSS.n4502 VSS.n38 4.5005
R7859 VSS.n4504 VSS.n38 4.5005
R7860 VSS.n193 VSS.n99 4.5005
R7861 VSS.n195 VSS.n99 4.5005
R7862 VSS.n192 VSS.n99 4.5005
R7863 VSS.n196 VSS.n99 4.5005
R7864 VSS.n191 VSS.n99 4.5005
R7865 VSS.n197 VSS.n99 4.5005
R7866 VSS.n190 VSS.n99 4.5005
R7867 VSS.n198 VSS.n99 4.5005
R7868 VSS.n189 VSS.n99 4.5005
R7869 VSS.n199 VSS.n99 4.5005
R7870 VSS.n188 VSS.n99 4.5005
R7871 VSS.n200 VSS.n99 4.5005
R7872 VSS.n187 VSS.n99 4.5005
R7873 VSS.n201 VSS.n99 4.5005
R7874 VSS.n186 VSS.n99 4.5005
R7875 VSS.n202 VSS.n99 4.5005
R7876 VSS.n185 VSS.n99 4.5005
R7877 VSS.n203 VSS.n99 4.5005
R7878 VSS.n184 VSS.n99 4.5005
R7879 VSS.n204 VSS.n99 4.5005
R7880 VSS.n183 VSS.n99 4.5005
R7881 VSS.n205 VSS.n99 4.5005
R7882 VSS.n182 VSS.n99 4.5005
R7883 VSS.n206 VSS.n99 4.5005
R7884 VSS.n181 VSS.n99 4.5005
R7885 VSS.n207 VSS.n99 4.5005
R7886 VSS.n180 VSS.n99 4.5005
R7887 VSS.n208 VSS.n99 4.5005
R7888 VSS.n179 VSS.n99 4.5005
R7889 VSS.n209 VSS.n99 4.5005
R7890 VSS.n178 VSS.n99 4.5005
R7891 VSS.n210 VSS.n99 4.5005
R7892 VSS.n177 VSS.n99 4.5005
R7893 VSS.n211 VSS.n99 4.5005
R7894 VSS.n176 VSS.n99 4.5005
R7895 VSS.n212 VSS.n99 4.5005
R7896 VSS.n175 VSS.n99 4.5005
R7897 VSS.n213 VSS.n99 4.5005
R7898 VSS.n174 VSS.n99 4.5005
R7899 VSS.n214 VSS.n99 4.5005
R7900 VSS.n173 VSS.n99 4.5005
R7901 VSS.n215 VSS.n99 4.5005
R7902 VSS.n172 VSS.n99 4.5005
R7903 VSS.n216 VSS.n99 4.5005
R7904 VSS.n171 VSS.n99 4.5005
R7905 VSS.n217 VSS.n99 4.5005
R7906 VSS.n170 VSS.n99 4.5005
R7907 VSS.n218 VSS.n99 4.5005
R7908 VSS.n169 VSS.n99 4.5005
R7909 VSS.n219 VSS.n99 4.5005
R7910 VSS.n168 VSS.n99 4.5005
R7911 VSS.n220 VSS.n99 4.5005
R7912 VSS.n167 VSS.n99 4.5005
R7913 VSS.n221 VSS.n99 4.5005
R7914 VSS.n166 VSS.n99 4.5005
R7915 VSS.n222 VSS.n99 4.5005
R7916 VSS.n165 VSS.n99 4.5005
R7917 VSS.n223 VSS.n99 4.5005
R7918 VSS.n164 VSS.n99 4.5005
R7919 VSS.n224 VSS.n99 4.5005
R7920 VSS.n163 VSS.n99 4.5005
R7921 VSS.n225 VSS.n99 4.5005
R7922 VSS.n162 VSS.n99 4.5005
R7923 VSS.n226 VSS.n99 4.5005
R7924 VSS.n161 VSS.n99 4.5005
R7925 VSS.n227 VSS.n99 4.5005
R7926 VSS.n160 VSS.n99 4.5005
R7927 VSS.n228 VSS.n99 4.5005
R7928 VSS.n159 VSS.n99 4.5005
R7929 VSS.n229 VSS.n99 4.5005
R7930 VSS.n158 VSS.n99 4.5005
R7931 VSS.n230 VSS.n99 4.5005
R7932 VSS.n157 VSS.n99 4.5005
R7933 VSS.n231 VSS.n99 4.5005
R7934 VSS.n156 VSS.n99 4.5005
R7935 VSS.n232 VSS.n99 4.5005
R7936 VSS.n155 VSS.n99 4.5005
R7937 VSS.n233 VSS.n99 4.5005
R7938 VSS.n154 VSS.n99 4.5005
R7939 VSS.n234 VSS.n99 4.5005
R7940 VSS.n153 VSS.n99 4.5005
R7941 VSS.n235 VSS.n99 4.5005
R7942 VSS.n4506 VSS.n99 4.5005
R7943 VSS.n236 VSS.n99 4.5005
R7944 VSS.n152 VSS.n99 4.5005
R7945 VSS.n237 VSS.n99 4.5005
R7946 VSS.n151 VSS.n99 4.5005
R7947 VSS.n238 VSS.n99 4.5005
R7948 VSS.n150 VSS.n99 4.5005
R7949 VSS.n239 VSS.n99 4.5005
R7950 VSS.n149 VSS.n99 4.5005
R7951 VSS.n240 VSS.n99 4.5005
R7952 VSS.n148 VSS.n99 4.5005
R7953 VSS.n241 VSS.n99 4.5005
R7954 VSS.n147 VSS.n99 4.5005
R7955 VSS.n242 VSS.n99 4.5005
R7956 VSS.n146 VSS.n99 4.5005
R7957 VSS.n243 VSS.n99 4.5005
R7958 VSS.n145 VSS.n99 4.5005
R7959 VSS.n244 VSS.n99 4.5005
R7960 VSS.n144 VSS.n99 4.5005
R7961 VSS.n245 VSS.n99 4.5005
R7962 VSS.n143 VSS.n99 4.5005
R7963 VSS.n246 VSS.n99 4.5005
R7964 VSS.n142 VSS.n99 4.5005
R7965 VSS.n247 VSS.n99 4.5005
R7966 VSS.n141 VSS.n99 4.5005
R7967 VSS.n248 VSS.n99 4.5005
R7968 VSS.n140 VSS.n99 4.5005
R7969 VSS.n249 VSS.n99 4.5005
R7970 VSS.n139 VSS.n99 4.5005
R7971 VSS.n250 VSS.n99 4.5005
R7972 VSS.n138 VSS.n99 4.5005
R7973 VSS.n251 VSS.n99 4.5005
R7974 VSS.n137 VSS.n99 4.5005
R7975 VSS.n252 VSS.n99 4.5005
R7976 VSS.n136 VSS.n99 4.5005
R7977 VSS.n253 VSS.n99 4.5005
R7978 VSS.n135 VSS.n99 4.5005
R7979 VSS.n254 VSS.n99 4.5005
R7980 VSS.n134 VSS.n99 4.5005
R7981 VSS.n255 VSS.n99 4.5005
R7982 VSS.n133 VSS.n99 4.5005
R7983 VSS.n256 VSS.n99 4.5005
R7984 VSS.n132 VSS.n99 4.5005
R7985 VSS.n4502 VSS.n99 4.5005
R7986 VSS.n4504 VSS.n99 4.5005
R7987 VSS.n193 VSS.n37 4.5005
R7988 VSS.n195 VSS.n37 4.5005
R7989 VSS.n192 VSS.n37 4.5005
R7990 VSS.n196 VSS.n37 4.5005
R7991 VSS.n191 VSS.n37 4.5005
R7992 VSS.n197 VSS.n37 4.5005
R7993 VSS.n190 VSS.n37 4.5005
R7994 VSS.n198 VSS.n37 4.5005
R7995 VSS.n189 VSS.n37 4.5005
R7996 VSS.n199 VSS.n37 4.5005
R7997 VSS.n188 VSS.n37 4.5005
R7998 VSS.n200 VSS.n37 4.5005
R7999 VSS.n187 VSS.n37 4.5005
R8000 VSS.n201 VSS.n37 4.5005
R8001 VSS.n186 VSS.n37 4.5005
R8002 VSS.n202 VSS.n37 4.5005
R8003 VSS.n185 VSS.n37 4.5005
R8004 VSS.n203 VSS.n37 4.5005
R8005 VSS.n184 VSS.n37 4.5005
R8006 VSS.n204 VSS.n37 4.5005
R8007 VSS.n183 VSS.n37 4.5005
R8008 VSS.n205 VSS.n37 4.5005
R8009 VSS.n182 VSS.n37 4.5005
R8010 VSS.n206 VSS.n37 4.5005
R8011 VSS.n181 VSS.n37 4.5005
R8012 VSS.n207 VSS.n37 4.5005
R8013 VSS.n180 VSS.n37 4.5005
R8014 VSS.n208 VSS.n37 4.5005
R8015 VSS.n179 VSS.n37 4.5005
R8016 VSS.n209 VSS.n37 4.5005
R8017 VSS.n178 VSS.n37 4.5005
R8018 VSS.n210 VSS.n37 4.5005
R8019 VSS.n177 VSS.n37 4.5005
R8020 VSS.n211 VSS.n37 4.5005
R8021 VSS.n176 VSS.n37 4.5005
R8022 VSS.n212 VSS.n37 4.5005
R8023 VSS.n175 VSS.n37 4.5005
R8024 VSS.n213 VSS.n37 4.5005
R8025 VSS.n174 VSS.n37 4.5005
R8026 VSS.n214 VSS.n37 4.5005
R8027 VSS.n173 VSS.n37 4.5005
R8028 VSS.n215 VSS.n37 4.5005
R8029 VSS.n172 VSS.n37 4.5005
R8030 VSS.n216 VSS.n37 4.5005
R8031 VSS.n171 VSS.n37 4.5005
R8032 VSS.n217 VSS.n37 4.5005
R8033 VSS.n170 VSS.n37 4.5005
R8034 VSS.n218 VSS.n37 4.5005
R8035 VSS.n169 VSS.n37 4.5005
R8036 VSS.n219 VSS.n37 4.5005
R8037 VSS.n168 VSS.n37 4.5005
R8038 VSS.n220 VSS.n37 4.5005
R8039 VSS.n167 VSS.n37 4.5005
R8040 VSS.n221 VSS.n37 4.5005
R8041 VSS.n166 VSS.n37 4.5005
R8042 VSS.n222 VSS.n37 4.5005
R8043 VSS.n165 VSS.n37 4.5005
R8044 VSS.n223 VSS.n37 4.5005
R8045 VSS.n164 VSS.n37 4.5005
R8046 VSS.n224 VSS.n37 4.5005
R8047 VSS.n163 VSS.n37 4.5005
R8048 VSS.n225 VSS.n37 4.5005
R8049 VSS.n162 VSS.n37 4.5005
R8050 VSS.n226 VSS.n37 4.5005
R8051 VSS.n161 VSS.n37 4.5005
R8052 VSS.n227 VSS.n37 4.5005
R8053 VSS.n160 VSS.n37 4.5005
R8054 VSS.n228 VSS.n37 4.5005
R8055 VSS.n159 VSS.n37 4.5005
R8056 VSS.n229 VSS.n37 4.5005
R8057 VSS.n158 VSS.n37 4.5005
R8058 VSS.n230 VSS.n37 4.5005
R8059 VSS.n157 VSS.n37 4.5005
R8060 VSS.n231 VSS.n37 4.5005
R8061 VSS.n156 VSS.n37 4.5005
R8062 VSS.n232 VSS.n37 4.5005
R8063 VSS.n155 VSS.n37 4.5005
R8064 VSS.n233 VSS.n37 4.5005
R8065 VSS.n154 VSS.n37 4.5005
R8066 VSS.n234 VSS.n37 4.5005
R8067 VSS.n153 VSS.n37 4.5005
R8068 VSS.n235 VSS.n37 4.5005
R8069 VSS.n4506 VSS.n37 4.5005
R8070 VSS.n236 VSS.n37 4.5005
R8071 VSS.n152 VSS.n37 4.5005
R8072 VSS.n237 VSS.n37 4.5005
R8073 VSS.n151 VSS.n37 4.5005
R8074 VSS.n238 VSS.n37 4.5005
R8075 VSS.n150 VSS.n37 4.5005
R8076 VSS.n239 VSS.n37 4.5005
R8077 VSS.n149 VSS.n37 4.5005
R8078 VSS.n240 VSS.n37 4.5005
R8079 VSS.n148 VSS.n37 4.5005
R8080 VSS.n241 VSS.n37 4.5005
R8081 VSS.n147 VSS.n37 4.5005
R8082 VSS.n242 VSS.n37 4.5005
R8083 VSS.n146 VSS.n37 4.5005
R8084 VSS.n243 VSS.n37 4.5005
R8085 VSS.n145 VSS.n37 4.5005
R8086 VSS.n244 VSS.n37 4.5005
R8087 VSS.n144 VSS.n37 4.5005
R8088 VSS.n245 VSS.n37 4.5005
R8089 VSS.n143 VSS.n37 4.5005
R8090 VSS.n246 VSS.n37 4.5005
R8091 VSS.n142 VSS.n37 4.5005
R8092 VSS.n247 VSS.n37 4.5005
R8093 VSS.n141 VSS.n37 4.5005
R8094 VSS.n248 VSS.n37 4.5005
R8095 VSS.n140 VSS.n37 4.5005
R8096 VSS.n249 VSS.n37 4.5005
R8097 VSS.n139 VSS.n37 4.5005
R8098 VSS.n250 VSS.n37 4.5005
R8099 VSS.n138 VSS.n37 4.5005
R8100 VSS.n251 VSS.n37 4.5005
R8101 VSS.n137 VSS.n37 4.5005
R8102 VSS.n252 VSS.n37 4.5005
R8103 VSS.n136 VSS.n37 4.5005
R8104 VSS.n253 VSS.n37 4.5005
R8105 VSS.n135 VSS.n37 4.5005
R8106 VSS.n254 VSS.n37 4.5005
R8107 VSS.n134 VSS.n37 4.5005
R8108 VSS.n255 VSS.n37 4.5005
R8109 VSS.n133 VSS.n37 4.5005
R8110 VSS.n256 VSS.n37 4.5005
R8111 VSS.n132 VSS.n37 4.5005
R8112 VSS.n4502 VSS.n37 4.5005
R8113 VSS.n4504 VSS.n37 4.5005
R8114 VSS.n193 VSS.n100 4.5005
R8115 VSS.n195 VSS.n100 4.5005
R8116 VSS.n192 VSS.n100 4.5005
R8117 VSS.n196 VSS.n100 4.5005
R8118 VSS.n191 VSS.n100 4.5005
R8119 VSS.n197 VSS.n100 4.5005
R8120 VSS.n190 VSS.n100 4.5005
R8121 VSS.n198 VSS.n100 4.5005
R8122 VSS.n189 VSS.n100 4.5005
R8123 VSS.n199 VSS.n100 4.5005
R8124 VSS.n188 VSS.n100 4.5005
R8125 VSS.n200 VSS.n100 4.5005
R8126 VSS.n187 VSS.n100 4.5005
R8127 VSS.n201 VSS.n100 4.5005
R8128 VSS.n186 VSS.n100 4.5005
R8129 VSS.n202 VSS.n100 4.5005
R8130 VSS.n185 VSS.n100 4.5005
R8131 VSS.n203 VSS.n100 4.5005
R8132 VSS.n184 VSS.n100 4.5005
R8133 VSS.n204 VSS.n100 4.5005
R8134 VSS.n183 VSS.n100 4.5005
R8135 VSS.n205 VSS.n100 4.5005
R8136 VSS.n182 VSS.n100 4.5005
R8137 VSS.n206 VSS.n100 4.5005
R8138 VSS.n181 VSS.n100 4.5005
R8139 VSS.n207 VSS.n100 4.5005
R8140 VSS.n180 VSS.n100 4.5005
R8141 VSS.n208 VSS.n100 4.5005
R8142 VSS.n179 VSS.n100 4.5005
R8143 VSS.n209 VSS.n100 4.5005
R8144 VSS.n178 VSS.n100 4.5005
R8145 VSS.n210 VSS.n100 4.5005
R8146 VSS.n177 VSS.n100 4.5005
R8147 VSS.n211 VSS.n100 4.5005
R8148 VSS.n176 VSS.n100 4.5005
R8149 VSS.n212 VSS.n100 4.5005
R8150 VSS.n175 VSS.n100 4.5005
R8151 VSS.n213 VSS.n100 4.5005
R8152 VSS.n174 VSS.n100 4.5005
R8153 VSS.n214 VSS.n100 4.5005
R8154 VSS.n173 VSS.n100 4.5005
R8155 VSS.n215 VSS.n100 4.5005
R8156 VSS.n172 VSS.n100 4.5005
R8157 VSS.n216 VSS.n100 4.5005
R8158 VSS.n171 VSS.n100 4.5005
R8159 VSS.n217 VSS.n100 4.5005
R8160 VSS.n170 VSS.n100 4.5005
R8161 VSS.n218 VSS.n100 4.5005
R8162 VSS.n169 VSS.n100 4.5005
R8163 VSS.n219 VSS.n100 4.5005
R8164 VSS.n168 VSS.n100 4.5005
R8165 VSS.n220 VSS.n100 4.5005
R8166 VSS.n167 VSS.n100 4.5005
R8167 VSS.n221 VSS.n100 4.5005
R8168 VSS.n166 VSS.n100 4.5005
R8169 VSS.n222 VSS.n100 4.5005
R8170 VSS.n165 VSS.n100 4.5005
R8171 VSS.n223 VSS.n100 4.5005
R8172 VSS.n164 VSS.n100 4.5005
R8173 VSS.n224 VSS.n100 4.5005
R8174 VSS.n163 VSS.n100 4.5005
R8175 VSS.n225 VSS.n100 4.5005
R8176 VSS.n162 VSS.n100 4.5005
R8177 VSS.n226 VSS.n100 4.5005
R8178 VSS.n161 VSS.n100 4.5005
R8179 VSS.n227 VSS.n100 4.5005
R8180 VSS.n160 VSS.n100 4.5005
R8181 VSS.n228 VSS.n100 4.5005
R8182 VSS.n159 VSS.n100 4.5005
R8183 VSS.n229 VSS.n100 4.5005
R8184 VSS.n158 VSS.n100 4.5005
R8185 VSS.n230 VSS.n100 4.5005
R8186 VSS.n157 VSS.n100 4.5005
R8187 VSS.n231 VSS.n100 4.5005
R8188 VSS.n156 VSS.n100 4.5005
R8189 VSS.n232 VSS.n100 4.5005
R8190 VSS.n155 VSS.n100 4.5005
R8191 VSS.n233 VSS.n100 4.5005
R8192 VSS.n154 VSS.n100 4.5005
R8193 VSS.n234 VSS.n100 4.5005
R8194 VSS.n153 VSS.n100 4.5005
R8195 VSS.n235 VSS.n100 4.5005
R8196 VSS.n4506 VSS.n100 4.5005
R8197 VSS.n236 VSS.n100 4.5005
R8198 VSS.n152 VSS.n100 4.5005
R8199 VSS.n237 VSS.n100 4.5005
R8200 VSS.n151 VSS.n100 4.5005
R8201 VSS.n238 VSS.n100 4.5005
R8202 VSS.n150 VSS.n100 4.5005
R8203 VSS.n239 VSS.n100 4.5005
R8204 VSS.n149 VSS.n100 4.5005
R8205 VSS.n240 VSS.n100 4.5005
R8206 VSS.n148 VSS.n100 4.5005
R8207 VSS.n241 VSS.n100 4.5005
R8208 VSS.n147 VSS.n100 4.5005
R8209 VSS.n242 VSS.n100 4.5005
R8210 VSS.n146 VSS.n100 4.5005
R8211 VSS.n243 VSS.n100 4.5005
R8212 VSS.n145 VSS.n100 4.5005
R8213 VSS.n244 VSS.n100 4.5005
R8214 VSS.n144 VSS.n100 4.5005
R8215 VSS.n245 VSS.n100 4.5005
R8216 VSS.n143 VSS.n100 4.5005
R8217 VSS.n246 VSS.n100 4.5005
R8218 VSS.n142 VSS.n100 4.5005
R8219 VSS.n247 VSS.n100 4.5005
R8220 VSS.n141 VSS.n100 4.5005
R8221 VSS.n248 VSS.n100 4.5005
R8222 VSS.n140 VSS.n100 4.5005
R8223 VSS.n249 VSS.n100 4.5005
R8224 VSS.n139 VSS.n100 4.5005
R8225 VSS.n250 VSS.n100 4.5005
R8226 VSS.n138 VSS.n100 4.5005
R8227 VSS.n251 VSS.n100 4.5005
R8228 VSS.n137 VSS.n100 4.5005
R8229 VSS.n252 VSS.n100 4.5005
R8230 VSS.n136 VSS.n100 4.5005
R8231 VSS.n253 VSS.n100 4.5005
R8232 VSS.n135 VSS.n100 4.5005
R8233 VSS.n254 VSS.n100 4.5005
R8234 VSS.n134 VSS.n100 4.5005
R8235 VSS.n255 VSS.n100 4.5005
R8236 VSS.n133 VSS.n100 4.5005
R8237 VSS.n256 VSS.n100 4.5005
R8238 VSS.n132 VSS.n100 4.5005
R8239 VSS.n4502 VSS.n100 4.5005
R8240 VSS.n4504 VSS.n100 4.5005
R8241 VSS.n193 VSS.n36 4.5005
R8242 VSS.n195 VSS.n36 4.5005
R8243 VSS.n192 VSS.n36 4.5005
R8244 VSS.n196 VSS.n36 4.5005
R8245 VSS.n191 VSS.n36 4.5005
R8246 VSS.n197 VSS.n36 4.5005
R8247 VSS.n190 VSS.n36 4.5005
R8248 VSS.n198 VSS.n36 4.5005
R8249 VSS.n189 VSS.n36 4.5005
R8250 VSS.n199 VSS.n36 4.5005
R8251 VSS.n188 VSS.n36 4.5005
R8252 VSS.n200 VSS.n36 4.5005
R8253 VSS.n187 VSS.n36 4.5005
R8254 VSS.n201 VSS.n36 4.5005
R8255 VSS.n186 VSS.n36 4.5005
R8256 VSS.n202 VSS.n36 4.5005
R8257 VSS.n185 VSS.n36 4.5005
R8258 VSS.n203 VSS.n36 4.5005
R8259 VSS.n184 VSS.n36 4.5005
R8260 VSS.n204 VSS.n36 4.5005
R8261 VSS.n183 VSS.n36 4.5005
R8262 VSS.n205 VSS.n36 4.5005
R8263 VSS.n182 VSS.n36 4.5005
R8264 VSS.n206 VSS.n36 4.5005
R8265 VSS.n181 VSS.n36 4.5005
R8266 VSS.n207 VSS.n36 4.5005
R8267 VSS.n180 VSS.n36 4.5005
R8268 VSS.n208 VSS.n36 4.5005
R8269 VSS.n179 VSS.n36 4.5005
R8270 VSS.n209 VSS.n36 4.5005
R8271 VSS.n178 VSS.n36 4.5005
R8272 VSS.n210 VSS.n36 4.5005
R8273 VSS.n177 VSS.n36 4.5005
R8274 VSS.n211 VSS.n36 4.5005
R8275 VSS.n176 VSS.n36 4.5005
R8276 VSS.n212 VSS.n36 4.5005
R8277 VSS.n175 VSS.n36 4.5005
R8278 VSS.n213 VSS.n36 4.5005
R8279 VSS.n174 VSS.n36 4.5005
R8280 VSS.n214 VSS.n36 4.5005
R8281 VSS.n173 VSS.n36 4.5005
R8282 VSS.n215 VSS.n36 4.5005
R8283 VSS.n172 VSS.n36 4.5005
R8284 VSS.n216 VSS.n36 4.5005
R8285 VSS.n171 VSS.n36 4.5005
R8286 VSS.n217 VSS.n36 4.5005
R8287 VSS.n170 VSS.n36 4.5005
R8288 VSS.n218 VSS.n36 4.5005
R8289 VSS.n169 VSS.n36 4.5005
R8290 VSS.n219 VSS.n36 4.5005
R8291 VSS.n168 VSS.n36 4.5005
R8292 VSS.n220 VSS.n36 4.5005
R8293 VSS.n167 VSS.n36 4.5005
R8294 VSS.n221 VSS.n36 4.5005
R8295 VSS.n166 VSS.n36 4.5005
R8296 VSS.n222 VSS.n36 4.5005
R8297 VSS.n165 VSS.n36 4.5005
R8298 VSS.n223 VSS.n36 4.5005
R8299 VSS.n164 VSS.n36 4.5005
R8300 VSS.n224 VSS.n36 4.5005
R8301 VSS.n163 VSS.n36 4.5005
R8302 VSS.n225 VSS.n36 4.5005
R8303 VSS.n162 VSS.n36 4.5005
R8304 VSS.n226 VSS.n36 4.5005
R8305 VSS.n161 VSS.n36 4.5005
R8306 VSS.n227 VSS.n36 4.5005
R8307 VSS.n160 VSS.n36 4.5005
R8308 VSS.n228 VSS.n36 4.5005
R8309 VSS.n159 VSS.n36 4.5005
R8310 VSS.n229 VSS.n36 4.5005
R8311 VSS.n158 VSS.n36 4.5005
R8312 VSS.n230 VSS.n36 4.5005
R8313 VSS.n157 VSS.n36 4.5005
R8314 VSS.n231 VSS.n36 4.5005
R8315 VSS.n156 VSS.n36 4.5005
R8316 VSS.n232 VSS.n36 4.5005
R8317 VSS.n155 VSS.n36 4.5005
R8318 VSS.n233 VSS.n36 4.5005
R8319 VSS.n154 VSS.n36 4.5005
R8320 VSS.n234 VSS.n36 4.5005
R8321 VSS.n153 VSS.n36 4.5005
R8322 VSS.n235 VSS.n36 4.5005
R8323 VSS.n4506 VSS.n36 4.5005
R8324 VSS.n236 VSS.n36 4.5005
R8325 VSS.n152 VSS.n36 4.5005
R8326 VSS.n237 VSS.n36 4.5005
R8327 VSS.n151 VSS.n36 4.5005
R8328 VSS.n238 VSS.n36 4.5005
R8329 VSS.n150 VSS.n36 4.5005
R8330 VSS.n239 VSS.n36 4.5005
R8331 VSS.n149 VSS.n36 4.5005
R8332 VSS.n240 VSS.n36 4.5005
R8333 VSS.n148 VSS.n36 4.5005
R8334 VSS.n241 VSS.n36 4.5005
R8335 VSS.n147 VSS.n36 4.5005
R8336 VSS.n242 VSS.n36 4.5005
R8337 VSS.n146 VSS.n36 4.5005
R8338 VSS.n243 VSS.n36 4.5005
R8339 VSS.n145 VSS.n36 4.5005
R8340 VSS.n244 VSS.n36 4.5005
R8341 VSS.n144 VSS.n36 4.5005
R8342 VSS.n245 VSS.n36 4.5005
R8343 VSS.n143 VSS.n36 4.5005
R8344 VSS.n246 VSS.n36 4.5005
R8345 VSS.n142 VSS.n36 4.5005
R8346 VSS.n247 VSS.n36 4.5005
R8347 VSS.n141 VSS.n36 4.5005
R8348 VSS.n248 VSS.n36 4.5005
R8349 VSS.n140 VSS.n36 4.5005
R8350 VSS.n249 VSS.n36 4.5005
R8351 VSS.n139 VSS.n36 4.5005
R8352 VSS.n250 VSS.n36 4.5005
R8353 VSS.n138 VSS.n36 4.5005
R8354 VSS.n251 VSS.n36 4.5005
R8355 VSS.n137 VSS.n36 4.5005
R8356 VSS.n252 VSS.n36 4.5005
R8357 VSS.n136 VSS.n36 4.5005
R8358 VSS.n253 VSS.n36 4.5005
R8359 VSS.n135 VSS.n36 4.5005
R8360 VSS.n254 VSS.n36 4.5005
R8361 VSS.n134 VSS.n36 4.5005
R8362 VSS.n255 VSS.n36 4.5005
R8363 VSS.n133 VSS.n36 4.5005
R8364 VSS.n256 VSS.n36 4.5005
R8365 VSS.n132 VSS.n36 4.5005
R8366 VSS.n4502 VSS.n36 4.5005
R8367 VSS.n4504 VSS.n36 4.5005
R8368 VSS.n193 VSS.n101 4.5005
R8369 VSS.n195 VSS.n101 4.5005
R8370 VSS.n192 VSS.n101 4.5005
R8371 VSS.n196 VSS.n101 4.5005
R8372 VSS.n191 VSS.n101 4.5005
R8373 VSS.n197 VSS.n101 4.5005
R8374 VSS.n190 VSS.n101 4.5005
R8375 VSS.n198 VSS.n101 4.5005
R8376 VSS.n189 VSS.n101 4.5005
R8377 VSS.n199 VSS.n101 4.5005
R8378 VSS.n188 VSS.n101 4.5005
R8379 VSS.n200 VSS.n101 4.5005
R8380 VSS.n187 VSS.n101 4.5005
R8381 VSS.n201 VSS.n101 4.5005
R8382 VSS.n186 VSS.n101 4.5005
R8383 VSS.n202 VSS.n101 4.5005
R8384 VSS.n185 VSS.n101 4.5005
R8385 VSS.n203 VSS.n101 4.5005
R8386 VSS.n184 VSS.n101 4.5005
R8387 VSS.n204 VSS.n101 4.5005
R8388 VSS.n183 VSS.n101 4.5005
R8389 VSS.n205 VSS.n101 4.5005
R8390 VSS.n182 VSS.n101 4.5005
R8391 VSS.n206 VSS.n101 4.5005
R8392 VSS.n181 VSS.n101 4.5005
R8393 VSS.n207 VSS.n101 4.5005
R8394 VSS.n180 VSS.n101 4.5005
R8395 VSS.n208 VSS.n101 4.5005
R8396 VSS.n179 VSS.n101 4.5005
R8397 VSS.n209 VSS.n101 4.5005
R8398 VSS.n178 VSS.n101 4.5005
R8399 VSS.n210 VSS.n101 4.5005
R8400 VSS.n177 VSS.n101 4.5005
R8401 VSS.n211 VSS.n101 4.5005
R8402 VSS.n176 VSS.n101 4.5005
R8403 VSS.n212 VSS.n101 4.5005
R8404 VSS.n175 VSS.n101 4.5005
R8405 VSS.n213 VSS.n101 4.5005
R8406 VSS.n174 VSS.n101 4.5005
R8407 VSS.n214 VSS.n101 4.5005
R8408 VSS.n173 VSS.n101 4.5005
R8409 VSS.n215 VSS.n101 4.5005
R8410 VSS.n172 VSS.n101 4.5005
R8411 VSS.n216 VSS.n101 4.5005
R8412 VSS.n171 VSS.n101 4.5005
R8413 VSS.n217 VSS.n101 4.5005
R8414 VSS.n170 VSS.n101 4.5005
R8415 VSS.n218 VSS.n101 4.5005
R8416 VSS.n169 VSS.n101 4.5005
R8417 VSS.n219 VSS.n101 4.5005
R8418 VSS.n168 VSS.n101 4.5005
R8419 VSS.n220 VSS.n101 4.5005
R8420 VSS.n167 VSS.n101 4.5005
R8421 VSS.n221 VSS.n101 4.5005
R8422 VSS.n166 VSS.n101 4.5005
R8423 VSS.n222 VSS.n101 4.5005
R8424 VSS.n165 VSS.n101 4.5005
R8425 VSS.n223 VSS.n101 4.5005
R8426 VSS.n164 VSS.n101 4.5005
R8427 VSS.n224 VSS.n101 4.5005
R8428 VSS.n163 VSS.n101 4.5005
R8429 VSS.n225 VSS.n101 4.5005
R8430 VSS.n162 VSS.n101 4.5005
R8431 VSS.n226 VSS.n101 4.5005
R8432 VSS.n161 VSS.n101 4.5005
R8433 VSS.n227 VSS.n101 4.5005
R8434 VSS.n160 VSS.n101 4.5005
R8435 VSS.n228 VSS.n101 4.5005
R8436 VSS.n159 VSS.n101 4.5005
R8437 VSS.n229 VSS.n101 4.5005
R8438 VSS.n158 VSS.n101 4.5005
R8439 VSS.n230 VSS.n101 4.5005
R8440 VSS.n157 VSS.n101 4.5005
R8441 VSS.n231 VSS.n101 4.5005
R8442 VSS.n156 VSS.n101 4.5005
R8443 VSS.n232 VSS.n101 4.5005
R8444 VSS.n155 VSS.n101 4.5005
R8445 VSS.n233 VSS.n101 4.5005
R8446 VSS.n154 VSS.n101 4.5005
R8447 VSS.n234 VSS.n101 4.5005
R8448 VSS.n153 VSS.n101 4.5005
R8449 VSS.n235 VSS.n101 4.5005
R8450 VSS.n4506 VSS.n101 4.5005
R8451 VSS.n236 VSS.n101 4.5005
R8452 VSS.n152 VSS.n101 4.5005
R8453 VSS.n237 VSS.n101 4.5005
R8454 VSS.n151 VSS.n101 4.5005
R8455 VSS.n238 VSS.n101 4.5005
R8456 VSS.n150 VSS.n101 4.5005
R8457 VSS.n239 VSS.n101 4.5005
R8458 VSS.n149 VSS.n101 4.5005
R8459 VSS.n240 VSS.n101 4.5005
R8460 VSS.n148 VSS.n101 4.5005
R8461 VSS.n241 VSS.n101 4.5005
R8462 VSS.n147 VSS.n101 4.5005
R8463 VSS.n242 VSS.n101 4.5005
R8464 VSS.n146 VSS.n101 4.5005
R8465 VSS.n243 VSS.n101 4.5005
R8466 VSS.n145 VSS.n101 4.5005
R8467 VSS.n244 VSS.n101 4.5005
R8468 VSS.n144 VSS.n101 4.5005
R8469 VSS.n245 VSS.n101 4.5005
R8470 VSS.n143 VSS.n101 4.5005
R8471 VSS.n246 VSS.n101 4.5005
R8472 VSS.n142 VSS.n101 4.5005
R8473 VSS.n247 VSS.n101 4.5005
R8474 VSS.n141 VSS.n101 4.5005
R8475 VSS.n248 VSS.n101 4.5005
R8476 VSS.n140 VSS.n101 4.5005
R8477 VSS.n249 VSS.n101 4.5005
R8478 VSS.n139 VSS.n101 4.5005
R8479 VSS.n250 VSS.n101 4.5005
R8480 VSS.n138 VSS.n101 4.5005
R8481 VSS.n251 VSS.n101 4.5005
R8482 VSS.n137 VSS.n101 4.5005
R8483 VSS.n252 VSS.n101 4.5005
R8484 VSS.n136 VSS.n101 4.5005
R8485 VSS.n253 VSS.n101 4.5005
R8486 VSS.n135 VSS.n101 4.5005
R8487 VSS.n254 VSS.n101 4.5005
R8488 VSS.n134 VSS.n101 4.5005
R8489 VSS.n255 VSS.n101 4.5005
R8490 VSS.n133 VSS.n101 4.5005
R8491 VSS.n256 VSS.n101 4.5005
R8492 VSS.n132 VSS.n101 4.5005
R8493 VSS.n4502 VSS.n101 4.5005
R8494 VSS.n4504 VSS.n101 4.5005
R8495 VSS.n193 VSS.n35 4.5005
R8496 VSS.n195 VSS.n35 4.5005
R8497 VSS.n192 VSS.n35 4.5005
R8498 VSS.n196 VSS.n35 4.5005
R8499 VSS.n191 VSS.n35 4.5005
R8500 VSS.n197 VSS.n35 4.5005
R8501 VSS.n190 VSS.n35 4.5005
R8502 VSS.n198 VSS.n35 4.5005
R8503 VSS.n189 VSS.n35 4.5005
R8504 VSS.n199 VSS.n35 4.5005
R8505 VSS.n188 VSS.n35 4.5005
R8506 VSS.n200 VSS.n35 4.5005
R8507 VSS.n187 VSS.n35 4.5005
R8508 VSS.n201 VSS.n35 4.5005
R8509 VSS.n186 VSS.n35 4.5005
R8510 VSS.n202 VSS.n35 4.5005
R8511 VSS.n185 VSS.n35 4.5005
R8512 VSS.n203 VSS.n35 4.5005
R8513 VSS.n184 VSS.n35 4.5005
R8514 VSS.n204 VSS.n35 4.5005
R8515 VSS.n183 VSS.n35 4.5005
R8516 VSS.n205 VSS.n35 4.5005
R8517 VSS.n182 VSS.n35 4.5005
R8518 VSS.n206 VSS.n35 4.5005
R8519 VSS.n181 VSS.n35 4.5005
R8520 VSS.n207 VSS.n35 4.5005
R8521 VSS.n180 VSS.n35 4.5005
R8522 VSS.n208 VSS.n35 4.5005
R8523 VSS.n179 VSS.n35 4.5005
R8524 VSS.n209 VSS.n35 4.5005
R8525 VSS.n178 VSS.n35 4.5005
R8526 VSS.n210 VSS.n35 4.5005
R8527 VSS.n177 VSS.n35 4.5005
R8528 VSS.n211 VSS.n35 4.5005
R8529 VSS.n176 VSS.n35 4.5005
R8530 VSS.n212 VSS.n35 4.5005
R8531 VSS.n175 VSS.n35 4.5005
R8532 VSS.n213 VSS.n35 4.5005
R8533 VSS.n174 VSS.n35 4.5005
R8534 VSS.n214 VSS.n35 4.5005
R8535 VSS.n173 VSS.n35 4.5005
R8536 VSS.n215 VSS.n35 4.5005
R8537 VSS.n172 VSS.n35 4.5005
R8538 VSS.n216 VSS.n35 4.5005
R8539 VSS.n171 VSS.n35 4.5005
R8540 VSS.n217 VSS.n35 4.5005
R8541 VSS.n170 VSS.n35 4.5005
R8542 VSS.n218 VSS.n35 4.5005
R8543 VSS.n169 VSS.n35 4.5005
R8544 VSS.n219 VSS.n35 4.5005
R8545 VSS.n168 VSS.n35 4.5005
R8546 VSS.n220 VSS.n35 4.5005
R8547 VSS.n167 VSS.n35 4.5005
R8548 VSS.n221 VSS.n35 4.5005
R8549 VSS.n166 VSS.n35 4.5005
R8550 VSS.n222 VSS.n35 4.5005
R8551 VSS.n165 VSS.n35 4.5005
R8552 VSS.n223 VSS.n35 4.5005
R8553 VSS.n164 VSS.n35 4.5005
R8554 VSS.n224 VSS.n35 4.5005
R8555 VSS.n163 VSS.n35 4.5005
R8556 VSS.n225 VSS.n35 4.5005
R8557 VSS.n162 VSS.n35 4.5005
R8558 VSS.n226 VSS.n35 4.5005
R8559 VSS.n161 VSS.n35 4.5005
R8560 VSS.n227 VSS.n35 4.5005
R8561 VSS.n160 VSS.n35 4.5005
R8562 VSS.n228 VSS.n35 4.5005
R8563 VSS.n159 VSS.n35 4.5005
R8564 VSS.n229 VSS.n35 4.5005
R8565 VSS.n158 VSS.n35 4.5005
R8566 VSS.n230 VSS.n35 4.5005
R8567 VSS.n157 VSS.n35 4.5005
R8568 VSS.n231 VSS.n35 4.5005
R8569 VSS.n156 VSS.n35 4.5005
R8570 VSS.n232 VSS.n35 4.5005
R8571 VSS.n155 VSS.n35 4.5005
R8572 VSS.n233 VSS.n35 4.5005
R8573 VSS.n154 VSS.n35 4.5005
R8574 VSS.n234 VSS.n35 4.5005
R8575 VSS.n153 VSS.n35 4.5005
R8576 VSS.n235 VSS.n35 4.5005
R8577 VSS.n4506 VSS.n35 4.5005
R8578 VSS.n236 VSS.n35 4.5005
R8579 VSS.n152 VSS.n35 4.5005
R8580 VSS.n237 VSS.n35 4.5005
R8581 VSS.n151 VSS.n35 4.5005
R8582 VSS.n238 VSS.n35 4.5005
R8583 VSS.n150 VSS.n35 4.5005
R8584 VSS.n239 VSS.n35 4.5005
R8585 VSS.n149 VSS.n35 4.5005
R8586 VSS.n240 VSS.n35 4.5005
R8587 VSS.n148 VSS.n35 4.5005
R8588 VSS.n241 VSS.n35 4.5005
R8589 VSS.n147 VSS.n35 4.5005
R8590 VSS.n242 VSS.n35 4.5005
R8591 VSS.n146 VSS.n35 4.5005
R8592 VSS.n243 VSS.n35 4.5005
R8593 VSS.n145 VSS.n35 4.5005
R8594 VSS.n244 VSS.n35 4.5005
R8595 VSS.n144 VSS.n35 4.5005
R8596 VSS.n245 VSS.n35 4.5005
R8597 VSS.n143 VSS.n35 4.5005
R8598 VSS.n246 VSS.n35 4.5005
R8599 VSS.n142 VSS.n35 4.5005
R8600 VSS.n247 VSS.n35 4.5005
R8601 VSS.n141 VSS.n35 4.5005
R8602 VSS.n248 VSS.n35 4.5005
R8603 VSS.n140 VSS.n35 4.5005
R8604 VSS.n249 VSS.n35 4.5005
R8605 VSS.n139 VSS.n35 4.5005
R8606 VSS.n250 VSS.n35 4.5005
R8607 VSS.n138 VSS.n35 4.5005
R8608 VSS.n251 VSS.n35 4.5005
R8609 VSS.n137 VSS.n35 4.5005
R8610 VSS.n252 VSS.n35 4.5005
R8611 VSS.n136 VSS.n35 4.5005
R8612 VSS.n253 VSS.n35 4.5005
R8613 VSS.n135 VSS.n35 4.5005
R8614 VSS.n254 VSS.n35 4.5005
R8615 VSS.n134 VSS.n35 4.5005
R8616 VSS.n255 VSS.n35 4.5005
R8617 VSS.n133 VSS.n35 4.5005
R8618 VSS.n256 VSS.n35 4.5005
R8619 VSS.n132 VSS.n35 4.5005
R8620 VSS.n4502 VSS.n35 4.5005
R8621 VSS.n4504 VSS.n35 4.5005
R8622 VSS.n193 VSS.n102 4.5005
R8623 VSS.n195 VSS.n102 4.5005
R8624 VSS.n192 VSS.n102 4.5005
R8625 VSS.n196 VSS.n102 4.5005
R8626 VSS.n191 VSS.n102 4.5005
R8627 VSS.n197 VSS.n102 4.5005
R8628 VSS.n190 VSS.n102 4.5005
R8629 VSS.n198 VSS.n102 4.5005
R8630 VSS.n189 VSS.n102 4.5005
R8631 VSS.n199 VSS.n102 4.5005
R8632 VSS.n188 VSS.n102 4.5005
R8633 VSS.n200 VSS.n102 4.5005
R8634 VSS.n187 VSS.n102 4.5005
R8635 VSS.n201 VSS.n102 4.5005
R8636 VSS.n186 VSS.n102 4.5005
R8637 VSS.n202 VSS.n102 4.5005
R8638 VSS.n185 VSS.n102 4.5005
R8639 VSS.n203 VSS.n102 4.5005
R8640 VSS.n184 VSS.n102 4.5005
R8641 VSS.n204 VSS.n102 4.5005
R8642 VSS.n183 VSS.n102 4.5005
R8643 VSS.n205 VSS.n102 4.5005
R8644 VSS.n182 VSS.n102 4.5005
R8645 VSS.n206 VSS.n102 4.5005
R8646 VSS.n181 VSS.n102 4.5005
R8647 VSS.n207 VSS.n102 4.5005
R8648 VSS.n180 VSS.n102 4.5005
R8649 VSS.n208 VSS.n102 4.5005
R8650 VSS.n179 VSS.n102 4.5005
R8651 VSS.n209 VSS.n102 4.5005
R8652 VSS.n178 VSS.n102 4.5005
R8653 VSS.n210 VSS.n102 4.5005
R8654 VSS.n177 VSS.n102 4.5005
R8655 VSS.n211 VSS.n102 4.5005
R8656 VSS.n176 VSS.n102 4.5005
R8657 VSS.n212 VSS.n102 4.5005
R8658 VSS.n175 VSS.n102 4.5005
R8659 VSS.n213 VSS.n102 4.5005
R8660 VSS.n174 VSS.n102 4.5005
R8661 VSS.n214 VSS.n102 4.5005
R8662 VSS.n173 VSS.n102 4.5005
R8663 VSS.n215 VSS.n102 4.5005
R8664 VSS.n172 VSS.n102 4.5005
R8665 VSS.n216 VSS.n102 4.5005
R8666 VSS.n171 VSS.n102 4.5005
R8667 VSS.n217 VSS.n102 4.5005
R8668 VSS.n170 VSS.n102 4.5005
R8669 VSS.n218 VSS.n102 4.5005
R8670 VSS.n169 VSS.n102 4.5005
R8671 VSS.n219 VSS.n102 4.5005
R8672 VSS.n168 VSS.n102 4.5005
R8673 VSS.n220 VSS.n102 4.5005
R8674 VSS.n167 VSS.n102 4.5005
R8675 VSS.n221 VSS.n102 4.5005
R8676 VSS.n166 VSS.n102 4.5005
R8677 VSS.n222 VSS.n102 4.5005
R8678 VSS.n165 VSS.n102 4.5005
R8679 VSS.n223 VSS.n102 4.5005
R8680 VSS.n164 VSS.n102 4.5005
R8681 VSS.n224 VSS.n102 4.5005
R8682 VSS.n163 VSS.n102 4.5005
R8683 VSS.n225 VSS.n102 4.5005
R8684 VSS.n162 VSS.n102 4.5005
R8685 VSS.n226 VSS.n102 4.5005
R8686 VSS.n161 VSS.n102 4.5005
R8687 VSS.n227 VSS.n102 4.5005
R8688 VSS.n160 VSS.n102 4.5005
R8689 VSS.n228 VSS.n102 4.5005
R8690 VSS.n159 VSS.n102 4.5005
R8691 VSS.n229 VSS.n102 4.5005
R8692 VSS.n158 VSS.n102 4.5005
R8693 VSS.n230 VSS.n102 4.5005
R8694 VSS.n157 VSS.n102 4.5005
R8695 VSS.n231 VSS.n102 4.5005
R8696 VSS.n156 VSS.n102 4.5005
R8697 VSS.n232 VSS.n102 4.5005
R8698 VSS.n155 VSS.n102 4.5005
R8699 VSS.n233 VSS.n102 4.5005
R8700 VSS.n154 VSS.n102 4.5005
R8701 VSS.n234 VSS.n102 4.5005
R8702 VSS.n153 VSS.n102 4.5005
R8703 VSS.n235 VSS.n102 4.5005
R8704 VSS.n4506 VSS.n102 4.5005
R8705 VSS.n236 VSS.n102 4.5005
R8706 VSS.n152 VSS.n102 4.5005
R8707 VSS.n237 VSS.n102 4.5005
R8708 VSS.n151 VSS.n102 4.5005
R8709 VSS.n238 VSS.n102 4.5005
R8710 VSS.n150 VSS.n102 4.5005
R8711 VSS.n239 VSS.n102 4.5005
R8712 VSS.n149 VSS.n102 4.5005
R8713 VSS.n240 VSS.n102 4.5005
R8714 VSS.n148 VSS.n102 4.5005
R8715 VSS.n241 VSS.n102 4.5005
R8716 VSS.n147 VSS.n102 4.5005
R8717 VSS.n242 VSS.n102 4.5005
R8718 VSS.n146 VSS.n102 4.5005
R8719 VSS.n243 VSS.n102 4.5005
R8720 VSS.n145 VSS.n102 4.5005
R8721 VSS.n244 VSS.n102 4.5005
R8722 VSS.n144 VSS.n102 4.5005
R8723 VSS.n245 VSS.n102 4.5005
R8724 VSS.n143 VSS.n102 4.5005
R8725 VSS.n246 VSS.n102 4.5005
R8726 VSS.n142 VSS.n102 4.5005
R8727 VSS.n247 VSS.n102 4.5005
R8728 VSS.n141 VSS.n102 4.5005
R8729 VSS.n248 VSS.n102 4.5005
R8730 VSS.n140 VSS.n102 4.5005
R8731 VSS.n249 VSS.n102 4.5005
R8732 VSS.n139 VSS.n102 4.5005
R8733 VSS.n250 VSS.n102 4.5005
R8734 VSS.n138 VSS.n102 4.5005
R8735 VSS.n251 VSS.n102 4.5005
R8736 VSS.n137 VSS.n102 4.5005
R8737 VSS.n252 VSS.n102 4.5005
R8738 VSS.n136 VSS.n102 4.5005
R8739 VSS.n253 VSS.n102 4.5005
R8740 VSS.n135 VSS.n102 4.5005
R8741 VSS.n254 VSS.n102 4.5005
R8742 VSS.n134 VSS.n102 4.5005
R8743 VSS.n255 VSS.n102 4.5005
R8744 VSS.n133 VSS.n102 4.5005
R8745 VSS.n256 VSS.n102 4.5005
R8746 VSS.n132 VSS.n102 4.5005
R8747 VSS.n4502 VSS.n102 4.5005
R8748 VSS.n4504 VSS.n102 4.5005
R8749 VSS.n193 VSS.n34 4.5005
R8750 VSS.n195 VSS.n34 4.5005
R8751 VSS.n192 VSS.n34 4.5005
R8752 VSS.n196 VSS.n34 4.5005
R8753 VSS.n191 VSS.n34 4.5005
R8754 VSS.n197 VSS.n34 4.5005
R8755 VSS.n190 VSS.n34 4.5005
R8756 VSS.n198 VSS.n34 4.5005
R8757 VSS.n189 VSS.n34 4.5005
R8758 VSS.n199 VSS.n34 4.5005
R8759 VSS.n188 VSS.n34 4.5005
R8760 VSS.n200 VSS.n34 4.5005
R8761 VSS.n187 VSS.n34 4.5005
R8762 VSS.n201 VSS.n34 4.5005
R8763 VSS.n186 VSS.n34 4.5005
R8764 VSS.n202 VSS.n34 4.5005
R8765 VSS.n185 VSS.n34 4.5005
R8766 VSS.n203 VSS.n34 4.5005
R8767 VSS.n184 VSS.n34 4.5005
R8768 VSS.n204 VSS.n34 4.5005
R8769 VSS.n183 VSS.n34 4.5005
R8770 VSS.n205 VSS.n34 4.5005
R8771 VSS.n182 VSS.n34 4.5005
R8772 VSS.n206 VSS.n34 4.5005
R8773 VSS.n181 VSS.n34 4.5005
R8774 VSS.n207 VSS.n34 4.5005
R8775 VSS.n180 VSS.n34 4.5005
R8776 VSS.n208 VSS.n34 4.5005
R8777 VSS.n179 VSS.n34 4.5005
R8778 VSS.n209 VSS.n34 4.5005
R8779 VSS.n178 VSS.n34 4.5005
R8780 VSS.n210 VSS.n34 4.5005
R8781 VSS.n177 VSS.n34 4.5005
R8782 VSS.n211 VSS.n34 4.5005
R8783 VSS.n176 VSS.n34 4.5005
R8784 VSS.n212 VSS.n34 4.5005
R8785 VSS.n175 VSS.n34 4.5005
R8786 VSS.n213 VSS.n34 4.5005
R8787 VSS.n174 VSS.n34 4.5005
R8788 VSS.n214 VSS.n34 4.5005
R8789 VSS.n173 VSS.n34 4.5005
R8790 VSS.n215 VSS.n34 4.5005
R8791 VSS.n172 VSS.n34 4.5005
R8792 VSS.n216 VSS.n34 4.5005
R8793 VSS.n171 VSS.n34 4.5005
R8794 VSS.n217 VSS.n34 4.5005
R8795 VSS.n170 VSS.n34 4.5005
R8796 VSS.n218 VSS.n34 4.5005
R8797 VSS.n169 VSS.n34 4.5005
R8798 VSS.n219 VSS.n34 4.5005
R8799 VSS.n168 VSS.n34 4.5005
R8800 VSS.n220 VSS.n34 4.5005
R8801 VSS.n167 VSS.n34 4.5005
R8802 VSS.n221 VSS.n34 4.5005
R8803 VSS.n166 VSS.n34 4.5005
R8804 VSS.n222 VSS.n34 4.5005
R8805 VSS.n165 VSS.n34 4.5005
R8806 VSS.n223 VSS.n34 4.5005
R8807 VSS.n164 VSS.n34 4.5005
R8808 VSS.n224 VSS.n34 4.5005
R8809 VSS.n163 VSS.n34 4.5005
R8810 VSS.n225 VSS.n34 4.5005
R8811 VSS.n162 VSS.n34 4.5005
R8812 VSS.n226 VSS.n34 4.5005
R8813 VSS.n161 VSS.n34 4.5005
R8814 VSS.n227 VSS.n34 4.5005
R8815 VSS.n160 VSS.n34 4.5005
R8816 VSS.n228 VSS.n34 4.5005
R8817 VSS.n159 VSS.n34 4.5005
R8818 VSS.n229 VSS.n34 4.5005
R8819 VSS.n158 VSS.n34 4.5005
R8820 VSS.n230 VSS.n34 4.5005
R8821 VSS.n157 VSS.n34 4.5005
R8822 VSS.n231 VSS.n34 4.5005
R8823 VSS.n156 VSS.n34 4.5005
R8824 VSS.n232 VSS.n34 4.5005
R8825 VSS.n155 VSS.n34 4.5005
R8826 VSS.n233 VSS.n34 4.5005
R8827 VSS.n154 VSS.n34 4.5005
R8828 VSS.n234 VSS.n34 4.5005
R8829 VSS.n153 VSS.n34 4.5005
R8830 VSS.n235 VSS.n34 4.5005
R8831 VSS.n4506 VSS.n34 4.5005
R8832 VSS.n236 VSS.n34 4.5005
R8833 VSS.n152 VSS.n34 4.5005
R8834 VSS.n237 VSS.n34 4.5005
R8835 VSS.n151 VSS.n34 4.5005
R8836 VSS.n238 VSS.n34 4.5005
R8837 VSS.n150 VSS.n34 4.5005
R8838 VSS.n239 VSS.n34 4.5005
R8839 VSS.n149 VSS.n34 4.5005
R8840 VSS.n240 VSS.n34 4.5005
R8841 VSS.n148 VSS.n34 4.5005
R8842 VSS.n241 VSS.n34 4.5005
R8843 VSS.n147 VSS.n34 4.5005
R8844 VSS.n242 VSS.n34 4.5005
R8845 VSS.n146 VSS.n34 4.5005
R8846 VSS.n243 VSS.n34 4.5005
R8847 VSS.n145 VSS.n34 4.5005
R8848 VSS.n244 VSS.n34 4.5005
R8849 VSS.n144 VSS.n34 4.5005
R8850 VSS.n245 VSS.n34 4.5005
R8851 VSS.n143 VSS.n34 4.5005
R8852 VSS.n246 VSS.n34 4.5005
R8853 VSS.n142 VSS.n34 4.5005
R8854 VSS.n247 VSS.n34 4.5005
R8855 VSS.n141 VSS.n34 4.5005
R8856 VSS.n248 VSS.n34 4.5005
R8857 VSS.n140 VSS.n34 4.5005
R8858 VSS.n249 VSS.n34 4.5005
R8859 VSS.n139 VSS.n34 4.5005
R8860 VSS.n250 VSS.n34 4.5005
R8861 VSS.n138 VSS.n34 4.5005
R8862 VSS.n251 VSS.n34 4.5005
R8863 VSS.n137 VSS.n34 4.5005
R8864 VSS.n252 VSS.n34 4.5005
R8865 VSS.n136 VSS.n34 4.5005
R8866 VSS.n253 VSS.n34 4.5005
R8867 VSS.n135 VSS.n34 4.5005
R8868 VSS.n254 VSS.n34 4.5005
R8869 VSS.n134 VSS.n34 4.5005
R8870 VSS.n255 VSS.n34 4.5005
R8871 VSS.n133 VSS.n34 4.5005
R8872 VSS.n256 VSS.n34 4.5005
R8873 VSS.n132 VSS.n34 4.5005
R8874 VSS.n4502 VSS.n34 4.5005
R8875 VSS.n4504 VSS.n34 4.5005
R8876 VSS.n193 VSS.n103 4.5005
R8877 VSS.n195 VSS.n103 4.5005
R8878 VSS.n192 VSS.n103 4.5005
R8879 VSS.n196 VSS.n103 4.5005
R8880 VSS.n191 VSS.n103 4.5005
R8881 VSS.n197 VSS.n103 4.5005
R8882 VSS.n190 VSS.n103 4.5005
R8883 VSS.n198 VSS.n103 4.5005
R8884 VSS.n189 VSS.n103 4.5005
R8885 VSS.n199 VSS.n103 4.5005
R8886 VSS.n188 VSS.n103 4.5005
R8887 VSS.n200 VSS.n103 4.5005
R8888 VSS.n187 VSS.n103 4.5005
R8889 VSS.n201 VSS.n103 4.5005
R8890 VSS.n186 VSS.n103 4.5005
R8891 VSS.n202 VSS.n103 4.5005
R8892 VSS.n185 VSS.n103 4.5005
R8893 VSS.n203 VSS.n103 4.5005
R8894 VSS.n184 VSS.n103 4.5005
R8895 VSS.n204 VSS.n103 4.5005
R8896 VSS.n183 VSS.n103 4.5005
R8897 VSS.n205 VSS.n103 4.5005
R8898 VSS.n182 VSS.n103 4.5005
R8899 VSS.n206 VSS.n103 4.5005
R8900 VSS.n181 VSS.n103 4.5005
R8901 VSS.n207 VSS.n103 4.5005
R8902 VSS.n180 VSS.n103 4.5005
R8903 VSS.n208 VSS.n103 4.5005
R8904 VSS.n179 VSS.n103 4.5005
R8905 VSS.n209 VSS.n103 4.5005
R8906 VSS.n178 VSS.n103 4.5005
R8907 VSS.n210 VSS.n103 4.5005
R8908 VSS.n177 VSS.n103 4.5005
R8909 VSS.n211 VSS.n103 4.5005
R8910 VSS.n176 VSS.n103 4.5005
R8911 VSS.n212 VSS.n103 4.5005
R8912 VSS.n175 VSS.n103 4.5005
R8913 VSS.n213 VSS.n103 4.5005
R8914 VSS.n174 VSS.n103 4.5005
R8915 VSS.n214 VSS.n103 4.5005
R8916 VSS.n173 VSS.n103 4.5005
R8917 VSS.n215 VSS.n103 4.5005
R8918 VSS.n172 VSS.n103 4.5005
R8919 VSS.n216 VSS.n103 4.5005
R8920 VSS.n171 VSS.n103 4.5005
R8921 VSS.n217 VSS.n103 4.5005
R8922 VSS.n170 VSS.n103 4.5005
R8923 VSS.n218 VSS.n103 4.5005
R8924 VSS.n169 VSS.n103 4.5005
R8925 VSS.n219 VSS.n103 4.5005
R8926 VSS.n168 VSS.n103 4.5005
R8927 VSS.n220 VSS.n103 4.5005
R8928 VSS.n167 VSS.n103 4.5005
R8929 VSS.n221 VSS.n103 4.5005
R8930 VSS.n166 VSS.n103 4.5005
R8931 VSS.n222 VSS.n103 4.5005
R8932 VSS.n165 VSS.n103 4.5005
R8933 VSS.n223 VSS.n103 4.5005
R8934 VSS.n164 VSS.n103 4.5005
R8935 VSS.n224 VSS.n103 4.5005
R8936 VSS.n163 VSS.n103 4.5005
R8937 VSS.n225 VSS.n103 4.5005
R8938 VSS.n162 VSS.n103 4.5005
R8939 VSS.n226 VSS.n103 4.5005
R8940 VSS.n161 VSS.n103 4.5005
R8941 VSS.n227 VSS.n103 4.5005
R8942 VSS.n160 VSS.n103 4.5005
R8943 VSS.n228 VSS.n103 4.5005
R8944 VSS.n159 VSS.n103 4.5005
R8945 VSS.n229 VSS.n103 4.5005
R8946 VSS.n158 VSS.n103 4.5005
R8947 VSS.n230 VSS.n103 4.5005
R8948 VSS.n157 VSS.n103 4.5005
R8949 VSS.n231 VSS.n103 4.5005
R8950 VSS.n156 VSS.n103 4.5005
R8951 VSS.n232 VSS.n103 4.5005
R8952 VSS.n155 VSS.n103 4.5005
R8953 VSS.n233 VSS.n103 4.5005
R8954 VSS.n154 VSS.n103 4.5005
R8955 VSS.n234 VSS.n103 4.5005
R8956 VSS.n153 VSS.n103 4.5005
R8957 VSS.n235 VSS.n103 4.5005
R8958 VSS.n4506 VSS.n103 4.5005
R8959 VSS.n236 VSS.n103 4.5005
R8960 VSS.n152 VSS.n103 4.5005
R8961 VSS.n237 VSS.n103 4.5005
R8962 VSS.n151 VSS.n103 4.5005
R8963 VSS.n238 VSS.n103 4.5005
R8964 VSS.n150 VSS.n103 4.5005
R8965 VSS.n239 VSS.n103 4.5005
R8966 VSS.n149 VSS.n103 4.5005
R8967 VSS.n240 VSS.n103 4.5005
R8968 VSS.n148 VSS.n103 4.5005
R8969 VSS.n241 VSS.n103 4.5005
R8970 VSS.n147 VSS.n103 4.5005
R8971 VSS.n242 VSS.n103 4.5005
R8972 VSS.n146 VSS.n103 4.5005
R8973 VSS.n243 VSS.n103 4.5005
R8974 VSS.n145 VSS.n103 4.5005
R8975 VSS.n244 VSS.n103 4.5005
R8976 VSS.n144 VSS.n103 4.5005
R8977 VSS.n245 VSS.n103 4.5005
R8978 VSS.n143 VSS.n103 4.5005
R8979 VSS.n246 VSS.n103 4.5005
R8980 VSS.n142 VSS.n103 4.5005
R8981 VSS.n247 VSS.n103 4.5005
R8982 VSS.n141 VSS.n103 4.5005
R8983 VSS.n248 VSS.n103 4.5005
R8984 VSS.n140 VSS.n103 4.5005
R8985 VSS.n249 VSS.n103 4.5005
R8986 VSS.n139 VSS.n103 4.5005
R8987 VSS.n250 VSS.n103 4.5005
R8988 VSS.n138 VSS.n103 4.5005
R8989 VSS.n251 VSS.n103 4.5005
R8990 VSS.n137 VSS.n103 4.5005
R8991 VSS.n252 VSS.n103 4.5005
R8992 VSS.n136 VSS.n103 4.5005
R8993 VSS.n253 VSS.n103 4.5005
R8994 VSS.n135 VSS.n103 4.5005
R8995 VSS.n254 VSS.n103 4.5005
R8996 VSS.n134 VSS.n103 4.5005
R8997 VSS.n255 VSS.n103 4.5005
R8998 VSS.n133 VSS.n103 4.5005
R8999 VSS.n256 VSS.n103 4.5005
R9000 VSS.n132 VSS.n103 4.5005
R9001 VSS.n4502 VSS.n103 4.5005
R9002 VSS.n4504 VSS.n103 4.5005
R9003 VSS.n193 VSS.n33 4.5005
R9004 VSS.n195 VSS.n33 4.5005
R9005 VSS.n192 VSS.n33 4.5005
R9006 VSS.n196 VSS.n33 4.5005
R9007 VSS.n191 VSS.n33 4.5005
R9008 VSS.n197 VSS.n33 4.5005
R9009 VSS.n190 VSS.n33 4.5005
R9010 VSS.n198 VSS.n33 4.5005
R9011 VSS.n189 VSS.n33 4.5005
R9012 VSS.n199 VSS.n33 4.5005
R9013 VSS.n188 VSS.n33 4.5005
R9014 VSS.n200 VSS.n33 4.5005
R9015 VSS.n187 VSS.n33 4.5005
R9016 VSS.n201 VSS.n33 4.5005
R9017 VSS.n186 VSS.n33 4.5005
R9018 VSS.n202 VSS.n33 4.5005
R9019 VSS.n185 VSS.n33 4.5005
R9020 VSS.n203 VSS.n33 4.5005
R9021 VSS.n184 VSS.n33 4.5005
R9022 VSS.n204 VSS.n33 4.5005
R9023 VSS.n183 VSS.n33 4.5005
R9024 VSS.n205 VSS.n33 4.5005
R9025 VSS.n182 VSS.n33 4.5005
R9026 VSS.n206 VSS.n33 4.5005
R9027 VSS.n181 VSS.n33 4.5005
R9028 VSS.n207 VSS.n33 4.5005
R9029 VSS.n180 VSS.n33 4.5005
R9030 VSS.n208 VSS.n33 4.5005
R9031 VSS.n179 VSS.n33 4.5005
R9032 VSS.n209 VSS.n33 4.5005
R9033 VSS.n178 VSS.n33 4.5005
R9034 VSS.n210 VSS.n33 4.5005
R9035 VSS.n177 VSS.n33 4.5005
R9036 VSS.n211 VSS.n33 4.5005
R9037 VSS.n176 VSS.n33 4.5005
R9038 VSS.n212 VSS.n33 4.5005
R9039 VSS.n175 VSS.n33 4.5005
R9040 VSS.n213 VSS.n33 4.5005
R9041 VSS.n174 VSS.n33 4.5005
R9042 VSS.n214 VSS.n33 4.5005
R9043 VSS.n173 VSS.n33 4.5005
R9044 VSS.n215 VSS.n33 4.5005
R9045 VSS.n172 VSS.n33 4.5005
R9046 VSS.n216 VSS.n33 4.5005
R9047 VSS.n171 VSS.n33 4.5005
R9048 VSS.n217 VSS.n33 4.5005
R9049 VSS.n170 VSS.n33 4.5005
R9050 VSS.n218 VSS.n33 4.5005
R9051 VSS.n169 VSS.n33 4.5005
R9052 VSS.n219 VSS.n33 4.5005
R9053 VSS.n168 VSS.n33 4.5005
R9054 VSS.n220 VSS.n33 4.5005
R9055 VSS.n167 VSS.n33 4.5005
R9056 VSS.n221 VSS.n33 4.5005
R9057 VSS.n166 VSS.n33 4.5005
R9058 VSS.n222 VSS.n33 4.5005
R9059 VSS.n165 VSS.n33 4.5005
R9060 VSS.n223 VSS.n33 4.5005
R9061 VSS.n164 VSS.n33 4.5005
R9062 VSS.n224 VSS.n33 4.5005
R9063 VSS.n163 VSS.n33 4.5005
R9064 VSS.n225 VSS.n33 4.5005
R9065 VSS.n162 VSS.n33 4.5005
R9066 VSS.n226 VSS.n33 4.5005
R9067 VSS.n161 VSS.n33 4.5005
R9068 VSS.n227 VSS.n33 4.5005
R9069 VSS.n160 VSS.n33 4.5005
R9070 VSS.n228 VSS.n33 4.5005
R9071 VSS.n159 VSS.n33 4.5005
R9072 VSS.n229 VSS.n33 4.5005
R9073 VSS.n158 VSS.n33 4.5005
R9074 VSS.n230 VSS.n33 4.5005
R9075 VSS.n157 VSS.n33 4.5005
R9076 VSS.n231 VSS.n33 4.5005
R9077 VSS.n156 VSS.n33 4.5005
R9078 VSS.n232 VSS.n33 4.5005
R9079 VSS.n155 VSS.n33 4.5005
R9080 VSS.n233 VSS.n33 4.5005
R9081 VSS.n154 VSS.n33 4.5005
R9082 VSS.n234 VSS.n33 4.5005
R9083 VSS.n153 VSS.n33 4.5005
R9084 VSS.n235 VSS.n33 4.5005
R9085 VSS.n4506 VSS.n33 4.5005
R9086 VSS.n236 VSS.n33 4.5005
R9087 VSS.n152 VSS.n33 4.5005
R9088 VSS.n237 VSS.n33 4.5005
R9089 VSS.n151 VSS.n33 4.5005
R9090 VSS.n238 VSS.n33 4.5005
R9091 VSS.n150 VSS.n33 4.5005
R9092 VSS.n239 VSS.n33 4.5005
R9093 VSS.n149 VSS.n33 4.5005
R9094 VSS.n240 VSS.n33 4.5005
R9095 VSS.n148 VSS.n33 4.5005
R9096 VSS.n241 VSS.n33 4.5005
R9097 VSS.n147 VSS.n33 4.5005
R9098 VSS.n242 VSS.n33 4.5005
R9099 VSS.n146 VSS.n33 4.5005
R9100 VSS.n243 VSS.n33 4.5005
R9101 VSS.n145 VSS.n33 4.5005
R9102 VSS.n244 VSS.n33 4.5005
R9103 VSS.n144 VSS.n33 4.5005
R9104 VSS.n245 VSS.n33 4.5005
R9105 VSS.n143 VSS.n33 4.5005
R9106 VSS.n246 VSS.n33 4.5005
R9107 VSS.n142 VSS.n33 4.5005
R9108 VSS.n247 VSS.n33 4.5005
R9109 VSS.n141 VSS.n33 4.5005
R9110 VSS.n248 VSS.n33 4.5005
R9111 VSS.n140 VSS.n33 4.5005
R9112 VSS.n249 VSS.n33 4.5005
R9113 VSS.n139 VSS.n33 4.5005
R9114 VSS.n250 VSS.n33 4.5005
R9115 VSS.n138 VSS.n33 4.5005
R9116 VSS.n251 VSS.n33 4.5005
R9117 VSS.n137 VSS.n33 4.5005
R9118 VSS.n252 VSS.n33 4.5005
R9119 VSS.n136 VSS.n33 4.5005
R9120 VSS.n253 VSS.n33 4.5005
R9121 VSS.n135 VSS.n33 4.5005
R9122 VSS.n254 VSS.n33 4.5005
R9123 VSS.n134 VSS.n33 4.5005
R9124 VSS.n255 VSS.n33 4.5005
R9125 VSS.n133 VSS.n33 4.5005
R9126 VSS.n256 VSS.n33 4.5005
R9127 VSS.n132 VSS.n33 4.5005
R9128 VSS.n4502 VSS.n33 4.5005
R9129 VSS.n4504 VSS.n33 4.5005
R9130 VSS.n193 VSS.n104 4.5005
R9131 VSS.n195 VSS.n104 4.5005
R9132 VSS.n192 VSS.n104 4.5005
R9133 VSS.n196 VSS.n104 4.5005
R9134 VSS.n191 VSS.n104 4.5005
R9135 VSS.n197 VSS.n104 4.5005
R9136 VSS.n190 VSS.n104 4.5005
R9137 VSS.n198 VSS.n104 4.5005
R9138 VSS.n189 VSS.n104 4.5005
R9139 VSS.n199 VSS.n104 4.5005
R9140 VSS.n188 VSS.n104 4.5005
R9141 VSS.n200 VSS.n104 4.5005
R9142 VSS.n187 VSS.n104 4.5005
R9143 VSS.n201 VSS.n104 4.5005
R9144 VSS.n186 VSS.n104 4.5005
R9145 VSS.n202 VSS.n104 4.5005
R9146 VSS.n185 VSS.n104 4.5005
R9147 VSS.n203 VSS.n104 4.5005
R9148 VSS.n184 VSS.n104 4.5005
R9149 VSS.n204 VSS.n104 4.5005
R9150 VSS.n183 VSS.n104 4.5005
R9151 VSS.n205 VSS.n104 4.5005
R9152 VSS.n182 VSS.n104 4.5005
R9153 VSS.n206 VSS.n104 4.5005
R9154 VSS.n181 VSS.n104 4.5005
R9155 VSS.n207 VSS.n104 4.5005
R9156 VSS.n180 VSS.n104 4.5005
R9157 VSS.n208 VSS.n104 4.5005
R9158 VSS.n179 VSS.n104 4.5005
R9159 VSS.n209 VSS.n104 4.5005
R9160 VSS.n178 VSS.n104 4.5005
R9161 VSS.n210 VSS.n104 4.5005
R9162 VSS.n177 VSS.n104 4.5005
R9163 VSS.n211 VSS.n104 4.5005
R9164 VSS.n176 VSS.n104 4.5005
R9165 VSS.n212 VSS.n104 4.5005
R9166 VSS.n175 VSS.n104 4.5005
R9167 VSS.n213 VSS.n104 4.5005
R9168 VSS.n174 VSS.n104 4.5005
R9169 VSS.n214 VSS.n104 4.5005
R9170 VSS.n173 VSS.n104 4.5005
R9171 VSS.n215 VSS.n104 4.5005
R9172 VSS.n172 VSS.n104 4.5005
R9173 VSS.n216 VSS.n104 4.5005
R9174 VSS.n171 VSS.n104 4.5005
R9175 VSS.n217 VSS.n104 4.5005
R9176 VSS.n170 VSS.n104 4.5005
R9177 VSS.n218 VSS.n104 4.5005
R9178 VSS.n169 VSS.n104 4.5005
R9179 VSS.n219 VSS.n104 4.5005
R9180 VSS.n168 VSS.n104 4.5005
R9181 VSS.n220 VSS.n104 4.5005
R9182 VSS.n167 VSS.n104 4.5005
R9183 VSS.n221 VSS.n104 4.5005
R9184 VSS.n166 VSS.n104 4.5005
R9185 VSS.n222 VSS.n104 4.5005
R9186 VSS.n165 VSS.n104 4.5005
R9187 VSS.n223 VSS.n104 4.5005
R9188 VSS.n164 VSS.n104 4.5005
R9189 VSS.n224 VSS.n104 4.5005
R9190 VSS.n163 VSS.n104 4.5005
R9191 VSS.n225 VSS.n104 4.5005
R9192 VSS.n162 VSS.n104 4.5005
R9193 VSS.n226 VSS.n104 4.5005
R9194 VSS.n161 VSS.n104 4.5005
R9195 VSS.n227 VSS.n104 4.5005
R9196 VSS.n160 VSS.n104 4.5005
R9197 VSS.n228 VSS.n104 4.5005
R9198 VSS.n159 VSS.n104 4.5005
R9199 VSS.n229 VSS.n104 4.5005
R9200 VSS.n158 VSS.n104 4.5005
R9201 VSS.n230 VSS.n104 4.5005
R9202 VSS.n157 VSS.n104 4.5005
R9203 VSS.n231 VSS.n104 4.5005
R9204 VSS.n156 VSS.n104 4.5005
R9205 VSS.n232 VSS.n104 4.5005
R9206 VSS.n155 VSS.n104 4.5005
R9207 VSS.n233 VSS.n104 4.5005
R9208 VSS.n154 VSS.n104 4.5005
R9209 VSS.n234 VSS.n104 4.5005
R9210 VSS.n153 VSS.n104 4.5005
R9211 VSS.n235 VSS.n104 4.5005
R9212 VSS.n4506 VSS.n104 4.5005
R9213 VSS.n236 VSS.n104 4.5005
R9214 VSS.n152 VSS.n104 4.5005
R9215 VSS.n237 VSS.n104 4.5005
R9216 VSS.n151 VSS.n104 4.5005
R9217 VSS.n238 VSS.n104 4.5005
R9218 VSS.n150 VSS.n104 4.5005
R9219 VSS.n239 VSS.n104 4.5005
R9220 VSS.n149 VSS.n104 4.5005
R9221 VSS.n240 VSS.n104 4.5005
R9222 VSS.n148 VSS.n104 4.5005
R9223 VSS.n241 VSS.n104 4.5005
R9224 VSS.n147 VSS.n104 4.5005
R9225 VSS.n242 VSS.n104 4.5005
R9226 VSS.n146 VSS.n104 4.5005
R9227 VSS.n243 VSS.n104 4.5005
R9228 VSS.n145 VSS.n104 4.5005
R9229 VSS.n244 VSS.n104 4.5005
R9230 VSS.n144 VSS.n104 4.5005
R9231 VSS.n245 VSS.n104 4.5005
R9232 VSS.n143 VSS.n104 4.5005
R9233 VSS.n246 VSS.n104 4.5005
R9234 VSS.n142 VSS.n104 4.5005
R9235 VSS.n247 VSS.n104 4.5005
R9236 VSS.n141 VSS.n104 4.5005
R9237 VSS.n248 VSS.n104 4.5005
R9238 VSS.n140 VSS.n104 4.5005
R9239 VSS.n249 VSS.n104 4.5005
R9240 VSS.n139 VSS.n104 4.5005
R9241 VSS.n250 VSS.n104 4.5005
R9242 VSS.n138 VSS.n104 4.5005
R9243 VSS.n251 VSS.n104 4.5005
R9244 VSS.n137 VSS.n104 4.5005
R9245 VSS.n252 VSS.n104 4.5005
R9246 VSS.n136 VSS.n104 4.5005
R9247 VSS.n253 VSS.n104 4.5005
R9248 VSS.n135 VSS.n104 4.5005
R9249 VSS.n254 VSS.n104 4.5005
R9250 VSS.n134 VSS.n104 4.5005
R9251 VSS.n255 VSS.n104 4.5005
R9252 VSS.n133 VSS.n104 4.5005
R9253 VSS.n256 VSS.n104 4.5005
R9254 VSS.n132 VSS.n104 4.5005
R9255 VSS.n4502 VSS.n104 4.5005
R9256 VSS.n4504 VSS.n104 4.5005
R9257 VSS.n193 VSS.n32 4.5005
R9258 VSS.n195 VSS.n32 4.5005
R9259 VSS.n192 VSS.n32 4.5005
R9260 VSS.n196 VSS.n32 4.5005
R9261 VSS.n191 VSS.n32 4.5005
R9262 VSS.n197 VSS.n32 4.5005
R9263 VSS.n190 VSS.n32 4.5005
R9264 VSS.n198 VSS.n32 4.5005
R9265 VSS.n189 VSS.n32 4.5005
R9266 VSS.n199 VSS.n32 4.5005
R9267 VSS.n188 VSS.n32 4.5005
R9268 VSS.n200 VSS.n32 4.5005
R9269 VSS.n187 VSS.n32 4.5005
R9270 VSS.n201 VSS.n32 4.5005
R9271 VSS.n186 VSS.n32 4.5005
R9272 VSS.n202 VSS.n32 4.5005
R9273 VSS.n185 VSS.n32 4.5005
R9274 VSS.n203 VSS.n32 4.5005
R9275 VSS.n184 VSS.n32 4.5005
R9276 VSS.n204 VSS.n32 4.5005
R9277 VSS.n183 VSS.n32 4.5005
R9278 VSS.n205 VSS.n32 4.5005
R9279 VSS.n182 VSS.n32 4.5005
R9280 VSS.n206 VSS.n32 4.5005
R9281 VSS.n181 VSS.n32 4.5005
R9282 VSS.n207 VSS.n32 4.5005
R9283 VSS.n180 VSS.n32 4.5005
R9284 VSS.n208 VSS.n32 4.5005
R9285 VSS.n179 VSS.n32 4.5005
R9286 VSS.n209 VSS.n32 4.5005
R9287 VSS.n178 VSS.n32 4.5005
R9288 VSS.n210 VSS.n32 4.5005
R9289 VSS.n177 VSS.n32 4.5005
R9290 VSS.n211 VSS.n32 4.5005
R9291 VSS.n176 VSS.n32 4.5005
R9292 VSS.n212 VSS.n32 4.5005
R9293 VSS.n175 VSS.n32 4.5005
R9294 VSS.n213 VSS.n32 4.5005
R9295 VSS.n174 VSS.n32 4.5005
R9296 VSS.n214 VSS.n32 4.5005
R9297 VSS.n173 VSS.n32 4.5005
R9298 VSS.n215 VSS.n32 4.5005
R9299 VSS.n172 VSS.n32 4.5005
R9300 VSS.n216 VSS.n32 4.5005
R9301 VSS.n171 VSS.n32 4.5005
R9302 VSS.n217 VSS.n32 4.5005
R9303 VSS.n170 VSS.n32 4.5005
R9304 VSS.n218 VSS.n32 4.5005
R9305 VSS.n169 VSS.n32 4.5005
R9306 VSS.n219 VSS.n32 4.5005
R9307 VSS.n168 VSS.n32 4.5005
R9308 VSS.n220 VSS.n32 4.5005
R9309 VSS.n167 VSS.n32 4.5005
R9310 VSS.n221 VSS.n32 4.5005
R9311 VSS.n166 VSS.n32 4.5005
R9312 VSS.n222 VSS.n32 4.5005
R9313 VSS.n165 VSS.n32 4.5005
R9314 VSS.n223 VSS.n32 4.5005
R9315 VSS.n164 VSS.n32 4.5005
R9316 VSS.n224 VSS.n32 4.5005
R9317 VSS.n163 VSS.n32 4.5005
R9318 VSS.n225 VSS.n32 4.5005
R9319 VSS.n162 VSS.n32 4.5005
R9320 VSS.n226 VSS.n32 4.5005
R9321 VSS.n161 VSS.n32 4.5005
R9322 VSS.n227 VSS.n32 4.5005
R9323 VSS.n160 VSS.n32 4.5005
R9324 VSS.n228 VSS.n32 4.5005
R9325 VSS.n159 VSS.n32 4.5005
R9326 VSS.n229 VSS.n32 4.5005
R9327 VSS.n158 VSS.n32 4.5005
R9328 VSS.n230 VSS.n32 4.5005
R9329 VSS.n157 VSS.n32 4.5005
R9330 VSS.n231 VSS.n32 4.5005
R9331 VSS.n156 VSS.n32 4.5005
R9332 VSS.n232 VSS.n32 4.5005
R9333 VSS.n155 VSS.n32 4.5005
R9334 VSS.n233 VSS.n32 4.5005
R9335 VSS.n154 VSS.n32 4.5005
R9336 VSS.n234 VSS.n32 4.5005
R9337 VSS.n153 VSS.n32 4.5005
R9338 VSS.n235 VSS.n32 4.5005
R9339 VSS.n4506 VSS.n32 4.5005
R9340 VSS.n236 VSS.n32 4.5005
R9341 VSS.n152 VSS.n32 4.5005
R9342 VSS.n237 VSS.n32 4.5005
R9343 VSS.n151 VSS.n32 4.5005
R9344 VSS.n238 VSS.n32 4.5005
R9345 VSS.n150 VSS.n32 4.5005
R9346 VSS.n239 VSS.n32 4.5005
R9347 VSS.n149 VSS.n32 4.5005
R9348 VSS.n240 VSS.n32 4.5005
R9349 VSS.n148 VSS.n32 4.5005
R9350 VSS.n241 VSS.n32 4.5005
R9351 VSS.n147 VSS.n32 4.5005
R9352 VSS.n242 VSS.n32 4.5005
R9353 VSS.n146 VSS.n32 4.5005
R9354 VSS.n243 VSS.n32 4.5005
R9355 VSS.n145 VSS.n32 4.5005
R9356 VSS.n244 VSS.n32 4.5005
R9357 VSS.n144 VSS.n32 4.5005
R9358 VSS.n245 VSS.n32 4.5005
R9359 VSS.n143 VSS.n32 4.5005
R9360 VSS.n246 VSS.n32 4.5005
R9361 VSS.n142 VSS.n32 4.5005
R9362 VSS.n247 VSS.n32 4.5005
R9363 VSS.n141 VSS.n32 4.5005
R9364 VSS.n248 VSS.n32 4.5005
R9365 VSS.n140 VSS.n32 4.5005
R9366 VSS.n249 VSS.n32 4.5005
R9367 VSS.n139 VSS.n32 4.5005
R9368 VSS.n250 VSS.n32 4.5005
R9369 VSS.n138 VSS.n32 4.5005
R9370 VSS.n251 VSS.n32 4.5005
R9371 VSS.n137 VSS.n32 4.5005
R9372 VSS.n252 VSS.n32 4.5005
R9373 VSS.n136 VSS.n32 4.5005
R9374 VSS.n253 VSS.n32 4.5005
R9375 VSS.n135 VSS.n32 4.5005
R9376 VSS.n254 VSS.n32 4.5005
R9377 VSS.n134 VSS.n32 4.5005
R9378 VSS.n255 VSS.n32 4.5005
R9379 VSS.n133 VSS.n32 4.5005
R9380 VSS.n256 VSS.n32 4.5005
R9381 VSS.n132 VSS.n32 4.5005
R9382 VSS.n4502 VSS.n32 4.5005
R9383 VSS.n4504 VSS.n32 4.5005
R9384 VSS.n193 VSS.n105 4.5005
R9385 VSS.n195 VSS.n105 4.5005
R9386 VSS.n192 VSS.n105 4.5005
R9387 VSS.n196 VSS.n105 4.5005
R9388 VSS.n191 VSS.n105 4.5005
R9389 VSS.n197 VSS.n105 4.5005
R9390 VSS.n190 VSS.n105 4.5005
R9391 VSS.n198 VSS.n105 4.5005
R9392 VSS.n189 VSS.n105 4.5005
R9393 VSS.n199 VSS.n105 4.5005
R9394 VSS.n188 VSS.n105 4.5005
R9395 VSS.n200 VSS.n105 4.5005
R9396 VSS.n187 VSS.n105 4.5005
R9397 VSS.n201 VSS.n105 4.5005
R9398 VSS.n186 VSS.n105 4.5005
R9399 VSS.n202 VSS.n105 4.5005
R9400 VSS.n185 VSS.n105 4.5005
R9401 VSS.n203 VSS.n105 4.5005
R9402 VSS.n184 VSS.n105 4.5005
R9403 VSS.n204 VSS.n105 4.5005
R9404 VSS.n183 VSS.n105 4.5005
R9405 VSS.n205 VSS.n105 4.5005
R9406 VSS.n182 VSS.n105 4.5005
R9407 VSS.n206 VSS.n105 4.5005
R9408 VSS.n181 VSS.n105 4.5005
R9409 VSS.n207 VSS.n105 4.5005
R9410 VSS.n180 VSS.n105 4.5005
R9411 VSS.n208 VSS.n105 4.5005
R9412 VSS.n179 VSS.n105 4.5005
R9413 VSS.n209 VSS.n105 4.5005
R9414 VSS.n178 VSS.n105 4.5005
R9415 VSS.n210 VSS.n105 4.5005
R9416 VSS.n177 VSS.n105 4.5005
R9417 VSS.n211 VSS.n105 4.5005
R9418 VSS.n176 VSS.n105 4.5005
R9419 VSS.n212 VSS.n105 4.5005
R9420 VSS.n175 VSS.n105 4.5005
R9421 VSS.n213 VSS.n105 4.5005
R9422 VSS.n174 VSS.n105 4.5005
R9423 VSS.n214 VSS.n105 4.5005
R9424 VSS.n173 VSS.n105 4.5005
R9425 VSS.n215 VSS.n105 4.5005
R9426 VSS.n172 VSS.n105 4.5005
R9427 VSS.n216 VSS.n105 4.5005
R9428 VSS.n171 VSS.n105 4.5005
R9429 VSS.n217 VSS.n105 4.5005
R9430 VSS.n170 VSS.n105 4.5005
R9431 VSS.n218 VSS.n105 4.5005
R9432 VSS.n169 VSS.n105 4.5005
R9433 VSS.n219 VSS.n105 4.5005
R9434 VSS.n168 VSS.n105 4.5005
R9435 VSS.n220 VSS.n105 4.5005
R9436 VSS.n167 VSS.n105 4.5005
R9437 VSS.n221 VSS.n105 4.5005
R9438 VSS.n166 VSS.n105 4.5005
R9439 VSS.n222 VSS.n105 4.5005
R9440 VSS.n165 VSS.n105 4.5005
R9441 VSS.n223 VSS.n105 4.5005
R9442 VSS.n164 VSS.n105 4.5005
R9443 VSS.n224 VSS.n105 4.5005
R9444 VSS.n163 VSS.n105 4.5005
R9445 VSS.n225 VSS.n105 4.5005
R9446 VSS.n162 VSS.n105 4.5005
R9447 VSS.n226 VSS.n105 4.5005
R9448 VSS.n161 VSS.n105 4.5005
R9449 VSS.n227 VSS.n105 4.5005
R9450 VSS.n160 VSS.n105 4.5005
R9451 VSS.n228 VSS.n105 4.5005
R9452 VSS.n159 VSS.n105 4.5005
R9453 VSS.n229 VSS.n105 4.5005
R9454 VSS.n158 VSS.n105 4.5005
R9455 VSS.n230 VSS.n105 4.5005
R9456 VSS.n157 VSS.n105 4.5005
R9457 VSS.n231 VSS.n105 4.5005
R9458 VSS.n156 VSS.n105 4.5005
R9459 VSS.n232 VSS.n105 4.5005
R9460 VSS.n155 VSS.n105 4.5005
R9461 VSS.n233 VSS.n105 4.5005
R9462 VSS.n154 VSS.n105 4.5005
R9463 VSS.n234 VSS.n105 4.5005
R9464 VSS.n153 VSS.n105 4.5005
R9465 VSS.n235 VSS.n105 4.5005
R9466 VSS.n4506 VSS.n105 4.5005
R9467 VSS.n236 VSS.n105 4.5005
R9468 VSS.n152 VSS.n105 4.5005
R9469 VSS.n237 VSS.n105 4.5005
R9470 VSS.n151 VSS.n105 4.5005
R9471 VSS.n238 VSS.n105 4.5005
R9472 VSS.n150 VSS.n105 4.5005
R9473 VSS.n239 VSS.n105 4.5005
R9474 VSS.n149 VSS.n105 4.5005
R9475 VSS.n240 VSS.n105 4.5005
R9476 VSS.n148 VSS.n105 4.5005
R9477 VSS.n241 VSS.n105 4.5005
R9478 VSS.n147 VSS.n105 4.5005
R9479 VSS.n242 VSS.n105 4.5005
R9480 VSS.n146 VSS.n105 4.5005
R9481 VSS.n243 VSS.n105 4.5005
R9482 VSS.n145 VSS.n105 4.5005
R9483 VSS.n244 VSS.n105 4.5005
R9484 VSS.n144 VSS.n105 4.5005
R9485 VSS.n245 VSS.n105 4.5005
R9486 VSS.n143 VSS.n105 4.5005
R9487 VSS.n246 VSS.n105 4.5005
R9488 VSS.n142 VSS.n105 4.5005
R9489 VSS.n247 VSS.n105 4.5005
R9490 VSS.n141 VSS.n105 4.5005
R9491 VSS.n248 VSS.n105 4.5005
R9492 VSS.n140 VSS.n105 4.5005
R9493 VSS.n249 VSS.n105 4.5005
R9494 VSS.n139 VSS.n105 4.5005
R9495 VSS.n250 VSS.n105 4.5005
R9496 VSS.n138 VSS.n105 4.5005
R9497 VSS.n251 VSS.n105 4.5005
R9498 VSS.n137 VSS.n105 4.5005
R9499 VSS.n252 VSS.n105 4.5005
R9500 VSS.n136 VSS.n105 4.5005
R9501 VSS.n253 VSS.n105 4.5005
R9502 VSS.n135 VSS.n105 4.5005
R9503 VSS.n254 VSS.n105 4.5005
R9504 VSS.n134 VSS.n105 4.5005
R9505 VSS.n255 VSS.n105 4.5005
R9506 VSS.n133 VSS.n105 4.5005
R9507 VSS.n256 VSS.n105 4.5005
R9508 VSS.n132 VSS.n105 4.5005
R9509 VSS.n4502 VSS.n105 4.5005
R9510 VSS.n4504 VSS.n105 4.5005
R9511 VSS.n193 VSS.n31 4.5005
R9512 VSS.n195 VSS.n31 4.5005
R9513 VSS.n192 VSS.n31 4.5005
R9514 VSS.n196 VSS.n31 4.5005
R9515 VSS.n191 VSS.n31 4.5005
R9516 VSS.n197 VSS.n31 4.5005
R9517 VSS.n190 VSS.n31 4.5005
R9518 VSS.n198 VSS.n31 4.5005
R9519 VSS.n189 VSS.n31 4.5005
R9520 VSS.n199 VSS.n31 4.5005
R9521 VSS.n188 VSS.n31 4.5005
R9522 VSS.n200 VSS.n31 4.5005
R9523 VSS.n187 VSS.n31 4.5005
R9524 VSS.n201 VSS.n31 4.5005
R9525 VSS.n186 VSS.n31 4.5005
R9526 VSS.n202 VSS.n31 4.5005
R9527 VSS.n185 VSS.n31 4.5005
R9528 VSS.n203 VSS.n31 4.5005
R9529 VSS.n184 VSS.n31 4.5005
R9530 VSS.n204 VSS.n31 4.5005
R9531 VSS.n183 VSS.n31 4.5005
R9532 VSS.n205 VSS.n31 4.5005
R9533 VSS.n182 VSS.n31 4.5005
R9534 VSS.n206 VSS.n31 4.5005
R9535 VSS.n181 VSS.n31 4.5005
R9536 VSS.n207 VSS.n31 4.5005
R9537 VSS.n180 VSS.n31 4.5005
R9538 VSS.n208 VSS.n31 4.5005
R9539 VSS.n179 VSS.n31 4.5005
R9540 VSS.n209 VSS.n31 4.5005
R9541 VSS.n178 VSS.n31 4.5005
R9542 VSS.n210 VSS.n31 4.5005
R9543 VSS.n177 VSS.n31 4.5005
R9544 VSS.n211 VSS.n31 4.5005
R9545 VSS.n176 VSS.n31 4.5005
R9546 VSS.n212 VSS.n31 4.5005
R9547 VSS.n175 VSS.n31 4.5005
R9548 VSS.n213 VSS.n31 4.5005
R9549 VSS.n174 VSS.n31 4.5005
R9550 VSS.n214 VSS.n31 4.5005
R9551 VSS.n173 VSS.n31 4.5005
R9552 VSS.n215 VSS.n31 4.5005
R9553 VSS.n172 VSS.n31 4.5005
R9554 VSS.n216 VSS.n31 4.5005
R9555 VSS.n171 VSS.n31 4.5005
R9556 VSS.n217 VSS.n31 4.5005
R9557 VSS.n170 VSS.n31 4.5005
R9558 VSS.n218 VSS.n31 4.5005
R9559 VSS.n169 VSS.n31 4.5005
R9560 VSS.n219 VSS.n31 4.5005
R9561 VSS.n168 VSS.n31 4.5005
R9562 VSS.n220 VSS.n31 4.5005
R9563 VSS.n167 VSS.n31 4.5005
R9564 VSS.n221 VSS.n31 4.5005
R9565 VSS.n166 VSS.n31 4.5005
R9566 VSS.n222 VSS.n31 4.5005
R9567 VSS.n165 VSS.n31 4.5005
R9568 VSS.n223 VSS.n31 4.5005
R9569 VSS.n164 VSS.n31 4.5005
R9570 VSS.n224 VSS.n31 4.5005
R9571 VSS.n163 VSS.n31 4.5005
R9572 VSS.n225 VSS.n31 4.5005
R9573 VSS.n162 VSS.n31 4.5005
R9574 VSS.n226 VSS.n31 4.5005
R9575 VSS.n161 VSS.n31 4.5005
R9576 VSS.n227 VSS.n31 4.5005
R9577 VSS.n160 VSS.n31 4.5005
R9578 VSS.n228 VSS.n31 4.5005
R9579 VSS.n159 VSS.n31 4.5005
R9580 VSS.n229 VSS.n31 4.5005
R9581 VSS.n158 VSS.n31 4.5005
R9582 VSS.n230 VSS.n31 4.5005
R9583 VSS.n157 VSS.n31 4.5005
R9584 VSS.n231 VSS.n31 4.5005
R9585 VSS.n156 VSS.n31 4.5005
R9586 VSS.n232 VSS.n31 4.5005
R9587 VSS.n155 VSS.n31 4.5005
R9588 VSS.n233 VSS.n31 4.5005
R9589 VSS.n154 VSS.n31 4.5005
R9590 VSS.n234 VSS.n31 4.5005
R9591 VSS.n153 VSS.n31 4.5005
R9592 VSS.n235 VSS.n31 4.5005
R9593 VSS.n4506 VSS.n31 4.5005
R9594 VSS.n236 VSS.n31 4.5005
R9595 VSS.n152 VSS.n31 4.5005
R9596 VSS.n237 VSS.n31 4.5005
R9597 VSS.n151 VSS.n31 4.5005
R9598 VSS.n238 VSS.n31 4.5005
R9599 VSS.n150 VSS.n31 4.5005
R9600 VSS.n239 VSS.n31 4.5005
R9601 VSS.n149 VSS.n31 4.5005
R9602 VSS.n240 VSS.n31 4.5005
R9603 VSS.n148 VSS.n31 4.5005
R9604 VSS.n241 VSS.n31 4.5005
R9605 VSS.n147 VSS.n31 4.5005
R9606 VSS.n242 VSS.n31 4.5005
R9607 VSS.n146 VSS.n31 4.5005
R9608 VSS.n243 VSS.n31 4.5005
R9609 VSS.n145 VSS.n31 4.5005
R9610 VSS.n244 VSS.n31 4.5005
R9611 VSS.n144 VSS.n31 4.5005
R9612 VSS.n245 VSS.n31 4.5005
R9613 VSS.n143 VSS.n31 4.5005
R9614 VSS.n246 VSS.n31 4.5005
R9615 VSS.n142 VSS.n31 4.5005
R9616 VSS.n247 VSS.n31 4.5005
R9617 VSS.n141 VSS.n31 4.5005
R9618 VSS.n248 VSS.n31 4.5005
R9619 VSS.n140 VSS.n31 4.5005
R9620 VSS.n249 VSS.n31 4.5005
R9621 VSS.n139 VSS.n31 4.5005
R9622 VSS.n250 VSS.n31 4.5005
R9623 VSS.n138 VSS.n31 4.5005
R9624 VSS.n251 VSS.n31 4.5005
R9625 VSS.n137 VSS.n31 4.5005
R9626 VSS.n252 VSS.n31 4.5005
R9627 VSS.n136 VSS.n31 4.5005
R9628 VSS.n253 VSS.n31 4.5005
R9629 VSS.n135 VSS.n31 4.5005
R9630 VSS.n254 VSS.n31 4.5005
R9631 VSS.n134 VSS.n31 4.5005
R9632 VSS.n255 VSS.n31 4.5005
R9633 VSS.n133 VSS.n31 4.5005
R9634 VSS.n256 VSS.n31 4.5005
R9635 VSS.n132 VSS.n31 4.5005
R9636 VSS.n4502 VSS.n31 4.5005
R9637 VSS.n4504 VSS.n31 4.5005
R9638 VSS.n193 VSS.n106 4.5005
R9639 VSS.n195 VSS.n106 4.5005
R9640 VSS.n192 VSS.n106 4.5005
R9641 VSS.n196 VSS.n106 4.5005
R9642 VSS.n191 VSS.n106 4.5005
R9643 VSS.n197 VSS.n106 4.5005
R9644 VSS.n190 VSS.n106 4.5005
R9645 VSS.n198 VSS.n106 4.5005
R9646 VSS.n189 VSS.n106 4.5005
R9647 VSS.n199 VSS.n106 4.5005
R9648 VSS.n188 VSS.n106 4.5005
R9649 VSS.n200 VSS.n106 4.5005
R9650 VSS.n187 VSS.n106 4.5005
R9651 VSS.n201 VSS.n106 4.5005
R9652 VSS.n186 VSS.n106 4.5005
R9653 VSS.n202 VSS.n106 4.5005
R9654 VSS.n185 VSS.n106 4.5005
R9655 VSS.n203 VSS.n106 4.5005
R9656 VSS.n184 VSS.n106 4.5005
R9657 VSS.n204 VSS.n106 4.5005
R9658 VSS.n183 VSS.n106 4.5005
R9659 VSS.n205 VSS.n106 4.5005
R9660 VSS.n182 VSS.n106 4.5005
R9661 VSS.n206 VSS.n106 4.5005
R9662 VSS.n181 VSS.n106 4.5005
R9663 VSS.n207 VSS.n106 4.5005
R9664 VSS.n180 VSS.n106 4.5005
R9665 VSS.n208 VSS.n106 4.5005
R9666 VSS.n179 VSS.n106 4.5005
R9667 VSS.n209 VSS.n106 4.5005
R9668 VSS.n178 VSS.n106 4.5005
R9669 VSS.n210 VSS.n106 4.5005
R9670 VSS.n177 VSS.n106 4.5005
R9671 VSS.n211 VSS.n106 4.5005
R9672 VSS.n176 VSS.n106 4.5005
R9673 VSS.n212 VSS.n106 4.5005
R9674 VSS.n175 VSS.n106 4.5005
R9675 VSS.n213 VSS.n106 4.5005
R9676 VSS.n174 VSS.n106 4.5005
R9677 VSS.n214 VSS.n106 4.5005
R9678 VSS.n173 VSS.n106 4.5005
R9679 VSS.n215 VSS.n106 4.5005
R9680 VSS.n172 VSS.n106 4.5005
R9681 VSS.n216 VSS.n106 4.5005
R9682 VSS.n171 VSS.n106 4.5005
R9683 VSS.n217 VSS.n106 4.5005
R9684 VSS.n170 VSS.n106 4.5005
R9685 VSS.n218 VSS.n106 4.5005
R9686 VSS.n169 VSS.n106 4.5005
R9687 VSS.n219 VSS.n106 4.5005
R9688 VSS.n168 VSS.n106 4.5005
R9689 VSS.n220 VSS.n106 4.5005
R9690 VSS.n167 VSS.n106 4.5005
R9691 VSS.n221 VSS.n106 4.5005
R9692 VSS.n166 VSS.n106 4.5005
R9693 VSS.n222 VSS.n106 4.5005
R9694 VSS.n165 VSS.n106 4.5005
R9695 VSS.n223 VSS.n106 4.5005
R9696 VSS.n164 VSS.n106 4.5005
R9697 VSS.n224 VSS.n106 4.5005
R9698 VSS.n163 VSS.n106 4.5005
R9699 VSS.n225 VSS.n106 4.5005
R9700 VSS.n162 VSS.n106 4.5005
R9701 VSS.n226 VSS.n106 4.5005
R9702 VSS.n161 VSS.n106 4.5005
R9703 VSS.n227 VSS.n106 4.5005
R9704 VSS.n160 VSS.n106 4.5005
R9705 VSS.n228 VSS.n106 4.5005
R9706 VSS.n159 VSS.n106 4.5005
R9707 VSS.n229 VSS.n106 4.5005
R9708 VSS.n158 VSS.n106 4.5005
R9709 VSS.n230 VSS.n106 4.5005
R9710 VSS.n157 VSS.n106 4.5005
R9711 VSS.n231 VSS.n106 4.5005
R9712 VSS.n156 VSS.n106 4.5005
R9713 VSS.n232 VSS.n106 4.5005
R9714 VSS.n155 VSS.n106 4.5005
R9715 VSS.n233 VSS.n106 4.5005
R9716 VSS.n154 VSS.n106 4.5005
R9717 VSS.n234 VSS.n106 4.5005
R9718 VSS.n153 VSS.n106 4.5005
R9719 VSS.n235 VSS.n106 4.5005
R9720 VSS.n4506 VSS.n106 4.5005
R9721 VSS.n236 VSS.n106 4.5005
R9722 VSS.n152 VSS.n106 4.5005
R9723 VSS.n237 VSS.n106 4.5005
R9724 VSS.n151 VSS.n106 4.5005
R9725 VSS.n238 VSS.n106 4.5005
R9726 VSS.n150 VSS.n106 4.5005
R9727 VSS.n239 VSS.n106 4.5005
R9728 VSS.n149 VSS.n106 4.5005
R9729 VSS.n240 VSS.n106 4.5005
R9730 VSS.n148 VSS.n106 4.5005
R9731 VSS.n241 VSS.n106 4.5005
R9732 VSS.n147 VSS.n106 4.5005
R9733 VSS.n242 VSS.n106 4.5005
R9734 VSS.n146 VSS.n106 4.5005
R9735 VSS.n243 VSS.n106 4.5005
R9736 VSS.n145 VSS.n106 4.5005
R9737 VSS.n244 VSS.n106 4.5005
R9738 VSS.n144 VSS.n106 4.5005
R9739 VSS.n245 VSS.n106 4.5005
R9740 VSS.n143 VSS.n106 4.5005
R9741 VSS.n246 VSS.n106 4.5005
R9742 VSS.n142 VSS.n106 4.5005
R9743 VSS.n247 VSS.n106 4.5005
R9744 VSS.n141 VSS.n106 4.5005
R9745 VSS.n248 VSS.n106 4.5005
R9746 VSS.n140 VSS.n106 4.5005
R9747 VSS.n249 VSS.n106 4.5005
R9748 VSS.n139 VSS.n106 4.5005
R9749 VSS.n250 VSS.n106 4.5005
R9750 VSS.n138 VSS.n106 4.5005
R9751 VSS.n251 VSS.n106 4.5005
R9752 VSS.n137 VSS.n106 4.5005
R9753 VSS.n252 VSS.n106 4.5005
R9754 VSS.n136 VSS.n106 4.5005
R9755 VSS.n253 VSS.n106 4.5005
R9756 VSS.n135 VSS.n106 4.5005
R9757 VSS.n254 VSS.n106 4.5005
R9758 VSS.n134 VSS.n106 4.5005
R9759 VSS.n255 VSS.n106 4.5005
R9760 VSS.n133 VSS.n106 4.5005
R9761 VSS.n256 VSS.n106 4.5005
R9762 VSS.n132 VSS.n106 4.5005
R9763 VSS.n4502 VSS.n106 4.5005
R9764 VSS.n4504 VSS.n106 4.5005
R9765 VSS.n193 VSS.n30 4.5005
R9766 VSS.n195 VSS.n30 4.5005
R9767 VSS.n192 VSS.n30 4.5005
R9768 VSS.n196 VSS.n30 4.5005
R9769 VSS.n191 VSS.n30 4.5005
R9770 VSS.n197 VSS.n30 4.5005
R9771 VSS.n190 VSS.n30 4.5005
R9772 VSS.n198 VSS.n30 4.5005
R9773 VSS.n189 VSS.n30 4.5005
R9774 VSS.n199 VSS.n30 4.5005
R9775 VSS.n188 VSS.n30 4.5005
R9776 VSS.n200 VSS.n30 4.5005
R9777 VSS.n187 VSS.n30 4.5005
R9778 VSS.n201 VSS.n30 4.5005
R9779 VSS.n186 VSS.n30 4.5005
R9780 VSS.n202 VSS.n30 4.5005
R9781 VSS.n185 VSS.n30 4.5005
R9782 VSS.n203 VSS.n30 4.5005
R9783 VSS.n184 VSS.n30 4.5005
R9784 VSS.n204 VSS.n30 4.5005
R9785 VSS.n183 VSS.n30 4.5005
R9786 VSS.n205 VSS.n30 4.5005
R9787 VSS.n182 VSS.n30 4.5005
R9788 VSS.n206 VSS.n30 4.5005
R9789 VSS.n181 VSS.n30 4.5005
R9790 VSS.n207 VSS.n30 4.5005
R9791 VSS.n180 VSS.n30 4.5005
R9792 VSS.n208 VSS.n30 4.5005
R9793 VSS.n179 VSS.n30 4.5005
R9794 VSS.n209 VSS.n30 4.5005
R9795 VSS.n178 VSS.n30 4.5005
R9796 VSS.n210 VSS.n30 4.5005
R9797 VSS.n177 VSS.n30 4.5005
R9798 VSS.n211 VSS.n30 4.5005
R9799 VSS.n176 VSS.n30 4.5005
R9800 VSS.n212 VSS.n30 4.5005
R9801 VSS.n175 VSS.n30 4.5005
R9802 VSS.n213 VSS.n30 4.5005
R9803 VSS.n174 VSS.n30 4.5005
R9804 VSS.n214 VSS.n30 4.5005
R9805 VSS.n173 VSS.n30 4.5005
R9806 VSS.n215 VSS.n30 4.5005
R9807 VSS.n172 VSS.n30 4.5005
R9808 VSS.n216 VSS.n30 4.5005
R9809 VSS.n171 VSS.n30 4.5005
R9810 VSS.n217 VSS.n30 4.5005
R9811 VSS.n170 VSS.n30 4.5005
R9812 VSS.n218 VSS.n30 4.5005
R9813 VSS.n169 VSS.n30 4.5005
R9814 VSS.n219 VSS.n30 4.5005
R9815 VSS.n168 VSS.n30 4.5005
R9816 VSS.n220 VSS.n30 4.5005
R9817 VSS.n167 VSS.n30 4.5005
R9818 VSS.n221 VSS.n30 4.5005
R9819 VSS.n166 VSS.n30 4.5005
R9820 VSS.n222 VSS.n30 4.5005
R9821 VSS.n165 VSS.n30 4.5005
R9822 VSS.n223 VSS.n30 4.5005
R9823 VSS.n164 VSS.n30 4.5005
R9824 VSS.n224 VSS.n30 4.5005
R9825 VSS.n163 VSS.n30 4.5005
R9826 VSS.n225 VSS.n30 4.5005
R9827 VSS.n162 VSS.n30 4.5005
R9828 VSS.n226 VSS.n30 4.5005
R9829 VSS.n161 VSS.n30 4.5005
R9830 VSS.n227 VSS.n30 4.5005
R9831 VSS.n160 VSS.n30 4.5005
R9832 VSS.n228 VSS.n30 4.5005
R9833 VSS.n159 VSS.n30 4.5005
R9834 VSS.n229 VSS.n30 4.5005
R9835 VSS.n158 VSS.n30 4.5005
R9836 VSS.n230 VSS.n30 4.5005
R9837 VSS.n157 VSS.n30 4.5005
R9838 VSS.n231 VSS.n30 4.5005
R9839 VSS.n156 VSS.n30 4.5005
R9840 VSS.n232 VSS.n30 4.5005
R9841 VSS.n155 VSS.n30 4.5005
R9842 VSS.n233 VSS.n30 4.5005
R9843 VSS.n154 VSS.n30 4.5005
R9844 VSS.n234 VSS.n30 4.5005
R9845 VSS.n153 VSS.n30 4.5005
R9846 VSS.n235 VSS.n30 4.5005
R9847 VSS.n4506 VSS.n30 4.5005
R9848 VSS.n236 VSS.n30 4.5005
R9849 VSS.n152 VSS.n30 4.5005
R9850 VSS.n237 VSS.n30 4.5005
R9851 VSS.n151 VSS.n30 4.5005
R9852 VSS.n238 VSS.n30 4.5005
R9853 VSS.n150 VSS.n30 4.5005
R9854 VSS.n239 VSS.n30 4.5005
R9855 VSS.n149 VSS.n30 4.5005
R9856 VSS.n240 VSS.n30 4.5005
R9857 VSS.n148 VSS.n30 4.5005
R9858 VSS.n241 VSS.n30 4.5005
R9859 VSS.n147 VSS.n30 4.5005
R9860 VSS.n242 VSS.n30 4.5005
R9861 VSS.n146 VSS.n30 4.5005
R9862 VSS.n243 VSS.n30 4.5005
R9863 VSS.n145 VSS.n30 4.5005
R9864 VSS.n244 VSS.n30 4.5005
R9865 VSS.n144 VSS.n30 4.5005
R9866 VSS.n245 VSS.n30 4.5005
R9867 VSS.n143 VSS.n30 4.5005
R9868 VSS.n246 VSS.n30 4.5005
R9869 VSS.n142 VSS.n30 4.5005
R9870 VSS.n247 VSS.n30 4.5005
R9871 VSS.n141 VSS.n30 4.5005
R9872 VSS.n248 VSS.n30 4.5005
R9873 VSS.n140 VSS.n30 4.5005
R9874 VSS.n249 VSS.n30 4.5005
R9875 VSS.n139 VSS.n30 4.5005
R9876 VSS.n250 VSS.n30 4.5005
R9877 VSS.n138 VSS.n30 4.5005
R9878 VSS.n251 VSS.n30 4.5005
R9879 VSS.n137 VSS.n30 4.5005
R9880 VSS.n252 VSS.n30 4.5005
R9881 VSS.n136 VSS.n30 4.5005
R9882 VSS.n253 VSS.n30 4.5005
R9883 VSS.n135 VSS.n30 4.5005
R9884 VSS.n254 VSS.n30 4.5005
R9885 VSS.n134 VSS.n30 4.5005
R9886 VSS.n255 VSS.n30 4.5005
R9887 VSS.n133 VSS.n30 4.5005
R9888 VSS.n256 VSS.n30 4.5005
R9889 VSS.n132 VSS.n30 4.5005
R9890 VSS.n4502 VSS.n30 4.5005
R9891 VSS.n4504 VSS.n30 4.5005
R9892 VSS.n193 VSS.n107 4.5005
R9893 VSS.n195 VSS.n107 4.5005
R9894 VSS.n192 VSS.n107 4.5005
R9895 VSS.n196 VSS.n107 4.5005
R9896 VSS.n191 VSS.n107 4.5005
R9897 VSS.n197 VSS.n107 4.5005
R9898 VSS.n190 VSS.n107 4.5005
R9899 VSS.n198 VSS.n107 4.5005
R9900 VSS.n189 VSS.n107 4.5005
R9901 VSS.n199 VSS.n107 4.5005
R9902 VSS.n188 VSS.n107 4.5005
R9903 VSS.n200 VSS.n107 4.5005
R9904 VSS.n187 VSS.n107 4.5005
R9905 VSS.n201 VSS.n107 4.5005
R9906 VSS.n186 VSS.n107 4.5005
R9907 VSS.n202 VSS.n107 4.5005
R9908 VSS.n185 VSS.n107 4.5005
R9909 VSS.n203 VSS.n107 4.5005
R9910 VSS.n184 VSS.n107 4.5005
R9911 VSS.n204 VSS.n107 4.5005
R9912 VSS.n183 VSS.n107 4.5005
R9913 VSS.n205 VSS.n107 4.5005
R9914 VSS.n182 VSS.n107 4.5005
R9915 VSS.n206 VSS.n107 4.5005
R9916 VSS.n181 VSS.n107 4.5005
R9917 VSS.n207 VSS.n107 4.5005
R9918 VSS.n180 VSS.n107 4.5005
R9919 VSS.n208 VSS.n107 4.5005
R9920 VSS.n179 VSS.n107 4.5005
R9921 VSS.n209 VSS.n107 4.5005
R9922 VSS.n178 VSS.n107 4.5005
R9923 VSS.n210 VSS.n107 4.5005
R9924 VSS.n177 VSS.n107 4.5005
R9925 VSS.n211 VSS.n107 4.5005
R9926 VSS.n176 VSS.n107 4.5005
R9927 VSS.n212 VSS.n107 4.5005
R9928 VSS.n175 VSS.n107 4.5005
R9929 VSS.n213 VSS.n107 4.5005
R9930 VSS.n174 VSS.n107 4.5005
R9931 VSS.n214 VSS.n107 4.5005
R9932 VSS.n173 VSS.n107 4.5005
R9933 VSS.n215 VSS.n107 4.5005
R9934 VSS.n172 VSS.n107 4.5005
R9935 VSS.n216 VSS.n107 4.5005
R9936 VSS.n171 VSS.n107 4.5005
R9937 VSS.n217 VSS.n107 4.5005
R9938 VSS.n170 VSS.n107 4.5005
R9939 VSS.n218 VSS.n107 4.5005
R9940 VSS.n169 VSS.n107 4.5005
R9941 VSS.n219 VSS.n107 4.5005
R9942 VSS.n168 VSS.n107 4.5005
R9943 VSS.n220 VSS.n107 4.5005
R9944 VSS.n167 VSS.n107 4.5005
R9945 VSS.n221 VSS.n107 4.5005
R9946 VSS.n166 VSS.n107 4.5005
R9947 VSS.n222 VSS.n107 4.5005
R9948 VSS.n165 VSS.n107 4.5005
R9949 VSS.n223 VSS.n107 4.5005
R9950 VSS.n164 VSS.n107 4.5005
R9951 VSS.n224 VSS.n107 4.5005
R9952 VSS.n163 VSS.n107 4.5005
R9953 VSS.n225 VSS.n107 4.5005
R9954 VSS.n162 VSS.n107 4.5005
R9955 VSS.n226 VSS.n107 4.5005
R9956 VSS.n161 VSS.n107 4.5005
R9957 VSS.n227 VSS.n107 4.5005
R9958 VSS.n160 VSS.n107 4.5005
R9959 VSS.n228 VSS.n107 4.5005
R9960 VSS.n159 VSS.n107 4.5005
R9961 VSS.n229 VSS.n107 4.5005
R9962 VSS.n158 VSS.n107 4.5005
R9963 VSS.n230 VSS.n107 4.5005
R9964 VSS.n157 VSS.n107 4.5005
R9965 VSS.n231 VSS.n107 4.5005
R9966 VSS.n156 VSS.n107 4.5005
R9967 VSS.n232 VSS.n107 4.5005
R9968 VSS.n155 VSS.n107 4.5005
R9969 VSS.n233 VSS.n107 4.5005
R9970 VSS.n154 VSS.n107 4.5005
R9971 VSS.n234 VSS.n107 4.5005
R9972 VSS.n153 VSS.n107 4.5005
R9973 VSS.n235 VSS.n107 4.5005
R9974 VSS.n4506 VSS.n107 4.5005
R9975 VSS.n236 VSS.n107 4.5005
R9976 VSS.n152 VSS.n107 4.5005
R9977 VSS.n237 VSS.n107 4.5005
R9978 VSS.n151 VSS.n107 4.5005
R9979 VSS.n238 VSS.n107 4.5005
R9980 VSS.n150 VSS.n107 4.5005
R9981 VSS.n239 VSS.n107 4.5005
R9982 VSS.n149 VSS.n107 4.5005
R9983 VSS.n240 VSS.n107 4.5005
R9984 VSS.n148 VSS.n107 4.5005
R9985 VSS.n241 VSS.n107 4.5005
R9986 VSS.n147 VSS.n107 4.5005
R9987 VSS.n242 VSS.n107 4.5005
R9988 VSS.n146 VSS.n107 4.5005
R9989 VSS.n243 VSS.n107 4.5005
R9990 VSS.n145 VSS.n107 4.5005
R9991 VSS.n244 VSS.n107 4.5005
R9992 VSS.n144 VSS.n107 4.5005
R9993 VSS.n245 VSS.n107 4.5005
R9994 VSS.n143 VSS.n107 4.5005
R9995 VSS.n246 VSS.n107 4.5005
R9996 VSS.n142 VSS.n107 4.5005
R9997 VSS.n247 VSS.n107 4.5005
R9998 VSS.n141 VSS.n107 4.5005
R9999 VSS.n248 VSS.n107 4.5005
R10000 VSS.n140 VSS.n107 4.5005
R10001 VSS.n249 VSS.n107 4.5005
R10002 VSS.n139 VSS.n107 4.5005
R10003 VSS.n250 VSS.n107 4.5005
R10004 VSS.n138 VSS.n107 4.5005
R10005 VSS.n251 VSS.n107 4.5005
R10006 VSS.n137 VSS.n107 4.5005
R10007 VSS.n252 VSS.n107 4.5005
R10008 VSS.n136 VSS.n107 4.5005
R10009 VSS.n253 VSS.n107 4.5005
R10010 VSS.n135 VSS.n107 4.5005
R10011 VSS.n254 VSS.n107 4.5005
R10012 VSS.n134 VSS.n107 4.5005
R10013 VSS.n255 VSS.n107 4.5005
R10014 VSS.n133 VSS.n107 4.5005
R10015 VSS.n256 VSS.n107 4.5005
R10016 VSS.n132 VSS.n107 4.5005
R10017 VSS.n4502 VSS.n107 4.5005
R10018 VSS.n4504 VSS.n107 4.5005
R10019 VSS.n193 VSS.n29 4.5005
R10020 VSS.n195 VSS.n29 4.5005
R10021 VSS.n192 VSS.n29 4.5005
R10022 VSS.n196 VSS.n29 4.5005
R10023 VSS.n191 VSS.n29 4.5005
R10024 VSS.n197 VSS.n29 4.5005
R10025 VSS.n190 VSS.n29 4.5005
R10026 VSS.n198 VSS.n29 4.5005
R10027 VSS.n189 VSS.n29 4.5005
R10028 VSS.n199 VSS.n29 4.5005
R10029 VSS.n188 VSS.n29 4.5005
R10030 VSS.n200 VSS.n29 4.5005
R10031 VSS.n187 VSS.n29 4.5005
R10032 VSS.n201 VSS.n29 4.5005
R10033 VSS.n186 VSS.n29 4.5005
R10034 VSS.n202 VSS.n29 4.5005
R10035 VSS.n185 VSS.n29 4.5005
R10036 VSS.n203 VSS.n29 4.5005
R10037 VSS.n184 VSS.n29 4.5005
R10038 VSS.n204 VSS.n29 4.5005
R10039 VSS.n183 VSS.n29 4.5005
R10040 VSS.n205 VSS.n29 4.5005
R10041 VSS.n182 VSS.n29 4.5005
R10042 VSS.n206 VSS.n29 4.5005
R10043 VSS.n181 VSS.n29 4.5005
R10044 VSS.n207 VSS.n29 4.5005
R10045 VSS.n180 VSS.n29 4.5005
R10046 VSS.n208 VSS.n29 4.5005
R10047 VSS.n179 VSS.n29 4.5005
R10048 VSS.n209 VSS.n29 4.5005
R10049 VSS.n178 VSS.n29 4.5005
R10050 VSS.n210 VSS.n29 4.5005
R10051 VSS.n177 VSS.n29 4.5005
R10052 VSS.n211 VSS.n29 4.5005
R10053 VSS.n176 VSS.n29 4.5005
R10054 VSS.n212 VSS.n29 4.5005
R10055 VSS.n175 VSS.n29 4.5005
R10056 VSS.n213 VSS.n29 4.5005
R10057 VSS.n174 VSS.n29 4.5005
R10058 VSS.n214 VSS.n29 4.5005
R10059 VSS.n173 VSS.n29 4.5005
R10060 VSS.n215 VSS.n29 4.5005
R10061 VSS.n172 VSS.n29 4.5005
R10062 VSS.n216 VSS.n29 4.5005
R10063 VSS.n171 VSS.n29 4.5005
R10064 VSS.n217 VSS.n29 4.5005
R10065 VSS.n170 VSS.n29 4.5005
R10066 VSS.n218 VSS.n29 4.5005
R10067 VSS.n169 VSS.n29 4.5005
R10068 VSS.n219 VSS.n29 4.5005
R10069 VSS.n168 VSS.n29 4.5005
R10070 VSS.n220 VSS.n29 4.5005
R10071 VSS.n167 VSS.n29 4.5005
R10072 VSS.n221 VSS.n29 4.5005
R10073 VSS.n166 VSS.n29 4.5005
R10074 VSS.n222 VSS.n29 4.5005
R10075 VSS.n165 VSS.n29 4.5005
R10076 VSS.n223 VSS.n29 4.5005
R10077 VSS.n164 VSS.n29 4.5005
R10078 VSS.n224 VSS.n29 4.5005
R10079 VSS.n163 VSS.n29 4.5005
R10080 VSS.n225 VSS.n29 4.5005
R10081 VSS.n162 VSS.n29 4.5005
R10082 VSS.n226 VSS.n29 4.5005
R10083 VSS.n161 VSS.n29 4.5005
R10084 VSS.n227 VSS.n29 4.5005
R10085 VSS.n160 VSS.n29 4.5005
R10086 VSS.n228 VSS.n29 4.5005
R10087 VSS.n159 VSS.n29 4.5005
R10088 VSS.n229 VSS.n29 4.5005
R10089 VSS.n158 VSS.n29 4.5005
R10090 VSS.n230 VSS.n29 4.5005
R10091 VSS.n157 VSS.n29 4.5005
R10092 VSS.n231 VSS.n29 4.5005
R10093 VSS.n156 VSS.n29 4.5005
R10094 VSS.n232 VSS.n29 4.5005
R10095 VSS.n155 VSS.n29 4.5005
R10096 VSS.n233 VSS.n29 4.5005
R10097 VSS.n154 VSS.n29 4.5005
R10098 VSS.n234 VSS.n29 4.5005
R10099 VSS.n153 VSS.n29 4.5005
R10100 VSS.n235 VSS.n29 4.5005
R10101 VSS.n4506 VSS.n29 4.5005
R10102 VSS.n236 VSS.n29 4.5005
R10103 VSS.n152 VSS.n29 4.5005
R10104 VSS.n237 VSS.n29 4.5005
R10105 VSS.n151 VSS.n29 4.5005
R10106 VSS.n238 VSS.n29 4.5005
R10107 VSS.n150 VSS.n29 4.5005
R10108 VSS.n239 VSS.n29 4.5005
R10109 VSS.n149 VSS.n29 4.5005
R10110 VSS.n240 VSS.n29 4.5005
R10111 VSS.n148 VSS.n29 4.5005
R10112 VSS.n241 VSS.n29 4.5005
R10113 VSS.n147 VSS.n29 4.5005
R10114 VSS.n242 VSS.n29 4.5005
R10115 VSS.n146 VSS.n29 4.5005
R10116 VSS.n243 VSS.n29 4.5005
R10117 VSS.n145 VSS.n29 4.5005
R10118 VSS.n244 VSS.n29 4.5005
R10119 VSS.n144 VSS.n29 4.5005
R10120 VSS.n245 VSS.n29 4.5005
R10121 VSS.n143 VSS.n29 4.5005
R10122 VSS.n246 VSS.n29 4.5005
R10123 VSS.n142 VSS.n29 4.5005
R10124 VSS.n247 VSS.n29 4.5005
R10125 VSS.n141 VSS.n29 4.5005
R10126 VSS.n248 VSS.n29 4.5005
R10127 VSS.n140 VSS.n29 4.5005
R10128 VSS.n249 VSS.n29 4.5005
R10129 VSS.n139 VSS.n29 4.5005
R10130 VSS.n250 VSS.n29 4.5005
R10131 VSS.n138 VSS.n29 4.5005
R10132 VSS.n251 VSS.n29 4.5005
R10133 VSS.n137 VSS.n29 4.5005
R10134 VSS.n252 VSS.n29 4.5005
R10135 VSS.n136 VSS.n29 4.5005
R10136 VSS.n253 VSS.n29 4.5005
R10137 VSS.n135 VSS.n29 4.5005
R10138 VSS.n254 VSS.n29 4.5005
R10139 VSS.n134 VSS.n29 4.5005
R10140 VSS.n255 VSS.n29 4.5005
R10141 VSS.n133 VSS.n29 4.5005
R10142 VSS.n256 VSS.n29 4.5005
R10143 VSS.n132 VSS.n29 4.5005
R10144 VSS.n4502 VSS.n29 4.5005
R10145 VSS.n4504 VSS.n29 4.5005
R10146 VSS.n193 VSS.n108 4.5005
R10147 VSS.n195 VSS.n108 4.5005
R10148 VSS.n192 VSS.n108 4.5005
R10149 VSS.n196 VSS.n108 4.5005
R10150 VSS.n191 VSS.n108 4.5005
R10151 VSS.n197 VSS.n108 4.5005
R10152 VSS.n190 VSS.n108 4.5005
R10153 VSS.n198 VSS.n108 4.5005
R10154 VSS.n189 VSS.n108 4.5005
R10155 VSS.n199 VSS.n108 4.5005
R10156 VSS.n188 VSS.n108 4.5005
R10157 VSS.n200 VSS.n108 4.5005
R10158 VSS.n187 VSS.n108 4.5005
R10159 VSS.n201 VSS.n108 4.5005
R10160 VSS.n186 VSS.n108 4.5005
R10161 VSS.n202 VSS.n108 4.5005
R10162 VSS.n185 VSS.n108 4.5005
R10163 VSS.n203 VSS.n108 4.5005
R10164 VSS.n184 VSS.n108 4.5005
R10165 VSS.n204 VSS.n108 4.5005
R10166 VSS.n183 VSS.n108 4.5005
R10167 VSS.n205 VSS.n108 4.5005
R10168 VSS.n182 VSS.n108 4.5005
R10169 VSS.n206 VSS.n108 4.5005
R10170 VSS.n181 VSS.n108 4.5005
R10171 VSS.n207 VSS.n108 4.5005
R10172 VSS.n180 VSS.n108 4.5005
R10173 VSS.n208 VSS.n108 4.5005
R10174 VSS.n179 VSS.n108 4.5005
R10175 VSS.n209 VSS.n108 4.5005
R10176 VSS.n178 VSS.n108 4.5005
R10177 VSS.n210 VSS.n108 4.5005
R10178 VSS.n177 VSS.n108 4.5005
R10179 VSS.n211 VSS.n108 4.5005
R10180 VSS.n176 VSS.n108 4.5005
R10181 VSS.n212 VSS.n108 4.5005
R10182 VSS.n175 VSS.n108 4.5005
R10183 VSS.n213 VSS.n108 4.5005
R10184 VSS.n174 VSS.n108 4.5005
R10185 VSS.n214 VSS.n108 4.5005
R10186 VSS.n173 VSS.n108 4.5005
R10187 VSS.n215 VSS.n108 4.5005
R10188 VSS.n172 VSS.n108 4.5005
R10189 VSS.n216 VSS.n108 4.5005
R10190 VSS.n171 VSS.n108 4.5005
R10191 VSS.n217 VSS.n108 4.5005
R10192 VSS.n170 VSS.n108 4.5005
R10193 VSS.n218 VSS.n108 4.5005
R10194 VSS.n169 VSS.n108 4.5005
R10195 VSS.n219 VSS.n108 4.5005
R10196 VSS.n168 VSS.n108 4.5005
R10197 VSS.n220 VSS.n108 4.5005
R10198 VSS.n167 VSS.n108 4.5005
R10199 VSS.n221 VSS.n108 4.5005
R10200 VSS.n166 VSS.n108 4.5005
R10201 VSS.n222 VSS.n108 4.5005
R10202 VSS.n165 VSS.n108 4.5005
R10203 VSS.n223 VSS.n108 4.5005
R10204 VSS.n164 VSS.n108 4.5005
R10205 VSS.n224 VSS.n108 4.5005
R10206 VSS.n163 VSS.n108 4.5005
R10207 VSS.n225 VSS.n108 4.5005
R10208 VSS.n162 VSS.n108 4.5005
R10209 VSS.n226 VSS.n108 4.5005
R10210 VSS.n161 VSS.n108 4.5005
R10211 VSS.n227 VSS.n108 4.5005
R10212 VSS.n160 VSS.n108 4.5005
R10213 VSS.n228 VSS.n108 4.5005
R10214 VSS.n159 VSS.n108 4.5005
R10215 VSS.n229 VSS.n108 4.5005
R10216 VSS.n158 VSS.n108 4.5005
R10217 VSS.n230 VSS.n108 4.5005
R10218 VSS.n157 VSS.n108 4.5005
R10219 VSS.n231 VSS.n108 4.5005
R10220 VSS.n156 VSS.n108 4.5005
R10221 VSS.n232 VSS.n108 4.5005
R10222 VSS.n155 VSS.n108 4.5005
R10223 VSS.n233 VSS.n108 4.5005
R10224 VSS.n154 VSS.n108 4.5005
R10225 VSS.n234 VSS.n108 4.5005
R10226 VSS.n153 VSS.n108 4.5005
R10227 VSS.n235 VSS.n108 4.5005
R10228 VSS.n4506 VSS.n108 4.5005
R10229 VSS.n236 VSS.n108 4.5005
R10230 VSS.n152 VSS.n108 4.5005
R10231 VSS.n237 VSS.n108 4.5005
R10232 VSS.n151 VSS.n108 4.5005
R10233 VSS.n238 VSS.n108 4.5005
R10234 VSS.n150 VSS.n108 4.5005
R10235 VSS.n239 VSS.n108 4.5005
R10236 VSS.n149 VSS.n108 4.5005
R10237 VSS.n240 VSS.n108 4.5005
R10238 VSS.n148 VSS.n108 4.5005
R10239 VSS.n241 VSS.n108 4.5005
R10240 VSS.n147 VSS.n108 4.5005
R10241 VSS.n242 VSS.n108 4.5005
R10242 VSS.n146 VSS.n108 4.5005
R10243 VSS.n243 VSS.n108 4.5005
R10244 VSS.n145 VSS.n108 4.5005
R10245 VSS.n244 VSS.n108 4.5005
R10246 VSS.n144 VSS.n108 4.5005
R10247 VSS.n245 VSS.n108 4.5005
R10248 VSS.n143 VSS.n108 4.5005
R10249 VSS.n246 VSS.n108 4.5005
R10250 VSS.n142 VSS.n108 4.5005
R10251 VSS.n247 VSS.n108 4.5005
R10252 VSS.n141 VSS.n108 4.5005
R10253 VSS.n248 VSS.n108 4.5005
R10254 VSS.n140 VSS.n108 4.5005
R10255 VSS.n249 VSS.n108 4.5005
R10256 VSS.n139 VSS.n108 4.5005
R10257 VSS.n250 VSS.n108 4.5005
R10258 VSS.n138 VSS.n108 4.5005
R10259 VSS.n251 VSS.n108 4.5005
R10260 VSS.n137 VSS.n108 4.5005
R10261 VSS.n252 VSS.n108 4.5005
R10262 VSS.n136 VSS.n108 4.5005
R10263 VSS.n253 VSS.n108 4.5005
R10264 VSS.n135 VSS.n108 4.5005
R10265 VSS.n254 VSS.n108 4.5005
R10266 VSS.n134 VSS.n108 4.5005
R10267 VSS.n255 VSS.n108 4.5005
R10268 VSS.n133 VSS.n108 4.5005
R10269 VSS.n256 VSS.n108 4.5005
R10270 VSS.n132 VSS.n108 4.5005
R10271 VSS.n4502 VSS.n108 4.5005
R10272 VSS.n4504 VSS.n108 4.5005
R10273 VSS.n193 VSS.n28 4.5005
R10274 VSS.n195 VSS.n28 4.5005
R10275 VSS.n192 VSS.n28 4.5005
R10276 VSS.n196 VSS.n28 4.5005
R10277 VSS.n191 VSS.n28 4.5005
R10278 VSS.n197 VSS.n28 4.5005
R10279 VSS.n190 VSS.n28 4.5005
R10280 VSS.n198 VSS.n28 4.5005
R10281 VSS.n189 VSS.n28 4.5005
R10282 VSS.n199 VSS.n28 4.5005
R10283 VSS.n188 VSS.n28 4.5005
R10284 VSS.n200 VSS.n28 4.5005
R10285 VSS.n187 VSS.n28 4.5005
R10286 VSS.n201 VSS.n28 4.5005
R10287 VSS.n186 VSS.n28 4.5005
R10288 VSS.n202 VSS.n28 4.5005
R10289 VSS.n185 VSS.n28 4.5005
R10290 VSS.n203 VSS.n28 4.5005
R10291 VSS.n184 VSS.n28 4.5005
R10292 VSS.n204 VSS.n28 4.5005
R10293 VSS.n183 VSS.n28 4.5005
R10294 VSS.n205 VSS.n28 4.5005
R10295 VSS.n182 VSS.n28 4.5005
R10296 VSS.n206 VSS.n28 4.5005
R10297 VSS.n181 VSS.n28 4.5005
R10298 VSS.n207 VSS.n28 4.5005
R10299 VSS.n180 VSS.n28 4.5005
R10300 VSS.n208 VSS.n28 4.5005
R10301 VSS.n179 VSS.n28 4.5005
R10302 VSS.n209 VSS.n28 4.5005
R10303 VSS.n178 VSS.n28 4.5005
R10304 VSS.n210 VSS.n28 4.5005
R10305 VSS.n177 VSS.n28 4.5005
R10306 VSS.n211 VSS.n28 4.5005
R10307 VSS.n176 VSS.n28 4.5005
R10308 VSS.n212 VSS.n28 4.5005
R10309 VSS.n175 VSS.n28 4.5005
R10310 VSS.n213 VSS.n28 4.5005
R10311 VSS.n174 VSS.n28 4.5005
R10312 VSS.n214 VSS.n28 4.5005
R10313 VSS.n173 VSS.n28 4.5005
R10314 VSS.n215 VSS.n28 4.5005
R10315 VSS.n172 VSS.n28 4.5005
R10316 VSS.n216 VSS.n28 4.5005
R10317 VSS.n171 VSS.n28 4.5005
R10318 VSS.n217 VSS.n28 4.5005
R10319 VSS.n170 VSS.n28 4.5005
R10320 VSS.n218 VSS.n28 4.5005
R10321 VSS.n169 VSS.n28 4.5005
R10322 VSS.n219 VSS.n28 4.5005
R10323 VSS.n168 VSS.n28 4.5005
R10324 VSS.n220 VSS.n28 4.5005
R10325 VSS.n167 VSS.n28 4.5005
R10326 VSS.n221 VSS.n28 4.5005
R10327 VSS.n166 VSS.n28 4.5005
R10328 VSS.n222 VSS.n28 4.5005
R10329 VSS.n165 VSS.n28 4.5005
R10330 VSS.n223 VSS.n28 4.5005
R10331 VSS.n164 VSS.n28 4.5005
R10332 VSS.n224 VSS.n28 4.5005
R10333 VSS.n163 VSS.n28 4.5005
R10334 VSS.n225 VSS.n28 4.5005
R10335 VSS.n162 VSS.n28 4.5005
R10336 VSS.n226 VSS.n28 4.5005
R10337 VSS.n161 VSS.n28 4.5005
R10338 VSS.n227 VSS.n28 4.5005
R10339 VSS.n160 VSS.n28 4.5005
R10340 VSS.n228 VSS.n28 4.5005
R10341 VSS.n159 VSS.n28 4.5005
R10342 VSS.n229 VSS.n28 4.5005
R10343 VSS.n158 VSS.n28 4.5005
R10344 VSS.n230 VSS.n28 4.5005
R10345 VSS.n157 VSS.n28 4.5005
R10346 VSS.n231 VSS.n28 4.5005
R10347 VSS.n156 VSS.n28 4.5005
R10348 VSS.n232 VSS.n28 4.5005
R10349 VSS.n155 VSS.n28 4.5005
R10350 VSS.n233 VSS.n28 4.5005
R10351 VSS.n154 VSS.n28 4.5005
R10352 VSS.n234 VSS.n28 4.5005
R10353 VSS.n153 VSS.n28 4.5005
R10354 VSS.n235 VSS.n28 4.5005
R10355 VSS.n4506 VSS.n28 4.5005
R10356 VSS.n236 VSS.n28 4.5005
R10357 VSS.n152 VSS.n28 4.5005
R10358 VSS.n237 VSS.n28 4.5005
R10359 VSS.n151 VSS.n28 4.5005
R10360 VSS.n238 VSS.n28 4.5005
R10361 VSS.n150 VSS.n28 4.5005
R10362 VSS.n239 VSS.n28 4.5005
R10363 VSS.n149 VSS.n28 4.5005
R10364 VSS.n240 VSS.n28 4.5005
R10365 VSS.n148 VSS.n28 4.5005
R10366 VSS.n241 VSS.n28 4.5005
R10367 VSS.n147 VSS.n28 4.5005
R10368 VSS.n242 VSS.n28 4.5005
R10369 VSS.n146 VSS.n28 4.5005
R10370 VSS.n243 VSS.n28 4.5005
R10371 VSS.n145 VSS.n28 4.5005
R10372 VSS.n244 VSS.n28 4.5005
R10373 VSS.n144 VSS.n28 4.5005
R10374 VSS.n245 VSS.n28 4.5005
R10375 VSS.n143 VSS.n28 4.5005
R10376 VSS.n246 VSS.n28 4.5005
R10377 VSS.n142 VSS.n28 4.5005
R10378 VSS.n247 VSS.n28 4.5005
R10379 VSS.n141 VSS.n28 4.5005
R10380 VSS.n248 VSS.n28 4.5005
R10381 VSS.n140 VSS.n28 4.5005
R10382 VSS.n249 VSS.n28 4.5005
R10383 VSS.n139 VSS.n28 4.5005
R10384 VSS.n250 VSS.n28 4.5005
R10385 VSS.n138 VSS.n28 4.5005
R10386 VSS.n251 VSS.n28 4.5005
R10387 VSS.n137 VSS.n28 4.5005
R10388 VSS.n252 VSS.n28 4.5005
R10389 VSS.n136 VSS.n28 4.5005
R10390 VSS.n253 VSS.n28 4.5005
R10391 VSS.n135 VSS.n28 4.5005
R10392 VSS.n254 VSS.n28 4.5005
R10393 VSS.n134 VSS.n28 4.5005
R10394 VSS.n255 VSS.n28 4.5005
R10395 VSS.n133 VSS.n28 4.5005
R10396 VSS.n256 VSS.n28 4.5005
R10397 VSS.n132 VSS.n28 4.5005
R10398 VSS.n4502 VSS.n28 4.5005
R10399 VSS.n4504 VSS.n28 4.5005
R10400 VSS.n193 VSS.n109 4.5005
R10401 VSS.n195 VSS.n109 4.5005
R10402 VSS.n192 VSS.n109 4.5005
R10403 VSS.n196 VSS.n109 4.5005
R10404 VSS.n191 VSS.n109 4.5005
R10405 VSS.n197 VSS.n109 4.5005
R10406 VSS.n190 VSS.n109 4.5005
R10407 VSS.n198 VSS.n109 4.5005
R10408 VSS.n189 VSS.n109 4.5005
R10409 VSS.n199 VSS.n109 4.5005
R10410 VSS.n188 VSS.n109 4.5005
R10411 VSS.n200 VSS.n109 4.5005
R10412 VSS.n187 VSS.n109 4.5005
R10413 VSS.n201 VSS.n109 4.5005
R10414 VSS.n186 VSS.n109 4.5005
R10415 VSS.n202 VSS.n109 4.5005
R10416 VSS.n185 VSS.n109 4.5005
R10417 VSS.n203 VSS.n109 4.5005
R10418 VSS.n184 VSS.n109 4.5005
R10419 VSS.n204 VSS.n109 4.5005
R10420 VSS.n183 VSS.n109 4.5005
R10421 VSS.n205 VSS.n109 4.5005
R10422 VSS.n182 VSS.n109 4.5005
R10423 VSS.n206 VSS.n109 4.5005
R10424 VSS.n181 VSS.n109 4.5005
R10425 VSS.n207 VSS.n109 4.5005
R10426 VSS.n180 VSS.n109 4.5005
R10427 VSS.n208 VSS.n109 4.5005
R10428 VSS.n179 VSS.n109 4.5005
R10429 VSS.n209 VSS.n109 4.5005
R10430 VSS.n178 VSS.n109 4.5005
R10431 VSS.n210 VSS.n109 4.5005
R10432 VSS.n177 VSS.n109 4.5005
R10433 VSS.n211 VSS.n109 4.5005
R10434 VSS.n176 VSS.n109 4.5005
R10435 VSS.n212 VSS.n109 4.5005
R10436 VSS.n175 VSS.n109 4.5005
R10437 VSS.n213 VSS.n109 4.5005
R10438 VSS.n174 VSS.n109 4.5005
R10439 VSS.n214 VSS.n109 4.5005
R10440 VSS.n173 VSS.n109 4.5005
R10441 VSS.n215 VSS.n109 4.5005
R10442 VSS.n172 VSS.n109 4.5005
R10443 VSS.n216 VSS.n109 4.5005
R10444 VSS.n171 VSS.n109 4.5005
R10445 VSS.n217 VSS.n109 4.5005
R10446 VSS.n170 VSS.n109 4.5005
R10447 VSS.n218 VSS.n109 4.5005
R10448 VSS.n169 VSS.n109 4.5005
R10449 VSS.n219 VSS.n109 4.5005
R10450 VSS.n168 VSS.n109 4.5005
R10451 VSS.n220 VSS.n109 4.5005
R10452 VSS.n167 VSS.n109 4.5005
R10453 VSS.n221 VSS.n109 4.5005
R10454 VSS.n166 VSS.n109 4.5005
R10455 VSS.n222 VSS.n109 4.5005
R10456 VSS.n165 VSS.n109 4.5005
R10457 VSS.n223 VSS.n109 4.5005
R10458 VSS.n164 VSS.n109 4.5005
R10459 VSS.n224 VSS.n109 4.5005
R10460 VSS.n163 VSS.n109 4.5005
R10461 VSS.n225 VSS.n109 4.5005
R10462 VSS.n162 VSS.n109 4.5005
R10463 VSS.n226 VSS.n109 4.5005
R10464 VSS.n161 VSS.n109 4.5005
R10465 VSS.n227 VSS.n109 4.5005
R10466 VSS.n160 VSS.n109 4.5005
R10467 VSS.n228 VSS.n109 4.5005
R10468 VSS.n159 VSS.n109 4.5005
R10469 VSS.n229 VSS.n109 4.5005
R10470 VSS.n158 VSS.n109 4.5005
R10471 VSS.n230 VSS.n109 4.5005
R10472 VSS.n157 VSS.n109 4.5005
R10473 VSS.n231 VSS.n109 4.5005
R10474 VSS.n156 VSS.n109 4.5005
R10475 VSS.n232 VSS.n109 4.5005
R10476 VSS.n155 VSS.n109 4.5005
R10477 VSS.n233 VSS.n109 4.5005
R10478 VSS.n154 VSS.n109 4.5005
R10479 VSS.n234 VSS.n109 4.5005
R10480 VSS.n153 VSS.n109 4.5005
R10481 VSS.n235 VSS.n109 4.5005
R10482 VSS.n4506 VSS.n109 4.5005
R10483 VSS.n236 VSS.n109 4.5005
R10484 VSS.n152 VSS.n109 4.5005
R10485 VSS.n237 VSS.n109 4.5005
R10486 VSS.n151 VSS.n109 4.5005
R10487 VSS.n238 VSS.n109 4.5005
R10488 VSS.n150 VSS.n109 4.5005
R10489 VSS.n239 VSS.n109 4.5005
R10490 VSS.n149 VSS.n109 4.5005
R10491 VSS.n240 VSS.n109 4.5005
R10492 VSS.n148 VSS.n109 4.5005
R10493 VSS.n241 VSS.n109 4.5005
R10494 VSS.n147 VSS.n109 4.5005
R10495 VSS.n242 VSS.n109 4.5005
R10496 VSS.n146 VSS.n109 4.5005
R10497 VSS.n243 VSS.n109 4.5005
R10498 VSS.n145 VSS.n109 4.5005
R10499 VSS.n244 VSS.n109 4.5005
R10500 VSS.n144 VSS.n109 4.5005
R10501 VSS.n245 VSS.n109 4.5005
R10502 VSS.n143 VSS.n109 4.5005
R10503 VSS.n246 VSS.n109 4.5005
R10504 VSS.n142 VSS.n109 4.5005
R10505 VSS.n247 VSS.n109 4.5005
R10506 VSS.n141 VSS.n109 4.5005
R10507 VSS.n248 VSS.n109 4.5005
R10508 VSS.n140 VSS.n109 4.5005
R10509 VSS.n249 VSS.n109 4.5005
R10510 VSS.n139 VSS.n109 4.5005
R10511 VSS.n250 VSS.n109 4.5005
R10512 VSS.n138 VSS.n109 4.5005
R10513 VSS.n251 VSS.n109 4.5005
R10514 VSS.n137 VSS.n109 4.5005
R10515 VSS.n252 VSS.n109 4.5005
R10516 VSS.n136 VSS.n109 4.5005
R10517 VSS.n253 VSS.n109 4.5005
R10518 VSS.n135 VSS.n109 4.5005
R10519 VSS.n254 VSS.n109 4.5005
R10520 VSS.n134 VSS.n109 4.5005
R10521 VSS.n255 VSS.n109 4.5005
R10522 VSS.n133 VSS.n109 4.5005
R10523 VSS.n256 VSS.n109 4.5005
R10524 VSS.n132 VSS.n109 4.5005
R10525 VSS.n4502 VSS.n109 4.5005
R10526 VSS.n4504 VSS.n109 4.5005
R10527 VSS.n193 VSS.n27 4.5005
R10528 VSS.n195 VSS.n27 4.5005
R10529 VSS.n192 VSS.n27 4.5005
R10530 VSS.n196 VSS.n27 4.5005
R10531 VSS.n191 VSS.n27 4.5005
R10532 VSS.n197 VSS.n27 4.5005
R10533 VSS.n190 VSS.n27 4.5005
R10534 VSS.n198 VSS.n27 4.5005
R10535 VSS.n189 VSS.n27 4.5005
R10536 VSS.n199 VSS.n27 4.5005
R10537 VSS.n188 VSS.n27 4.5005
R10538 VSS.n200 VSS.n27 4.5005
R10539 VSS.n187 VSS.n27 4.5005
R10540 VSS.n201 VSS.n27 4.5005
R10541 VSS.n186 VSS.n27 4.5005
R10542 VSS.n202 VSS.n27 4.5005
R10543 VSS.n185 VSS.n27 4.5005
R10544 VSS.n203 VSS.n27 4.5005
R10545 VSS.n184 VSS.n27 4.5005
R10546 VSS.n204 VSS.n27 4.5005
R10547 VSS.n183 VSS.n27 4.5005
R10548 VSS.n205 VSS.n27 4.5005
R10549 VSS.n182 VSS.n27 4.5005
R10550 VSS.n206 VSS.n27 4.5005
R10551 VSS.n181 VSS.n27 4.5005
R10552 VSS.n207 VSS.n27 4.5005
R10553 VSS.n180 VSS.n27 4.5005
R10554 VSS.n208 VSS.n27 4.5005
R10555 VSS.n179 VSS.n27 4.5005
R10556 VSS.n209 VSS.n27 4.5005
R10557 VSS.n178 VSS.n27 4.5005
R10558 VSS.n210 VSS.n27 4.5005
R10559 VSS.n177 VSS.n27 4.5005
R10560 VSS.n211 VSS.n27 4.5005
R10561 VSS.n176 VSS.n27 4.5005
R10562 VSS.n212 VSS.n27 4.5005
R10563 VSS.n175 VSS.n27 4.5005
R10564 VSS.n213 VSS.n27 4.5005
R10565 VSS.n174 VSS.n27 4.5005
R10566 VSS.n214 VSS.n27 4.5005
R10567 VSS.n173 VSS.n27 4.5005
R10568 VSS.n215 VSS.n27 4.5005
R10569 VSS.n172 VSS.n27 4.5005
R10570 VSS.n216 VSS.n27 4.5005
R10571 VSS.n171 VSS.n27 4.5005
R10572 VSS.n217 VSS.n27 4.5005
R10573 VSS.n170 VSS.n27 4.5005
R10574 VSS.n218 VSS.n27 4.5005
R10575 VSS.n169 VSS.n27 4.5005
R10576 VSS.n219 VSS.n27 4.5005
R10577 VSS.n168 VSS.n27 4.5005
R10578 VSS.n220 VSS.n27 4.5005
R10579 VSS.n167 VSS.n27 4.5005
R10580 VSS.n221 VSS.n27 4.5005
R10581 VSS.n166 VSS.n27 4.5005
R10582 VSS.n222 VSS.n27 4.5005
R10583 VSS.n165 VSS.n27 4.5005
R10584 VSS.n223 VSS.n27 4.5005
R10585 VSS.n164 VSS.n27 4.5005
R10586 VSS.n224 VSS.n27 4.5005
R10587 VSS.n163 VSS.n27 4.5005
R10588 VSS.n225 VSS.n27 4.5005
R10589 VSS.n162 VSS.n27 4.5005
R10590 VSS.n226 VSS.n27 4.5005
R10591 VSS.n161 VSS.n27 4.5005
R10592 VSS.n227 VSS.n27 4.5005
R10593 VSS.n160 VSS.n27 4.5005
R10594 VSS.n228 VSS.n27 4.5005
R10595 VSS.n159 VSS.n27 4.5005
R10596 VSS.n229 VSS.n27 4.5005
R10597 VSS.n158 VSS.n27 4.5005
R10598 VSS.n230 VSS.n27 4.5005
R10599 VSS.n157 VSS.n27 4.5005
R10600 VSS.n231 VSS.n27 4.5005
R10601 VSS.n156 VSS.n27 4.5005
R10602 VSS.n232 VSS.n27 4.5005
R10603 VSS.n155 VSS.n27 4.5005
R10604 VSS.n233 VSS.n27 4.5005
R10605 VSS.n154 VSS.n27 4.5005
R10606 VSS.n234 VSS.n27 4.5005
R10607 VSS.n153 VSS.n27 4.5005
R10608 VSS.n235 VSS.n27 4.5005
R10609 VSS.n4506 VSS.n27 4.5005
R10610 VSS.n236 VSS.n27 4.5005
R10611 VSS.n152 VSS.n27 4.5005
R10612 VSS.n237 VSS.n27 4.5005
R10613 VSS.n151 VSS.n27 4.5005
R10614 VSS.n238 VSS.n27 4.5005
R10615 VSS.n150 VSS.n27 4.5005
R10616 VSS.n239 VSS.n27 4.5005
R10617 VSS.n149 VSS.n27 4.5005
R10618 VSS.n240 VSS.n27 4.5005
R10619 VSS.n148 VSS.n27 4.5005
R10620 VSS.n241 VSS.n27 4.5005
R10621 VSS.n147 VSS.n27 4.5005
R10622 VSS.n242 VSS.n27 4.5005
R10623 VSS.n146 VSS.n27 4.5005
R10624 VSS.n243 VSS.n27 4.5005
R10625 VSS.n145 VSS.n27 4.5005
R10626 VSS.n244 VSS.n27 4.5005
R10627 VSS.n144 VSS.n27 4.5005
R10628 VSS.n245 VSS.n27 4.5005
R10629 VSS.n143 VSS.n27 4.5005
R10630 VSS.n246 VSS.n27 4.5005
R10631 VSS.n142 VSS.n27 4.5005
R10632 VSS.n247 VSS.n27 4.5005
R10633 VSS.n141 VSS.n27 4.5005
R10634 VSS.n248 VSS.n27 4.5005
R10635 VSS.n140 VSS.n27 4.5005
R10636 VSS.n249 VSS.n27 4.5005
R10637 VSS.n139 VSS.n27 4.5005
R10638 VSS.n250 VSS.n27 4.5005
R10639 VSS.n138 VSS.n27 4.5005
R10640 VSS.n251 VSS.n27 4.5005
R10641 VSS.n137 VSS.n27 4.5005
R10642 VSS.n252 VSS.n27 4.5005
R10643 VSS.n136 VSS.n27 4.5005
R10644 VSS.n253 VSS.n27 4.5005
R10645 VSS.n135 VSS.n27 4.5005
R10646 VSS.n254 VSS.n27 4.5005
R10647 VSS.n134 VSS.n27 4.5005
R10648 VSS.n255 VSS.n27 4.5005
R10649 VSS.n133 VSS.n27 4.5005
R10650 VSS.n256 VSS.n27 4.5005
R10651 VSS.n132 VSS.n27 4.5005
R10652 VSS.n4502 VSS.n27 4.5005
R10653 VSS.n4504 VSS.n27 4.5005
R10654 VSS.n193 VSS.n110 4.5005
R10655 VSS.n195 VSS.n110 4.5005
R10656 VSS.n192 VSS.n110 4.5005
R10657 VSS.n196 VSS.n110 4.5005
R10658 VSS.n191 VSS.n110 4.5005
R10659 VSS.n197 VSS.n110 4.5005
R10660 VSS.n190 VSS.n110 4.5005
R10661 VSS.n198 VSS.n110 4.5005
R10662 VSS.n189 VSS.n110 4.5005
R10663 VSS.n199 VSS.n110 4.5005
R10664 VSS.n188 VSS.n110 4.5005
R10665 VSS.n200 VSS.n110 4.5005
R10666 VSS.n187 VSS.n110 4.5005
R10667 VSS.n201 VSS.n110 4.5005
R10668 VSS.n186 VSS.n110 4.5005
R10669 VSS.n202 VSS.n110 4.5005
R10670 VSS.n185 VSS.n110 4.5005
R10671 VSS.n203 VSS.n110 4.5005
R10672 VSS.n184 VSS.n110 4.5005
R10673 VSS.n204 VSS.n110 4.5005
R10674 VSS.n183 VSS.n110 4.5005
R10675 VSS.n205 VSS.n110 4.5005
R10676 VSS.n182 VSS.n110 4.5005
R10677 VSS.n206 VSS.n110 4.5005
R10678 VSS.n181 VSS.n110 4.5005
R10679 VSS.n207 VSS.n110 4.5005
R10680 VSS.n180 VSS.n110 4.5005
R10681 VSS.n208 VSS.n110 4.5005
R10682 VSS.n179 VSS.n110 4.5005
R10683 VSS.n209 VSS.n110 4.5005
R10684 VSS.n178 VSS.n110 4.5005
R10685 VSS.n210 VSS.n110 4.5005
R10686 VSS.n177 VSS.n110 4.5005
R10687 VSS.n211 VSS.n110 4.5005
R10688 VSS.n176 VSS.n110 4.5005
R10689 VSS.n212 VSS.n110 4.5005
R10690 VSS.n175 VSS.n110 4.5005
R10691 VSS.n213 VSS.n110 4.5005
R10692 VSS.n174 VSS.n110 4.5005
R10693 VSS.n214 VSS.n110 4.5005
R10694 VSS.n173 VSS.n110 4.5005
R10695 VSS.n215 VSS.n110 4.5005
R10696 VSS.n172 VSS.n110 4.5005
R10697 VSS.n216 VSS.n110 4.5005
R10698 VSS.n171 VSS.n110 4.5005
R10699 VSS.n217 VSS.n110 4.5005
R10700 VSS.n170 VSS.n110 4.5005
R10701 VSS.n218 VSS.n110 4.5005
R10702 VSS.n169 VSS.n110 4.5005
R10703 VSS.n219 VSS.n110 4.5005
R10704 VSS.n168 VSS.n110 4.5005
R10705 VSS.n220 VSS.n110 4.5005
R10706 VSS.n167 VSS.n110 4.5005
R10707 VSS.n221 VSS.n110 4.5005
R10708 VSS.n166 VSS.n110 4.5005
R10709 VSS.n222 VSS.n110 4.5005
R10710 VSS.n165 VSS.n110 4.5005
R10711 VSS.n223 VSS.n110 4.5005
R10712 VSS.n164 VSS.n110 4.5005
R10713 VSS.n224 VSS.n110 4.5005
R10714 VSS.n163 VSS.n110 4.5005
R10715 VSS.n225 VSS.n110 4.5005
R10716 VSS.n162 VSS.n110 4.5005
R10717 VSS.n226 VSS.n110 4.5005
R10718 VSS.n161 VSS.n110 4.5005
R10719 VSS.n227 VSS.n110 4.5005
R10720 VSS.n160 VSS.n110 4.5005
R10721 VSS.n228 VSS.n110 4.5005
R10722 VSS.n159 VSS.n110 4.5005
R10723 VSS.n229 VSS.n110 4.5005
R10724 VSS.n158 VSS.n110 4.5005
R10725 VSS.n230 VSS.n110 4.5005
R10726 VSS.n157 VSS.n110 4.5005
R10727 VSS.n231 VSS.n110 4.5005
R10728 VSS.n156 VSS.n110 4.5005
R10729 VSS.n232 VSS.n110 4.5005
R10730 VSS.n155 VSS.n110 4.5005
R10731 VSS.n233 VSS.n110 4.5005
R10732 VSS.n154 VSS.n110 4.5005
R10733 VSS.n234 VSS.n110 4.5005
R10734 VSS.n153 VSS.n110 4.5005
R10735 VSS.n235 VSS.n110 4.5005
R10736 VSS.n4506 VSS.n110 4.5005
R10737 VSS.n236 VSS.n110 4.5005
R10738 VSS.n152 VSS.n110 4.5005
R10739 VSS.n237 VSS.n110 4.5005
R10740 VSS.n151 VSS.n110 4.5005
R10741 VSS.n238 VSS.n110 4.5005
R10742 VSS.n150 VSS.n110 4.5005
R10743 VSS.n239 VSS.n110 4.5005
R10744 VSS.n149 VSS.n110 4.5005
R10745 VSS.n240 VSS.n110 4.5005
R10746 VSS.n148 VSS.n110 4.5005
R10747 VSS.n241 VSS.n110 4.5005
R10748 VSS.n147 VSS.n110 4.5005
R10749 VSS.n242 VSS.n110 4.5005
R10750 VSS.n146 VSS.n110 4.5005
R10751 VSS.n243 VSS.n110 4.5005
R10752 VSS.n145 VSS.n110 4.5005
R10753 VSS.n244 VSS.n110 4.5005
R10754 VSS.n144 VSS.n110 4.5005
R10755 VSS.n245 VSS.n110 4.5005
R10756 VSS.n143 VSS.n110 4.5005
R10757 VSS.n246 VSS.n110 4.5005
R10758 VSS.n142 VSS.n110 4.5005
R10759 VSS.n247 VSS.n110 4.5005
R10760 VSS.n141 VSS.n110 4.5005
R10761 VSS.n248 VSS.n110 4.5005
R10762 VSS.n140 VSS.n110 4.5005
R10763 VSS.n249 VSS.n110 4.5005
R10764 VSS.n139 VSS.n110 4.5005
R10765 VSS.n250 VSS.n110 4.5005
R10766 VSS.n138 VSS.n110 4.5005
R10767 VSS.n251 VSS.n110 4.5005
R10768 VSS.n137 VSS.n110 4.5005
R10769 VSS.n252 VSS.n110 4.5005
R10770 VSS.n136 VSS.n110 4.5005
R10771 VSS.n253 VSS.n110 4.5005
R10772 VSS.n135 VSS.n110 4.5005
R10773 VSS.n254 VSS.n110 4.5005
R10774 VSS.n134 VSS.n110 4.5005
R10775 VSS.n255 VSS.n110 4.5005
R10776 VSS.n133 VSS.n110 4.5005
R10777 VSS.n256 VSS.n110 4.5005
R10778 VSS.n132 VSS.n110 4.5005
R10779 VSS.n4502 VSS.n110 4.5005
R10780 VSS.n4504 VSS.n110 4.5005
R10781 VSS.n193 VSS.n26 4.5005
R10782 VSS.n195 VSS.n26 4.5005
R10783 VSS.n192 VSS.n26 4.5005
R10784 VSS.n196 VSS.n26 4.5005
R10785 VSS.n191 VSS.n26 4.5005
R10786 VSS.n197 VSS.n26 4.5005
R10787 VSS.n190 VSS.n26 4.5005
R10788 VSS.n198 VSS.n26 4.5005
R10789 VSS.n189 VSS.n26 4.5005
R10790 VSS.n199 VSS.n26 4.5005
R10791 VSS.n188 VSS.n26 4.5005
R10792 VSS.n200 VSS.n26 4.5005
R10793 VSS.n187 VSS.n26 4.5005
R10794 VSS.n201 VSS.n26 4.5005
R10795 VSS.n186 VSS.n26 4.5005
R10796 VSS.n202 VSS.n26 4.5005
R10797 VSS.n185 VSS.n26 4.5005
R10798 VSS.n203 VSS.n26 4.5005
R10799 VSS.n184 VSS.n26 4.5005
R10800 VSS.n204 VSS.n26 4.5005
R10801 VSS.n183 VSS.n26 4.5005
R10802 VSS.n205 VSS.n26 4.5005
R10803 VSS.n182 VSS.n26 4.5005
R10804 VSS.n206 VSS.n26 4.5005
R10805 VSS.n181 VSS.n26 4.5005
R10806 VSS.n207 VSS.n26 4.5005
R10807 VSS.n180 VSS.n26 4.5005
R10808 VSS.n208 VSS.n26 4.5005
R10809 VSS.n179 VSS.n26 4.5005
R10810 VSS.n209 VSS.n26 4.5005
R10811 VSS.n178 VSS.n26 4.5005
R10812 VSS.n210 VSS.n26 4.5005
R10813 VSS.n177 VSS.n26 4.5005
R10814 VSS.n211 VSS.n26 4.5005
R10815 VSS.n176 VSS.n26 4.5005
R10816 VSS.n212 VSS.n26 4.5005
R10817 VSS.n175 VSS.n26 4.5005
R10818 VSS.n213 VSS.n26 4.5005
R10819 VSS.n174 VSS.n26 4.5005
R10820 VSS.n214 VSS.n26 4.5005
R10821 VSS.n173 VSS.n26 4.5005
R10822 VSS.n215 VSS.n26 4.5005
R10823 VSS.n172 VSS.n26 4.5005
R10824 VSS.n216 VSS.n26 4.5005
R10825 VSS.n171 VSS.n26 4.5005
R10826 VSS.n217 VSS.n26 4.5005
R10827 VSS.n170 VSS.n26 4.5005
R10828 VSS.n218 VSS.n26 4.5005
R10829 VSS.n169 VSS.n26 4.5005
R10830 VSS.n219 VSS.n26 4.5005
R10831 VSS.n168 VSS.n26 4.5005
R10832 VSS.n220 VSS.n26 4.5005
R10833 VSS.n167 VSS.n26 4.5005
R10834 VSS.n221 VSS.n26 4.5005
R10835 VSS.n166 VSS.n26 4.5005
R10836 VSS.n222 VSS.n26 4.5005
R10837 VSS.n165 VSS.n26 4.5005
R10838 VSS.n223 VSS.n26 4.5005
R10839 VSS.n164 VSS.n26 4.5005
R10840 VSS.n224 VSS.n26 4.5005
R10841 VSS.n163 VSS.n26 4.5005
R10842 VSS.n225 VSS.n26 4.5005
R10843 VSS.n162 VSS.n26 4.5005
R10844 VSS.n226 VSS.n26 4.5005
R10845 VSS.n161 VSS.n26 4.5005
R10846 VSS.n227 VSS.n26 4.5005
R10847 VSS.n160 VSS.n26 4.5005
R10848 VSS.n228 VSS.n26 4.5005
R10849 VSS.n159 VSS.n26 4.5005
R10850 VSS.n229 VSS.n26 4.5005
R10851 VSS.n158 VSS.n26 4.5005
R10852 VSS.n230 VSS.n26 4.5005
R10853 VSS.n157 VSS.n26 4.5005
R10854 VSS.n231 VSS.n26 4.5005
R10855 VSS.n156 VSS.n26 4.5005
R10856 VSS.n232 VSS.n26 4.5005
R10857 VSS.n155 VSS.n26 4.5005
R10858 VSS.n233 VSS.n26 4.5005
R10859 VSS.n154 VSS.n26 4.5005
R10860 VSS.n234 VSS.n26 4.5005
R10861 VSS.n153 VSS.n26 4.5005
R10862 VSS.n235 VSS.n26 4.5005
R10863 VSS.n4506 VSS.n26 4.5005
R10864 VSS.n236 VSS.n26 4.5005
R10865 VSS.n152 VSS.n26 4.5005
R10866 VSS.n237 VSS.n26 4.5005
R10867 VSS.n151 VSS.n26 4.5005
R10868 VSS.n238 VSS.n26 4.5005
R10869 VSS.n150 VSS.n26 4.5005
R10870 VSS.n239 VSS.n26 4.5005
R10871 VSS.n149 VSS.n26 4.5005
R10872 VSS.n240 VSS.n26 4.5005
R10873 VSS.n148 VSS.n26 4.5005
R10874 VSS.n241 VSS.n26 4.5005
R10875 VSS.n147 VSS.n26 4.5005
R10876 VSS.n242 VSS.n26 4.5005
R10877 VSS.n146 VSS.n26 4.5005
R10878 VSS.n243 VSS.n26 4.5005
R10879 VSS.n145 VSS.n26 4.5005
R10880 VSS.n244 VSS.n26 4.5005
R10881 VSS.n144 VSS.n26 4.5005
R10882 VSS.n245 VSS.n26 4.5005
R10883 VSS.n143 VSS.n26 4.5005
R10884 VSS.n246 VSS.n26 4.5005
R10885 VSS.n142 VSS.n26 4.5005
R10886 VSS.n247 VSS.n26 4.5005
R10887 VSS.n141 VSS.n26 4.5005
R10888 VSS.n248 VSS.n26 4.5005
R10889 VSS.n140 VSS.n26 4.5005
R10890 VSS.n249 VSS.n26 4.5005
R10891 VSS.n139 VSS.n26 4.5005
R10892 VSS.n250 VSS.n26 4.5005
R10893 VSS.n138 VSS.n26 4.5005
R10894 VSS.n251 VSS.n26 4.5005
R10895 VSS.n137 VSS.n26 4.5005
R10896 VSS.n252 VSS.n26 4.5005
R10897 VSS.n136 VSS.n26 4.5005
R10898 VSS.n253 VSS.n26 4.5005
R10899 VSS.n135 VSS.n26 4.5005
R10900 VSS.n254 VSS.n26 4.5005
R10901 VSS.n134 VSS.n26 4.5005
R10902 VSS.n255 VSS.n26 4.5005
R10903 VSS.n133 VSS.n26 4.5005
R10904 VSS.n256 VSS.n26 4.5005
R10905 VSS.n132 VSS.n26 4.5005
R10906 VSS.n4502 VSS.n26 4.5005
R10907 VSS.n4504 VSS.n26 4.5005
R10908 VSS.n193 VSS.n111 4.5005
R10909 VSS.n195 VSS.n111 4.5005
R10910 VSS.n192 VSS.n111 4.5005
R10911 VSS.n196 VSS.n111 4.5005
R10912 VSS.n191 VSS.n111 4.5005
R10913 VSS.n197 VSS.n111 4.5005
R10914 VSS.n190 VSS.n111 4.5005
R10915 VSS.n198 VSS.n111 4.5005
R10916 VSS.n189 VSS.n111 4.5005
R10917 VSS.n199 VSS.n111 4.5005
R10918 VSS.n188 VSS.n111 4.5005
R10919 VSS.n200 VSS.n111 4.5005
R10920 VSS.n187 VSS.n111 4.5005
R10921 VSS.n201 VSS.n111 4.5005
R10922 VSS.n186 VSS.n111 4.5005
R10923 VSS.n202 VSS.n111 4.5005
R10924 VSS.n185 VSS.n111 4.5005
R10925 VSS.n203 VSS.n111 4.5005
R10926 VSS.n184 VSS.n111 4.5005
R10927 VSS.n204 VSS.n111 4.5005
R10928 VSS.n183 VSS.n111 4.5005
R10929 VSS.n205 VSS.n111 4.5005
R10930 VSS.n182 VSS.n111 4.5005
R10931 VSS.n206 VSS.n111 4.5005
R10932 VSS.n181 VSS.n111 4.5005
R10933 VSS.n207 VSS.n111 4.5005
R10934 VSS.n180 VSS.n111 4.5005
R10935 VSS.n208 VSS.n111 4.5005
R10936 VSS.n179 VSS.n111 4.5005
R10937 VSS.n209 VSS.n111 4.5005
R10938 VSS.n178 VSS.n111 4.5005
R10939 VSS.n210 VSS.n111 4.5005
R10940 VSS.n177 VSS.n111 4.5005
R10941 VSS.n211 VSS.n111 4.5005
R10942 VSS.n176 VSS.n111 4.5005
R10943 VSS.n212 VSS.n111 4.5005
R10944 VSS.n175 VSS.n111 4.5005
R10945 VSS.n213 VSS.n111 4.5005
R10946 VSS.n174 VSS.n111 4.5005
R10947 VSS.n214 VSS.n111 4.5005
R10948 VSS.n173 VSS.n111 4.5005
R10949 VSS.n215 VSS.n111 4.5005
R10950 VSS.n172 VSS.n111 4.5005
R10951 VSS.n216 VSS.n111 4.5005
R10952 VSS.n171 VSS.n111 4.5005
R10953 VSS.n217 VSS.n111 4.5005
R10954 VSS.n170 VSS.n111 4.5005
R10955 VSS.n218 VSS.n111 4.5005
R10956 VSS.n169 VSS.n111 4.5005
R10957 VSS.n219 VSS.n111 4.5005
R10958 VSS.n168 VSS.n111 4.5005
R10959 VSS.n220 VSS.n111 4.5005
R10960 VSS.n167 VSS.n111 4.5005
R10961 VSS.n221 VSS.n111 4.5005
R10962 VSS.n166 VSS.n111 4.5005
R10963 VSS.n222 VSS.n111 4.5005
R10964 VSS.n165 VSS.n111 4.5005
R10965 VSS.n223 VSS.n111 4.5005
R10966 VSS.n164 VSS.n111 4.5005
R10967 VSS.n224 VSS.n111 4.5005
R10968 VSS.n163 VSS.n111 4.5005
R10969 VSS.n225 VSS.n111 4.5005
R10970 VSS.n162 VSS.n111 4.5005
R10971 VSS.n226 VSS.n111 4.5005
R10972 VSS.n161 VSS.n111 4.5005
R10973 VSS.n227 VSS.n111 4.5005
R10974 VSS.n160 VSS.n111 4.5005
R10975 VSS.n228 VSS.n111 4.5005
R10976 VSS.n159 VSS.n111 4.5005
R10977 VSS.n229 VSS.n111 4.5005
R10978 VSS.n158 VSS.n111 4.5005
R10979 VSS.n230 VSS.n111 4.5005
R10980 VSS.n157 VSS.n111 4.5005
R10981 VSS.n231 VSS.n111 4.5005
R10982 VSS.n156 VSS.n111 4.5005
R10983 VSS.n232 VSS.n111 4.5005
R10984 VSS.n155 VSS.n111 4.5005
R10985 VSS.n233 VSS.n111 4.5005
R10986 VSS.n154 VSS.n111 4.5005
R10987 VSS.n234 VSS.n111 4.5005
R10988 VSS.n153 VSS.n111 4.5005
R10989 VSS.n235 VSS.n111 4.5005
R10990 VSS.n4506 VSS.n111 4.5005
R10991 VSS.n236 VSS.n111 4.5005
R10992 VSS.n152 VSS.n111 4.5005
R10993 VSS.n237 VSS.n111 4.5005
R10994 VSS.n151 VSS.n111 4.5005
R10995 VSS.n238 VSS.n111 4.5005
R10996 VSS.n150 VSS.n111 4.5005
R10997 VSS.n239 VSS.n111 4.5005
R10998 VSS.n149 VSS.n111 4.5005
R10999 VSS.n240 VSS.n111 4.5005
R11000 VSS.n148 VSS.n111 4.5005
R11001 VSS.n241 VSS.n111 4.5005
R11002 VSS.n147 VSS.n111 4.5005
R11003 VSS.n242 VSS.n111 4.5005
R11004 VSS.n146 VSS.n111 4.5005
R11005 VSS.n243 VSS.n111 4.5005
R11006 VSS.n145 VSS.n111 4.5005
R11007 VSS.n244 VSS.n111 4.5005
R11008 VSS.n144 VSS.n111 4.5005
R11009 VSS.n245 VSS.n111 4.5005
R11010 VSS.n143 VSS.n111 4.5005
R11011 VSS.n246 VSS.n111 4.5005
R11012 VSS.n142 VSS.n111 4.5005
R11013 VSS.n247 VSS.n111 4.5005
R11014 VSS.n141 VSS.n111 4.5005
R11015 VSS.n248 VSS.n111 4.5005
R11016 VSS.n140 VSS.n111 4.5005
R11017 VSS.n249 VSS.n111 4.5005
R11018 VSS.n139 VSS.n111 4.5005
R11019 VSS.n250 VSS.n111 4.5005
R11020 VSS.n138 VSS.n111 4.5005
R11021 VSS.n251 VSS.n111 4.5005
R11022 VSS.n137 VSS.n111 4.5005
R11023 VSS.n252 VSS.n111 4.5005
R11024 VSS.n136 VSS.n111 4.5005
R11025 VSS.n253 VSS.n111 4.5005
R11026 VSS.n135 VSS.n111 4.5005
R11027 VSS.n254 VSS.n111 4.5005
R11028 VSS.n134 VSS.n111 4.5005
R11029 VSS.n255 VSS.n111 4.5005
R11030 VSS.n133 VSS.n111 4.5005
R11031 VSS.n256 VSS.n111 4.5005
R11032 VSS.n132 VSS.n111 4.5005
R11033 VSS.n4502 VSS.n111 4.5005
R11034 VSS.n4504 VSS.n111 4.5005
R11035 VSS.n193 VSS.n25 4.5005
R11036 VSS.n195 VSS.n25 4.5005
R11037 VSS.n192 VSS.n25 4.5005
R11038 VSS.n196 VSS.n25 4.5005
R11039 VSS.n191 VSS.n25 4.5005
R11040 VSS.n197 VSS.n25 4.5005
R11041 VSS.n190 VSS.n25 4.5005
R11042 VSS.n198 VSS.n25 4.5005
R11043 VSS.n189 VSS.n25 4.5005
R11044 VSS.n199 VSS.n25 4.5005
R11045 VSS.n188 VSS.n25 4.5005
R11046 VSS.n200 VSS.n25 4.5005
R11047 VSS.n187 VSS.n25 4.5005
R11048 VSS.n201 VSS.n25 4.5005
R11049 VSS.n186 VSS.n25 4.5005
R11050 VSS.n202 VSS.n25 4.5005
R11051 VSS.n185 VSS.n25 4.5005
R11052 VSS.n203 VSS.n25 4.5005
R11053 VSS.n184 VSS.n25 4.5005
R11054 VSS.n204 VSS.n25 4.5005
R11055 VSS.n183 VSS.n25 4.5005
R11056 VSS.n205 VSS.n25 4.5005
R11057 VSS.n182 VSS.n25 4.5005
R11058 VSS.n206 VSS.n25 4.5005
R11059 VSS.n181 VSS.n25 4.5005
R11060 VSS.n207 VSS.n25 4.5005
R11061 VSS.n180 VSS.n25 4.5005
R11062 VSS.n208 VSS.n25 4.5005
R11063 VSS.n179 VSS.n25 4.5005
R11064 VSS.n209 VSS.n25 4.5005
R11065 VSS.n178 VSS.n25 4.5005
R11066 VSS.n210 VSS.n25 4.5005
R11067 VSS.n177 VSS.n25 4.5005
R11068 VSS.n211 VSS.n25 4.5005
R11069 VSS.n176 VSS.n25 4.5005
R11070 VSS.n212 VSS.n25 4.5005
R11071 VSS.n175 VSS.n25 4.5005
R11072 VSS.n213 VSS.n25 4.5005
R11073 VSS.n174 VSS.n25 4.5005
R11074 VSS.n214 VSS.n25 4.5005
R11075 VSS.n173 VSS.n25 4.5005
R11076 VSS.n215 VSS.n25 4.5005
R11077 VSS.n172 VSS.n25 4.5005
R11078 VSS.n216 VSS.n25 4.5005
R11079 VSS.n171 VSS.n25 4.5005
R11080 VSS.n217 VSS.n25 4.5005
R11081 VSS.n170 VSS.n25 4.5005
R11082 VSS.n218 VSS.n25 4.5005
R11083 VSS.n169 VSS.n25 4.5005
R11084 VSS.n219 VSS.n25 4.5005
R11085 VSS.n168 VSS.n25 4.5005
R11086 VSS.n220 VSS.n25 4.5005
R11087 VSS.n167 VSS.n25 4.5005
R11088 VSS.n221 VSS.n25 4.5005
R11089 VSS.n166 VSS.n25 4.5005
R11090 VSS.n222 VSS.n25 4.5005
R11091 VSS.n165 VSS.n25 4.5005
R11092 VSS.n223 VSS.n25 4.5005
R11093 VSS.n164 VSS.n25 4.5005
R11094 VSS.n224 VSS.n25 4.5005
R11095 VSS.n163 VSS.n25 4.5005
R11096 VSS.n225 VSS.n25 4.5005
R11097 VSS.n162 VSS.n25 4.5005
R11098 VSS.n226 VSS.n25 4.5005
R11099 VSS.n161 VSS.n25 4.5005
R11100 VSS.n227 VSS.n25 4.5005
R11101 VSS.n160 VSS.n25 4.5005
R11102 VSS.n228 VSS.n25 4.5005
R11103 VSS.n159 VSS.n25 4.5005
R11104 VSS.n229 VSS.n25 4.5005
R11105 VSS.n158 VSS.n25 4.5005
R11106 VSS.n230 VSS.n25 4.5005
R11107 VSS.n157 VSS.n25 4.5005
R11108 VSS.n231 VSS.n25 4.5005
R11109 VSS.n156 VSS.n25 4.5005
R11110 VSS.n232 VSS.n25 4.5005
R11111 VSS.n155 VSS.n25 4.5005
R11112 VSS.n233 VSS.n25 4.5005
R11113 VSS.n154 VSS.n25 4.5005
R11114 VSS.n234 VSS.n25 4.5005
R11115 VSS.n153 VSS.n25 4.5005
R11116 VSS.n235 VSS.n25 4.5005
R11117 VSS.n4506 VSS.n25 4.5005
R11118 VSS.n236 VSS.n25 4.5005
R11119 VSS.n152 VSS.n25 4.5005
R11120 VSS.n237 VSS.n25 4.5005
R11121 VSS.n151 VSS.n25 4.5005
R11122 VSS.n238 VSS.n25 4.5005
R11123 VSS.n150 VSS.n25 4.5005
R11124 VSS.n239 VSS.n25 4.5005
R11125 VSS.n149 VSS.n25 4.5005
R11126 VSS.n240 VSS.n25 4.5005
R11127 VSS.n148 VSS.n25 4.5005
R11128 VSS.n241 VSS.n25 4.5005
R11129 VSS.n147 VSS.n25 4.5005
R11130 VSS.n242 VSS.n25 4.5005
R11131 VSS.n146 VSS.n25 4.5005
R11132 VSS.n243 VSS.n25 4.5005
R11133 VSS.n145 VSS.n25 4.5005
R11134 VSS.n244 VSS.n25 4.5005
R11135 VSS.n144 VSS.n25 4.5005
R11136 VSS.n245 VSS.n25 4.5005
R11137 VSS.n143 VSS.n25 4.5005
R11138 VSS.n246 VSS.n25 4.5005
R11139 VSS.n142 VSS.n25 4.5005
R11140 VSS.n247 VSS.n25 4.5005
R11141 VSS.n141 VSS.n25 4.5005
R11142 VSS.n248 VSS.n25 4.5005
R11143 VSS.n140 VSS.n25 4.5005
R11144 VSS.n249 VSS.n25 4.5005
R11145 VSS.n139 VSS.n25 4.5005
R11146 VSS.n250 VSS.n25 4.5005
R11147 VSS.n138 VSS.n25 4.5005
R11148 VSS.n251 VSS.n25 4.5005
R11149 VSS.n137 VSS.n25 4.5005
R11150 VSS.n252 VSS.n25 4.5005
R11151 VSS.n136 VSS.n25 4.5005
R11152 VSS.n253 VSS.n25 4.5005
R11153 VSS.n135 VSS.n25 4.5005
R11154 VSS.n254 VSS.n25 4.5005
R11155 VSS.n134 VSS.n25 4.5005
R11156 VSS.n255 VSS.n25 4.5005
R11157 VSS.n133 VSS.n25 4.5005
R11158 VSS.n256 VSS.n25 4.5005
R11159 VSS.n132 VSS.n25 4.5005
R11160 VSS.n4502 VSS.n25 4.5005
R11161 VSS.n4504 VSS.n25 4.5005
R11162 VSS.n193 VSS.n112 4.5005
R11163 VSS.n195 VSS.n112 4.5005
R11164 VSS.n192 VSS.n112 4.5005
R11165 VSS.n196 VSS.n112 4.5005
R11166 VSS.n191 VSS.n112 4.5005
R11167 VSS.n197 VSS.n112 4.5005
R11168 VSS.n190 VSS.n112 4.5005
R11169 VSS.n198 VSS.n112 4.5005
R11170 VSS.n189 VSS.n112 4.5005
R11171 VSS.n199 VSS.n112 4.5005
R11172 VSS.n188 VSS.n112 4.5005
R11173 VSS.n200 VSS.n112 4.5005
R11174 VSS.n187 VSS.n112 4.5005
R11175 VSS.n201 VSS.n112 4.5005
R11176 VSS.n186 VSS.n112 4.5005
R11177 VSS.n202 VSS.n112 4.5005
R11178 VSS.n185 VSS.n112 4.5005
R11179 VSS.n203 VSS.n112 4.5005
R11180 VSS.n184 VSS.n112 4.5005
R11181 VSS.n204 VSS.n112 4.5005
R11182 VSS.n183 VSS.n112 4.5005
R11183 VSS.n205 VSS.n112 4.5005
R11184 VSS.n182 VSS.n112 4.5005
R11185 VSS.n206 VSS.n112 4.5005
R11186 VSS.n181 VSS.n112 4.5005
R11187 VSS.n207 VSS.n112 4.5005
R11188 VSS.n180 VSS.n112 4.5005
R11189 VSS.n208 VSS.n112 4.5005
R11190 VSS.n179 VSS.n112 4.5005
R11191 VSS.n209 VSS.n112 4.5005
R11192 VSS.n178 VSS.n112 4.5005
R11193 VSS.n210 VSS.n112 4.5005
R11194 VSS.n177 VSS.n112 4.5005
R11195 VSS.n211 VSS.n112 4.5005
R11196 VSS.n176 VSS.n112 4.5005
R11197 VSS.n212 VSS.n112 4.5005
R11198 VSS.n175 VSS.n112 4.5005
R11199 VSS.n213 VSS.n112 4.5005
R11200 VSS.n174 VSS.n112 4.5005
R11201 VSS.n214 VSS.n112 4.5005
R11202 VSS.n173 VSS.n112 4.5005
R11203 VSS.n215 VSS.n112 4.5005
R11204 VSS.n172 VSS.n112 4.5005
R11205 VSS.n216 VSS.n112 4.5005
R11206 VSS.n171 VSS.n112 4.5005
R11207 VSS.n217 VSS.n112 4.5005
R11208 VSS.n170 VSS.n112 4.5005
R11209 VSS.n218 VSS.n112 4.5005
R11210 VSS.n169 VSS.n112 4.5005
R11211 VSS.n219 VSS.n112 4.5005
R11212 VSS.n168 VSS.n112 4.5005
R11213 VSS.n220 VSS.n112 4.5005
R11214 VSS.n167 VSS.n112 4.5005
R11215 VSS.n221 VSS.n112 4.5005
R11216 VSS.n166 VSS.n112 4.5005
R11217 VSS.n222 VSS.n112 4.5005
R11218 VSS.n165 VSS.n112 4.5005
R11219 VSS.n223 VSS.n112 4.5005
R11220 VSS.n164 VSS.n112 4.5005
R11221 VSS.n224 VSS.n112 4.5005
R11222 VSS.n163 VSS.n112 4.5005
R11223 VSS.n225 VSS.n112 4.5005
R11224 VSS.n162 VSS.n112 4.5005
R11225 VSS.n226 VSS.n112 4.5005
R11226 VSS.n161 VSS.n112 4.5005
R11227 VSS.n227 VSS.n112 4.5005
R11228 VSS.n160 VSS.n112 4.5005
R11229 VSS.n228 VSS.n112 4.5005
R11230 VSS.n159 VSS.n112 4.5005
R11231 VSS.n229 VSS.n112 4.5005
R11232 VSS.n158 VSS.n112 4.5005
R11233 VSS.n230 VSS.n112 4.5005
R11234 VSS.n157 VSS.n112 4.5005
R11235 VSS.n231 VSS.n112 4.5005
R11236 VSS.n156 VSS.n112 4.5005
R11237 VSS.n232 VSS.n112 4.5005
R11238 VSS.n155 VSS.n112 4.5005
R11239 VSS.n233 VSS.n112 4.5005
R11240 VSS.n154 VSS.n112 4.5005
R11241 VSS.n234 VSS.n112 4.5005
R11242 VSS.n153 VSS.n112 4.5005
R11243 VSS.n235 VSS.n112 4.5005
R11244 VSS.n4506 VSS.n112 4.5005
R11245 VSS.n236 VSS.n112 4.5005
R11246 VSS.n152 VSS.n112 4.5005
R11247 VSS.n237 VSS.n112 4.5005
R11248 VSS.n151 VSS.n112 4.5005
R11249 VSS.n238 VSS.n112 4.5005
R11250 VSS.n150 VSS.n112 4.5005
R11251 VSS.n239 VSS.n112 4.5005
R11252 VSS.n149 VSS.n112 4.5005
R11253 VSS.n240 VSS.n112 4.5005
R11254 VSS.n148 VSS.n112 4.5005
R11255 VSS.n241 VSS.n112 4.5005
R11256 VSS.n147 VSS.n112 4.5005
R11257 VSS.n242 VSS.n112 4.5005
R11258 VSS.n146 VSS.n112 4.5005
R11259 VSS.n243 VSS.n112 4.5005
R11260 VSS.n145 VSS.n112 4.5005
R11261 VSS.n244 VSS.n112 4.5005
R11262 VSS.n144 VSS.n112 4.5005
R11263 VSS.n245 VSS.n112 4.5005
R11264 VSS.n143 VSS.n112 4.5005
R11265 VSS.n246 VSS.n112 4.5005
R11266 VSS.n142 VSS.n112 4.5005
R11267 VSS.n247 VSS.n112 4.5005
R11268 VSS.n141 VSS.n112 4.5005
R11269 VSS.n248 VSS.n112 4.5005
R11270 VSS.n140 VSS.n112 4.5005
R11271 VSS.n249 VSS.n112 4.5005
R11272 VSS.n139 VSS.n112 4.5005
R11273 VSS.n250 VSS.n112 4.5005
R11274 VSS.n138 VSS.n112 4.5005
R11275 VSS.n251 VSS.n112 4.5005
R11276 VSS.n137 VSS.n112 4.5005
R11277 VSS.n252 VSS.n112 4.5005
R11278 VSS.n136 VSS.n112 4.5005
R11279 VSS.n253 VSS.n112 4.5005
R11280 VSS.n135 VSS.n112 4.5005
R11281 VSS.n254 VSS.n112 4.5005
R11282 VSS.n134 VSS.n112 4.5005
R11283 VSS.n255 VSS.n112 4.5005
R11284 VSS.n133 VSS.n112 4.5005
R11285 VSS.n256 VSS.n112 4.5005
R11286 VSS.n132 VSS.n112 4.5005
R11287 VSS.n4502 VSS.n112 4.5005
R11288 VSS.n4504 VSS.n112 4.5005
R11289 VSS.n193 VSS.n24 4.5005
R11290 VSS.n195 VSS.n24 4.5005
R11291 VSS.n192 VSS.n24 4.5005
R11292 VSS.n196 VSS.n24 4.5005
R11293 VSS.n191 VSS.n24 4.5005
R11294 VSS.n197 VSS.n24 4.5005
R11295 VSS.n190 VSS.n24 4.5005
R11296 VSS.n198 VSS.n24 4.5005
R11297 VSS.n189 VSS.n24 4.5005
R11298 VSS.n199 VSS.n24 4.5005
R11299 VSS.n188 VSS.n24 4.5005
R11300 VSS.n200 VSS.n24 4.5005
R11301 VSS.n187 VSS.n24 4.5005
R11302 VSS.n201 VSS.n24 4.5005
R11303 VSS.n186 VSS.n24 4.5005
R11304 VSS.n202 VSS.n24 4.5005
R11305 VSS.n185 VSS.n24 4.5005
R11306 VSS.n203 VSS.n24 4.5005
R11307 VSS.n184 VSS.n24 4.5005
R11308 VSS.n204 VSS.n24 4.5005
R11309 VSS.n183 VSS.n24 4.5005
R11310 VSS.n205 VSS.n24 4.5005
R11311 VSS.n182 VSS.n24 4.5005
R11312 VSS.n206 VSS.n24 4.5005
R11313 VSS.n181 VSS.n24 4.5005
R11314 VSS.n207 VSS.n24 4.5005
R11315 VSS.n180 VSS.n24 4.5005
R11316 VSS.n208 VSS.n24 4.5005
R11317 VSS.n179 VSS.n24 4.5005
R11318 VSS.n209 VSS.n24 4.5005
R11319 VSS.n178 VSS.n24 4.5005
R11320 VSS.n210 VSS.n24 4.5005
R11321 VSS.n177 VSS.n24 4.5005
R11322 VSS.n211 VSS.n24 4.5005
R11323 VSS.n176 VSS.n24 4.5005
R11324 VSS.n212 VSS.n24 4.5005
R11325 VSS.n175 VSS.n24 4.5005
R11326 VSS.n213 VSS.n24 4.5005
R11327 VSS.n174 VSS.n24 4.5005
R11328 VSS.n214 VSS.n24 4.5005
R11329 VSS.n173 VSS.n24 4.5005
R11330 VSS.n215 VSS.n24 4.5005
R11331 VSS.n172 VSS.n24 4.5005
R11332 VSS.n216 VSS.n24 4.5005
R11333 VSS.n171 VSS.n24 4.5005
R11334 VSS.n217 VSS.n24 4.5005
R11335 VSS.n170 VSS.n24 4.5005
R11336 VSS.n218 VSS.n24 4.5005
R11337 VSS.n169 VSS.n24 4.5005
R11338 VSS.n219 VSS.n24 4.5005
R11339 VSS.n168 VSS.n24 4.5005
R11340 VSS.n220 VSS.n24 4.5005
R11341 VSS.n167 VSS.n24 4.5005
R11342 VSS.n221 VSS.n24 4.5005
R11343 VSS.n166 VSS.n24 4.5005
R11344 VSS.n222 VSS.n24 4.5005
R11345 VSS.n165 VSS.n24 4.5005
R11346 VSS.n223 VSS.n24 4.5005
R11347 VSS.n164 VSS.n24 4.5005
R11348 VSS.n224 VSS.n24 4.5005
R11349 VSS.n163 VSS.n24 4.5005
R11350 VSS.n225 VSS.n24 4.5005
R11351 VSS.n162 VSS.n24 4.5005
R11352 VSS.n226 VSS.n24 4.5005
R11353 VSS.n161 VSS.n24 4.5005
R11354 VSS.n227 VSS.n24 4.5005
R11355 VSS.n160 VSS.n24 4.5005
R11356 VSS.n228 VSS.n24 4.5005
R11357 VSS.n159 VSS.n24 4.5005
R11358 VSS.n229 VSS.n24 4.5005
R11359 VSS.n158 VSS.n24 4.5005
R11360 VSS.n230 VSS.n24 4.5005
R11361 VSS.n157 VSS.n24 4.5005
R11362 VSS.n231 VSS.n24 4.5005
R11363 VSS.n156 VSS.n24 4.5005
R11364 VSS.n232 VSS.n24 4.5005
R11365 VSS.n155 VSS.n24 4.5005
R11366 VSS.n233 VSS.n24 4.5005
R11367 VSS.n154 VSS.n24 4.5005
R11368 VSS.n234 VSS.n24 4.5005
R11369 VSS.n153 VSS.n24 4.5005
R11370 VSS.n235 VSS.n24 4.5005
R11371 VSS.n4506 VSS.n24 4.5005
R11372 VSS.n236 VSS.n24 4.5005
R11373 VSS.n152 VSS.n24 4.5005
R11374 VSS.n237 VSS.n24 4.5005
R11375 VSS.n151 VSS.n24 4.5005
R11376 VSS.n238 VSS.n24 4.5005
R11377 VSS.n150 VSS.n24 4.5005
R11378 VSS.n239 VSS.n24 4.5005
R11379 VSS.n149 VSS.n24 4.5005
R11380 VSS.n240 VSS.n24 4.5005
R11381 VSS.n148 VSS.n24 4.5005
R11382 VSS.n241 VSS.n24 4.5005
R11383 VSS.n147 VSS.n24 4.5005
R11384 VSS.n242 VSS.n24 4.5005
R11385 VSS.n146 VSS.n24 4.5005
R11386 VSS.n243 VSS.n24 4.5005
R11387 VSS.n145 VSS.n24 4.5005
R11388 VSS.n244 VSS.n24 4.5005
R11389 VSS.n144 VSS.n24 4.5005
R11390 VSS.n245 VSS.n24 4.5005
R11391 VSS.n143 VSS.n24 4.5005
R11392 VSS.n246 VSS.n24 4.5005
R11393 VSS.n142 VSS.n24 4.5005
R11394 VSS.n247 VSS.n24 4.5005
R11395 VSS.n141 VSS.n24 4.5005
R11396 VSS.n248 VSS.n24 4.5005
R11397 VSS.n140 VSS.n24 4.5005
R11398 VSS.n249 VSS.n24 4.5005
R11399 VSS.n139 VSS.n24 4.5005
R11400 VSS.n250 VSS.n24 4.5005
R11401 VSS.n138 VSS.n24 4.5005
R11402 VSS.n251 VSS.n24 4.5005
R11403 VSS.n137 VSS.n24 4.5005
R11404 VSS.n252 VSS.n24 4.5005
R11405 VSS.n136 VSS.n24 4.5005
R11406 VSS.n253 VSS.n24 4.5005
R11407 VSS.n135 VSS.n24 4.5005
R11408 VSS.n254 VSS.n24 4.5005
R11409 VSS.n134 VSS.n24 4.5005
R11410 VSS.n255 VSS.n24 4.5005
R11411 VSS.n133 VSS.n24 4.5005
R11412 VSS.n256 VSS.n24 4.5005
R11413 VSS.n132 VSS.n24 4.5005
R11414 VSS.n4502 VSS.n24 4.5005
R11415 VSS.n4504 VSS.n24 4.5005
R11416 VSS.n193 VSS.n113 4.5005
R11417 VSS.n195 VSS.n113 4.5005
R11418 VSS.n192 VSS.n113 4.5005
R11419 VSS.n196 VSS.n113 4.5005
R11420 VSS.n191 VSS.n113 4.5005
R11421 VSS.n197 VSS.n113 4.5005
R11422 VSS.n190 VSS.n113 4.5005
R11423 VSS.n198 VSS.n113 4.5005
R11424 VSS.n189 VSS.n113 4.5005
R11425 VSS.n199 VSS.n113 4.5005
R11426 VSS.n188 VSS.n113 4.5005
R11427 VSS.n200 VSS.n113 4.5005
R11428 VSS.n187 VSS.n113 4.5005
R11429 VSS.n201 VSS.n113 4.5005
R11430 VSS.n186 VSS.n113 4.5005
R11431 VSS.n202 VSS.n113 4.5005
R11432 VSS.n185 VSS.n113 4.5005
R11433 VSS.n203 VSS.n113 4.5005
R11434 VSS.n184 VSS.n113 4.5005
R11435 VSS.n204 VSS.n113 4.5005
R11436 VSS.n183 VSS.n113 4.5005
R11437 VSS.n205 VSS.n113 4.5005
R11438 VSS.n182 VSS.n113 4.5005
R11439 VSS.n206 VSS.n113 4.5005
R11440 VSS.n181 VSS.n113 4.5005
R11441 VSS.n207 VSS.n113 4.5005
R11442 VSS.n180 VSS.n113 4.5005
R11443 VSS.n208 VSS.n113 4.5005
R11444 VSS.n179 VSS.n113 4.5005
R11445 VSS.n209 VSS.n113 4.5005
R11446 VSS.n178 VSS.n113 4.5005
R11447 VSS.n210 VSS.n113 4.5005
R11448 VSS.n177 VSS.n113 4.5005
R11449 VSS.n211 VSS.n113 4.5005
R11450 VSS.n176 VSS.n113 4.5005
R11451 VSS.n212 VSS.n113 4.5005
R11452 VSS.n175 VSS.n113 4.5005
R11453 VSS.n213 VSS.n113 4.5005
R11454 VSS.n174 VSS.n113 4.5005
R11455 VSS.n214 VSS.n113 4.5005
R11456 VSS.n173 VSS.n113 4.5005
R11457 VSS.n215 VSS.n113 4.5005
R11458 VSS.n172 VSS.n113 4.5005
R11459 VSS.n216 VSS.n113 4.5005
R11460 VSS.n171 VSS.n113 4.5005
R11461 VSS.n217 VSS.n113 4.5005
R11462 VSS.n170 VSS.n113 4.5005
R11463 VSS.n218 VSS.n113 4.5005
R11464 VSS.n169 VSS.n113 4.5005
R11465 VSS.n219 VSS.n113 4.5005
R11466 VSS.n168 VSS.n113 4.5005
R11467 VSS.n220 VSS.n113 4.5005
R11468 VSS.n167 VSS.n113 4.5005
R11469 VSS.n221 VSS.n113 4.5005
R11470 VSS.n166 VSS.n113 4.5005
R11471 VSS.n222 VSS.n113 4.5005
R11472 VSS.n165 VSS.n113 4.5005
R11473 VSS.n223 VSS.n113 4.5005
R11474 VSS.n164 VSS.n113 4.5005
R11475 VSS.n224 VSS.n113 4.5005
R11476 VSS.n163 VSS.n113 4.5005
R11477 VSS.n225 VSS.n113 4.5005
R11478 VSS.n162 VSS.n113 4.5005
R11479 VSS.n226 VSS.n113 4.5005
R11480 VSS.n161 VSS.n113 4.5005
R11481 VSS.n227 VSS.n113 4.5005
R11482 VSS.n160 VSS.n113 4.5005
R11483 VSS.n228 VSS.n113 4.5005
R11484 VSS.n159 VSS.n113 4.5005
R11485 VSS.n229 VSS.n113 4.5005
R11486 VSS.n158 VSS.n113 4.5005
R11487 VSS.n230 VSS.n113 4.5005
R11488 VSS.n157 VSS.n113 4.5005
R11489 VSS.n231 VSS.n113 4.5005
R11490 VSS.n156 VSS.n113 4.5005
R11491 VSS.n232 VSS.n113 4.5005
R11492 VSS.n155 VSS.n113 4.5005
R11493 VSS.n233 VSS.n113 4.5005
R11494 VSS.n154 VSS.n113 4.5005
R11495 VSS.n234 VSS.n113 4.5005
R11496 VSS.n153 VSS.n113 4.5005
R11497 VSS.n235 VSS.n113 4.5005
R11498 VSS.n4506 VSS.n113 4.5005
R11499 VSS.n236 VSS.n113 4.5005
R11500 VSS.n152 VSS.n113 4.5005
R11501 VSS.n237 VSS.n113 4.5005
R11502 VSS.n151 VSS.n113 4.5005
R11503 VSS.n238 VSS.n113 4.5005
R11504 VSS.n150 VSS.n113 4.5005
R11505 VSS.n239 VSS.n113 4.5005
R11506 VSS.n149 VSS.n113 4.5005
R11507 VSS.n240 VSS.n113 4.5005
R11508 VSS.n148 VSS.n113 4.5005
R11509 VSS.n241 VSS.n113 4.5005
R11510 VSS.n147 VSS.n113 4.5005
R11511 VSS.n242 VSS.n113 4.5005
R11512 VSS.n146 VSS.n113 4.5005
R11513 VSS.n243 VSS.n113 4.5005
R11514 VSS.n145 VSS.n113 4.5005
R11515 VSS.n244 VSS.n113 4.5005
R11516 VSS.n144 VSS.n113 4.5005
R11517 VSS.n245 VSS.n113 4.5005
R11518 VSS.n143 VSS.n113 4.5005
R11519 VSS.n246 VSS.n113 4.5005
R11520 VSS.n142 VSS.n113 4.5005
R11521 VSS.n247 VSS.n113 4.5005
R11522 VSS.n141 VSS.n113 4.5005
R11523 VSS.n248 VSS.n113 4.5005
R11524 VSS.n140 VSS.n113 4.5005
R11525 VSS.n249 VSS.n113 4.5005
R11526 VSS.n139 VSS.n113 4.5005
R11527 VSS.n250 VSS.n113 4.5005
R11528 VSS.n138 VSS.n113 4.5005
R11529 VSS.n251 VSS.n113 4.5005
R11530 VSS.n137 VSS.n113 4.5005
R11531 VSS.n252 VSS.n113 4.5005
R11532 VSS.n136 VSS.n113 4.5005
R11533 VSS.n253 VSS.n113 4.5005
R11534 VSS.n135 VSS.n113 4.5005
R11535 VSS.n254 VSS.n113 4.5005
R11536 VSS.n134 VSS.n113 4.5005
R11537 VSS.n255 VSS.n113 4.5005
R11538 VSS.n133 VSS.n113 4.5005
R11539 VSS.n256 VSS.n113 4.5005
R11540 VSS.n132 VSS.n113 4.5005
R11541 VSS.n4502 VSS.n113 4.5005
R11542 VSS.n4504 VSS.n113 4.5005
R11543 VSS.n193 VSS.n23 4.5005
R11544 VSS.n195 VSS.n23 4.5005
R11545 VSS.n192 VSS.n23 4.5005
R11546 VSS.n196 VSS.n23 4.5005
R11547 VSS.n191 VSS.n23 4.5005
R11548 VSS.n197 VSS.n23 4.5005
R11549 VSS.n190 VSS.n23 4.5005
R11550 VSS.n198 VSS.n23 4.5005
R11551 VSS.n189 VSS.n23 4.5005
R11552 VSS.n199 VSS.n23 4.5005
R11553 VSS.n188 VSS.n23 4.5005
R11554 VSS.n200 VSS.n23 4.5005
R11555 VSS.n187 VSS.n23 4.5005
R11556 VSS.n201 VSS.n23 4.5005
R11557 VSS.n186 VSS.n23 4.5005
R11558 VSS.n202 VSS.n23 4.5005
R11559 VSS.n185 VSS.n23 4.5005
R11560 VSS.n203 VSS.n23 4.5005
R11561 VSS.n184 VSS.n23 4.5005
R11562 VSS.n204 VSS.n23 4.5005
R11563 VSS.n183 VSS.n23 4.5005
R11564 VSS.n205 VSS.n23 4.5005
R11565 VSS.n182 VSS.n23 4.5005
R11566 VSS.n206 VSS.n23 4.5005
R11567 VSS.n181 VSS.n23 4.5005
R11568 VSS.n207 VSS.n23 4.5005
R11569 VSS.n180 VSS.n23 4.5005
R11570 VSS.n208 VSS.n23 4.5005
R11571 VSS.n179 VSS.n23 4.5005
R11572 VSS.n209 VSS.n23 4.5005
R11573 VSS.n178 VSS.n23 4.5005
R11574 VSS.n210 VSS.n23 4.5005
R11575 VSS.n177 VSS.n23 4.5005
R11576 VSS.n211 VSS.n23 4.5005
R11577 VSS.n176 VSS.n23 4.5005
R11578 VSS.n212 VSS.n23 4.5005
R11579 VSS.n175 VSS.n23 4.5005
R11580 VSS.n213 VSS.n23 4.5005
R11581 VSS.n174 VSS.n23 4.5005
R11582 VSS.n214 VSS.n23 4.5005
R11583 VSS.n173 VSS.n23 4.5005
R11584 VSS.n215 VSS.n23 4.5005
R11585 VSS.n172 VSS.n23 4.5005
R11586 VSS.n216 VSS.n23 4.5005
R11587 VSS.n171 VSS.n23 4.5005
R11588 VSS.n217 VSS.n23 4.5005
R11589 VSS.n170 VSS.n23 4.5005
R11590 VSS.n218 VSS.n23 4.5005
R11591 VSS.n169 VSS.n23 4.5005
R11592 VSS.n219 VSS.n23 4.5005
R11593 VSS.n168 VSS.n23 4.5005
R11594 VSS.n220 VSS.n23 4.5005
R11595 VSS.n167 VSS.n23 4.5005
R11596 VSS.n221 VSS.n23 4.5005
R11597 VSS.n166 VSS.n23 4.5005
R11598 VSS.n222 VSS.n23 4.5005
R11599 VSS.n165 VSS.n23 4.5005
R11600 VSS.n223 VSS.n23 4.5005
R11601 VSS.n164 VSS.n23 4.5005
R11602 VSS.n224 VSS.n23 4.5005
R11603 VSS.n163 VSS.n23 4.5005
R11604 VSS.n225 VSS.n23 4.5005
R11605 VSS.n162 VSS.n23 4.5005
R11606 VSS.n226 VSS.n23 4.5005
R11607 VSS.n161 VSS.n23 4.5005
R11608 VSS.n227 VSS.n23 4.5005
R11609 VSS.n160 VSS.n23 4.5005
R11610 VSS.n228 VSS.n23 4.5005
R11611 VSS.n159 VSS.n23 4.5005
R11612 VSS.n229 VSS.n23 4.5005
R11613 VSS.n158 VSS.n23 4.5005
R11614 VSS.n230 VSS.n23 4.5005
R11615 VSS.n157 VSS.n23 4.5005
R11616 VSS.n231 VSS.n23 4.5005
R11617 VSS.n156 VSS.n23 4.5005
R11618 VSS.n232 VSS.n23 4.5005
R11619 VSS.n155 VSS.n23 4.5005
R11620 VSS.n233 VSS.n23 4.5005
R11621 VSS.n154 VSS.n23 4.5005
R11622 VSS.n234 VSS.n23 4.5005
R11623 VSS.n153 VSS.n23 4.5005
R11624 VSS.n235 VSS.n23 4.5005
R11625 VSS.n4506 VSS.n23 4.5005
R11626 VSS.n236 VSS.n23 4.5005
R11627 VSS.n152 VSS.n23 4.5005
R11628 VSS.n237 VSS.n23 4.5005
R11629 VSS.n151 VSS.n23 4.5005
R11630 VSS.n238 VSS.n23 4.5005
R11631 VSS.n150 VSS.n23 4.5005
R11632 VSS.n239 VSS.n23 4.5005
R11633 VSS.n149 VSS.n23 4.5005
R11634 VSS.n240 VSS.n23 4.5005
R11635 VSS.n148 VSS.n23 4.5005
R11636 VSS.n241 VSS.n23 4.5005
R11637 VSS.n147 VSS.n23 4.5005
R11638 VSS.n242 VSS.n23 4.5005
R11639 VSS.n146 VSS.n23 4.5005
R11640 VSS.n243 VSS.n23 4.5005
R11641 VSS.n145 VSS.n23 4.5005
R11642 VSS.n244 VSS.n23 4.5005
R11643 VSS.n144 VSS.n23 4.5005
R11644 VSS.n245 VSS.n23 4.5005
R11645 VSS.n143 VSS.n23 4.5005
R11646 VSS.n246 VSS.n23 4.5005
R11647 VSS.n142 VSS.n23 4.5005
R11648 VSS.n247 VSS.n23 4.5005
R11649 VSS.n141 VSS.n23 4.5005
R11650 VSS.n248 VSS.n23 4.5005
R11651 VSS.n140 VSS.n23 4.5005
R11652 VSS.n249 VSS.n23 4.5005
R11653 VSS.n139 VSS.n23 4.5005
R11654 VSS.n250 VSS.n23 4.5005
R11655 VSS.n138 VSS.n23 4.5005
R11656 VSS.n251 VSS.n23 4.5005
R11657 VSS.n137 VSS.n23 4.5005
R11658 VSS.n252 VSS.n23 4.5005
R11659 VSS.n136 VSS.n23 4.5005
R11660 VSS.n253 VSS.n23 4.5005
R11661 VSS.n135 VSS.n23 4.5005
R11662 VSS.n254 VSS.n23 4.5005
R11663 VSS.n134 VSS.n23 4.5005
R11664 VSS.n255 VSS.n23 4.5005
R11665 VSS.n133 VSS.n23 4.5005
R11666 VSS.n256 VSS.n23 4.5005
R11667 VSS.n132 VSS.n23 4.5005
R11668 VSS.n4502 VSS.n23 4.5005
R11669 VSS.n4504 VSS.n23 4.5005
R11670 VSS.n193 VSS.n114 4.5005
R11671 VSS.n195 VSS.n114 4.5005
R11672 VSS.n192 VSS.n114 4.5005
R11673 VSS.n196 VSS.n114 4.5005
R11674 VSS.n191 VSS.n114 4.5005
R11675 VSS.n197 VSS.n114 4.5005
R11676 VSS.n190 VSS.n114 4.5005
R11677 VSS.n198 VSS.n114 4.5005
R11678 VSS.n189 VSS.n114 4.5005
R11679 VSS.n199 VSS.n114 4.5005
R11680 VSS.n188 VSS.n114 4.5005
R11681 VSS.n200 VSS.n114 4.5005
R11682 VSS.n187 VSS.n114 4.5005
R11683 VSS.n201 VSS.n114 4.5005
R11684 VSS.n186 VSS.n114 4.5005
R11685 VSS.n202 VSS.n114 4.5005
R11686 VSS.n185 VSS.n114 4.5005
R11687 VSS.n203 VSS.n114 4.5005
R11688 VSS.n184 VSS.n114 4.5005
R11689 VSS.n204 VSS.n114 4.5005
R11690 VSS.n183 VSS.n114 4.5005
R11691 VSS.n205 VSS.n114 4.5005
R11692 VSS.n182 VSS.n114 4.5005
R11693 VSS.n206 VSS.n114 4.5005
R11694 VSS.n181 VSS.n114 4.5005
R11695 VSS.n207 VSS.n114 4.5005
R11696 VSS.n180 VSS.n114 4.5005
R11697 VSS.n208 VSS.n114 4.5005
R11698 VSS.n179 VSS.n114 4.5005
R11699 VSS.n209 VSS.n114 4.5005
R11700 VSS.n178 VSS.n114 4.5005
R11701 VSS.n210 VSS.n114 4.5005
R11702 VSS.n177 VSS.n114 4.5005
R11703 VSS.n211 VSS.n114 4.5005
R11704 VSS.n176 VSS.n114 4.5005
R11705 VSS.n212 VSS.n114 4.5005
R11706 VSS.n175 VSS.n114 4.5005
R11707 VSS.n213 VSS.n114 4.5005
R11708 VSS.n174 VSS.n114 4.5005
R11709 VSS.n214 VSS.n114 4.5005
R11710 VSS.n173 VSS.n114 4.5005
R11711 VSS.n215 VSS.n114 4.5005
R11712 VSS.n172 VSS.n114 4.5005
R11713 VSS.n216 VSS.n114 4.5005
R11714 VSS.n171 VSS.n114 4.5005
R11715 VSS.n217 VSS.n114 4.5005
R11716 VSS.n170 VSS.n114 4.5005
R11717 VSS.n218 VSS.n114 4.5005
R11718 VSS.n169 VSS.n114 4.5005
R11719 VSS.n219 VSS.n114 4.5005
R11720 VSS.n168 VSS.n114 4.5005
R11721 VSS.n220 VSS.n114 4.5005
R11722 VSS.n167 VSS.n114 4.5005
R11723 VSS.n221 VSS.n114 4.5005
R11724 VSS.n166 VSS.n114 4.5005
R11725 VSS.n222 VSS.n114 4.5005
R11726 VSS.n165 VSS.n114 4.5005
R11727 VSS.n223 VSS.n114 4.5005
R11728 VSS.n164 VSS.n114 4.5005
R11729 VSS.n224 VSS.n114 4.5005
R11730 VSS.n163 VSS.n114 4.5005
R11731 VSS.n225 VSS.n114 4.5005
R11732 VSS.n162 VSS.n114 4.5005
R11733 VSS.n226 VSS.n114 4.5005
R11734 VSS.n161 VSS.n114 4.5005
R11735 VSS.n227 VSS.n114 4.5005
R11736 VSS.n160 VSS.n114 4.5005
R11737 VSS.n228 VSS.n114 4.5005
R11738 VSS.n159 VSS.n114 4.5005
R11739 VSS.n229 VSS.n114 4.5005
R11740 VSS.n158 VSS.n114 4.5005
R11741 VSS.n230 VSS.n114 4.5005
R11742 VSS.n157 VSS.n114 4.5005
R11743 VSS.n231 VSS.n114 4.5005
R11744 VSS.n156 VSS.n114 4.5005
R11745 VSS.n232 VSS.n114 4.5005
R11746 VSS.n155 VSS.n114 4.5005
R11747 VSS.n233 VSS.n114 4.5005
R11748 VSS.n154 VSS.n114 4.5005
R11749 VSS.n234 VSS.n114 4.5005
R11750 VSS.n153 VSS.n114 4.5005
R11751 VSS.n235 VSS.n114 4.5005
R11752 VSS.n4506 VSS.n114 4.5005
R11753 VSS.n236 VSS.n114 4.5005
R11754 VSS.n152 VSS.n114 4.5005
R11755 VSS.n237 VSS.n114 4.5005
R11756 VSS.n151 VSS.n114 4.5005
R11757 VSS.n238 VSS.n114 4.5005
R11758 VSS.n150 VSS.n114 4.5005
R11759 VSS.n239 VSS.n114 4.5005
R11760 VSS.n149 VSS.n114 4.5005
R11761 VSS.n240 VSS.n114 4.5005
R11762 VSS.n148 VSS.n114 4.5005
R11763 VSS.n241 VSS.n114 4.5005
R11764 VSS.n147 VSS.n114 4.5005
R11765 VSS.n242 VSS.n114 4.5005
R11766 VSS.n146 VSS.n114 4.5005
R11767 VSS.n243 VSS.n114 4.5005
R11768 VSS.n145 VSS.n114 4.5005
R11769 VSS.n244 VSS.n114 4.5005
R11770 VSS.n144 VSS.n114 4.5005
R11771 VSS.n245 VSS.n114 4.5005
R11772 VSS.n143 VSS.n114 4.5005
R11773 VSS.n246 VSS.n114 4.5005
R11774 VSS.n142 VSS.n114 4.5005
R11775 VSS.n247 VSS.n114 4.5005
R11776 VSS.n141 VSS.n114 4.5005
R11777 VSS.n248 VSS.n114 4.5005
R11778 VSS.n140 VSS.n114 4.5005
R11779 VSS.n249 VSS.n114 4.5005
R11780 VSS.n139 VSS.n114 4.5005
R11781 VSS.n250 VSS.n114 4.5005
R11782 VSS.n138 VSS.n114 4.5005
R11783 VSS.n251 VSS.n114 4.5005
R11784 VSS.n137 VSS.n114 4.5005
R11785 VSS.n252 VSS.n114 4.5005
R11786 VSS.n136 VSS.n114 4.5005
R11787 VSS.n253 VSS.n114 4.5005
R11788 VSS.n135 VSS.n114 4.5005
R11789 VSS.n254 VSS.n114 4.5005
R11790 VSS.n134 VSS.n114 4.5005
R11791 VSS.n255 VSS.n114 4.5005
R11792 VSS.n133 VSS.n114 4.5005
R11793 VSS.n256 VSS.n114 4.5005
R11794 VSS.n132 VSS.n114 4.5005
R11795 VSS.n4502 VSS.n114 4.5005
R11796 VSS.n4504 VSS.n114 4.5005
R11797 VSS.n193 VSS.n22 4.5005
R11798 VSS.n195 VSS.n22 4.5005
R11799 VSS.n192 VSS.n22 4.5005
R11800 VSS.n196 VSS.n22 4.5005
R11801 VSS.n191 VSS.n22 4.5005
R11802 VSS.n197 VSS.n22 4.5005
R11803 VSS.n190 VSS.n22 4.5005
R11804 VSS.n198 VSS.n22 4.5005
R11805 VSS.n189 VSS.n22 4.5005
R11806 VSS.n199 VSS.n22 4.5005
R11807 VSS.n188 VSS.n22 4.5005
R11808 VSS.n200 VSS.n22 4.5005
R11809 VSS.n187 VSS.n22 4.5005
R11810 VSS.n201 VSS.n22 4.5005
R11811 VSS.n186 VSS.n22 4.5005
R11812 VSS.n202 VSS.n22 4.5005
R11813 VSS.n185 VSS.n22 4.5005
R11814 VSS.n203 VSS.n22 4.5005
R11815 VSS.n184 VSS.n22 4.5005
R11816 VSS.n204 VSS.n22 4.5005
R11817 VSS.n183 VSS.n22 4.5005
R11818 VSS.n205 VSS.n22 4.5005
R11819 VSS.n182 VSS.n22 4.5005
R11820 VSS.n206 VSS.n22 4.5005
R11821 VSS.n181 VSS.n22 4.5005
R11822 VSS.n207 VSS.n22 4.5005
R11823 VSS.n180 VSS.n22 4.5005
R11824 VSS.n208 VSS.n22 4.5005
R11825 VSS.n179 VSS.n22 4.5005
R11826 VSS.n209 VSS.n22 4.5005
R11827 VSS.n178 VSS.n22 4.5005
R11828 VSS.n210 VSS.n22 4.5005
R11829 VSS.n177 VSS.n22 4.5005
R11830 VSS.n211 VSS.n22 4.5005
R11831 VSS.n176 VSS.n22 4.5005
R11832 VSS.n212 VSS.n22 4.5005
R11833 VSS.n175 VSS.n22 4.5005
R11834 VSS.n213 VSS.n22 4.5005
R11835 VSS.n174 VSS.n22 4.5005
R11836 VSS.n214 VSS.n22 4.5005
R11837 VSS.n173 VSS.n22 4.5005
R11838 VSS.n215 VSS.n22 4.5005
R11839 VSS.n172 VSS.n22 4.5005
R11840 VSS.n216 VSS.n22 4.5005
R11841 VSS.n171 VSS.n22 4.5005
R11842 VSS.n217 VSS.n22 4.5005
R11843 VSS.n170 VSS.n22 4.5005
R11844 VSS.n218 VSS.n22 4.5005
R11845 VSS.n169 VSS.n22 4.5005
R11846 VSS.n219 VSS.n22 4.5005
R11847 VSS.n168 VSS.n22 4.5005
R11848 VSS.n220 VSS.n22 4.5005
R11849 VSS.n167 VSS.n22 4.5005
R11850 VSS.n221 VSS.n22 4.5005
R11851 VSS.n166 VSS.n22 4.5005
R11852 VSS.n222 VSS.n22 4.5005
R11853 VSS.n165 VSS.n22 4.5005
R11854 VSS.n223 VSS.n22 4.5005
R11855 VSS.n164 VSS.n22 4.5005
R11856 VSS.n224 VSS.n22 4.5005
R11857 VSS.n163 VSS.n22 4.5005
R11858 VSS.n225 VSS.n22 4.5005
R11859 VSS.n162 VSS.n22 4.5005
R11860 VSS.n226 VSS.n22 4.5005
R11861 VSS.n161 VSS.n22 4.5005
R11862 VSS.n227 VSS.n22 4.5005
R11863 VSS.n160 VSS.n22 4.5005
R11864 VSS.n228 VSS.n22 4.5005
R11865 VSS.n159 VSS.n22 4.5005
R11866 VSS.n229 VSS.n22 4.5005
R11867 VSS.n158 VSS.n22 4.5005
R11868 VSS.n230 VSS.n22 4.5005
R11869 VSS.n157 VSS.n22 4.5005
R11870 VSS.n231 VSS.n22 4.5005
R11871 VSS.n156 VSS.n22 4.5005
R11872 VSS.n232 VSS.n22 4.5005
R11873 VSS.n155 VSS.n22 4.5005
R11874 VSS.n233 VSS.n22 4.5005
R11875 VSS.n154 VSS.n22 4.5005
R11876 VSS.n234 VSS.n22 4.5005
R11877 VSS.n153 VSS.n22 4.5005
R11878 VSS.n235 VSS.n22 4.5005
R11879 VSS.n4506 VSS.n22 4.5005
R11880 VSS.n236 VSS.n22 4.5005
R11881 VSS.n152 VSS.n22 4.5005
R11882 VSS.n237 VSS.n22 4.5005
R11883 VSS.n151 VSS.n22 4.5005
R11884 VSS.n238 VSS.n22 4.5005
R11885 VSS.n150 VSS.n22 4.5005
R11886 VSS.n239 VSS.n22 4.5005
R11887 VSS.n149 VSS.n22 4.5005
R11888 VSS.n240 VSS.n22 4.5005
R11889 VSS.n148 VSS.n22 4.5005
R11890 VSS.n241 VSS.n22 4.5005
R11891 VSS.n147 VSS.n22 4.5005
R11892 VSS.n242 VSS.n22 4.5005
R11893 VSS.n146 VSS.n22 4.5005
R11894 VSS.n243 VSS.n22 4.5005
R11895 VSS.n145 VSS.n22 4.5005
R11896 VSS.n244 VSS.n22 4.5005
R11897 VSS.n144 VSS.n22 4.5005
R11898 VSS.n245 VSS.n22 4.5005
R11899 VSS.n143 VSS.n22 4.5005
R11900 VSS.n246 VSS.n22 4.5005
R11901 VSS.n142 VSS.n22 4.5005
R11902 VSS.n247 VSS.n22 4.5005
R11903 VSS.n141 VSS.n22 4.5005
R11904 VSS.n248 VSS.n22 4.5005
R11905 VSS.n140 VSS.n22 4.5005
R11906 VSS.n249 VSS.n22 4.5005
R11907 VSS.n139 VSS.n22 4.5005
R11908 VSS.n250 VSS.n22 4.5005
R11909 VSS.n138 VSS.n22 4.5005
R11910 VSS.n251 VSS.n22 4.5005
R11911 VSS.n137 VSS.n22 4.5005
R11912 VSS.n252 VSS.n22 4.5005
R11913 VSS.n136 VSS.n22 4.5005
R11914 VSS.n253 VSS.n22 4.5005
R11915 VSS.n135 VSS.n22 4.5005
R11916 VSS.n254 VSS.n22 4.5005
R11917 VSS.n134 VSS.n22 4.5005
R11918 VSS.n255 VSS.n22 4.5005
R11919 VSS.n133 VSS.n22 4.5005
R11920 VSS.n256 VSS.n22 4.5005
R11921 VSS.n132 VSS.n22 4.5005
R11922 VSS.n4502 VSS.n22 4.5005
R11923 VSS.n4504 VSS.n22 4.5005
R11924 VSS.n193 VSS.n115 4.5005
R11925 VSS.n195 VSS.n115 4.5005
R11926 VSS.n192 VSS.n115 4.5005
R11927 VSS.n196 VSS.n115 4.5005
R11928 VSS.n191 VSS.n115 4.5005
R11929 VSS.n197 VSS.n115 4.5005
R11930 VSS.n190 VSS.n115 4.5005
R11931 VSS.n198 VSS.n115 4.5005
R11932 VSS.n189 VSS.n115 4.5005
R11933 VSS.n199 VSS.n115 4.5005
R11934 VSS.n188 VSS.n115 4.5005
R11935 VSS.n200 VSS.n115 4.5005
R11936 VSS.n187 VSS.n115 4.5005
R11937 VSS.n201 VSS.n115 4.5005
R11938 VSS.n186 VSS.n115 4.5005
R11939 VSS.n202 VSS.n115 4.5005
R11940 VSS.n185 VSS.n115 4.5005
R11941 VSS.n203 VSS.n115 4.5005
R11942 VSS.n184 VSS.n115 4.5005
R11943 VSS.n204 VSS.n115 4.5005
R11944 VSS.n183 VSS.n115 4.5005
R11945 VSS.n205 VSS.n115 4.5005
R11946 VSS.n182 VSS.n115 4.5005
R11947 VSS.n206 VSS.n115 4.5005
R11948 VSS.n181 VSS.n115 4.5005
R11949 VSS.n207 VSS.n115 4.5005
R11950 VSS.n180 VSS.n115 4.5005
R11951 VSS.n208 VSS.n115 4.5005
R11952 VSS.n179 VSS.n115 4.5005
R11953 VSS.n209 VSS.n115 4.5005
R11954 VSS.n178 VSS.n115 4.5005
R11955 VSS.n210 VSS.n115 4.5005
R11956 VSS.n177 VSS.n115 4.5005
R11957 VSS.n211 VSS.n115 4.5005
R11958 VSS.n176 VSS.n115 4.5005
R11959 VSS.n212 VSS.n115 4.5005
R11960 VSS.n175 VSS.n115 4.5005
R11961 VSS.n213 VSS.n115 4.5005
R11962 VSS.n174 VSS.n115 4.5005
R11963 VSS.n214 VSS.n115 4.5005
R11964 VSS.n173 VSS.n115 4.5005
R11965 VSS.n215 VSS.n115 4.5005
R11966 VSS.n172 VSS.n115 4.5005
R11967 VSS.n216 VSS.n115 4.5005
R11968 VSS.n171 VSS.n115 4.5005
R11969 VSS.n217 VSS.n115 4.5005
R11970 VSS.n170 VSS.n115 4.5005
R11971 VSS.n218 VSS.n115 4.5005
R11972 VSS.n169 VSS.n115 4.5005
R11973 VSS.n219 VSS.n115 4.5005
R11974 VSS.n168 VSS.n115 4.5005
R11975 VSS.n220 VSS.n115 4.5005
R11976 VSS.n167 VSS.n115 4.5005
R11977 VSS.n221 VSS.n115 4.5005
R11978 VSS.n166 VSS.n115 4.5005
R11979 VSS.n222 VSS.n115 4.5005
R11980 VSS.n165 VSS.n115 4.5005
R11981 VSS.n223 VSS.n115 4.5005
R11982 VSS.n164 VSS.n115 4.5005
R11983 VSS.n224 VSS.n115 4.5005
R11984 VSS.n163 VSS.n115 4.5005
R11985 VSS.n225 VSS.n115 4.5005
R11986 VSS.n162 VSS.n115 4.5005
R11987 VSS.n226 VSS.n115 4.5005
R11988 VSS.n161 VSS.n115 4.5005
R11989 VSS.n227 VSS.n115 4.5005
R11990 VSS.n160 VSS.n115 4.5005
R11991 VSS.n228 VSS.n115 4.5005
R11992 VSS.n159 VSS.n115 4.5005
R11993 VSS.n229 VSS.n115 4.5005
R11994 VSS.n158 VSS.n115 4.5005
R11995 VSS.n230 VSS.n115 4.5005
R11996 VSS.n157 VSS.n115 4.5005
R11997 VSS.n231 VSS.n115 4.5005
R11998 VSS.n156 VSS.n115 4.5005
R11999 VSS.n232 VSS.n115 4.5005
R12000 VSS.n155 VSS.n115 4.5005
R12001 VSS.n233 VSS.n115 4.5005
R12002 VSS.n154 VSS.n115 4.5005
R12003 VSS.n234 VSS.n115 4.5005
R12004 VSS.n153 VSS.n115 4.5005
R12005 VSS.n235 VSS.n115 4.5005
R12006 VSS.n4506 VSS.n115 4.5005
R12007 VSS.n236 VSS.n115 4.5005
R12008 VSS.n152 VSS.n115 4.5005
R12009 VSS.n237 VSS.n115 4.5005
R12010 VSS.n151 VSS.n115 4.5005
R12011 VSS.n238 VSS.n115 4.5005
R12012 VSS.n150 VSS.n115 4.5005
R12013 VSS.n239 VSS.n115 4.5005
R12014 VSS.n149 VSS.n115 4.5005
R12015 VSS.n240 VSS.n115 4.5005
R12016 VSS.n148 VSS.n115 4.5005
R12017 VSS.n241 VSS.n115 4.5005
R12018 VSS.n147 VSS.n115 4.5005
R12019 VSS.n242 VSS.n115 4.5005
R12020 VSS.n146 VSS.n115 4.5005
R12021 VSS.n243 VSS.n115 4.5005
R12022 VSS.n145 VSS.n115 4.5005
R12023 VSS.n244 VSS.n115 4.5005
R12024 VSS.n144 VSS.n115 4.5005
R12025 VSS.n245 VSS.n115 4.5005
R12026 VSS.n143 VSS.n115 4.5005
R12027 VSS.n246 VSS.n115 4.5005
R12028 VSS.n142 VSS.n115 4.5005
R12029 VSS.n247 VSS.n115 4.5005
R12030 VSS.n141 VSS.n115 4.5005
R12031 VSS.n248 VSS.n115 4.5005
R12032 VSS.n140 VSS.n115 4.5005
R12033 VSS.n249 VSS.n115 4.5005
R12034 VSS.n139 VSS.n115 4.5005
R12035 VSS.n250 VSS.n115 4.5005
R12036 VSS.n138 VSS.n115 4.5005
R12037 VSS.n251 VSS.n115 4.5005
R12038 VSS.n137 VSS.n115 4.5005
R12039 VSS.n252 VSS.n115 4.5005
R12040 VSS.n136 VSS.n115 4.5005
R12041 VSS.n253 VSS.n115 4.5005
R12042 VSS.n135 VSS.n115 4.5005
R12043 VSS.n254 VSS.n115 4.5005
R12044 VSS.n134 VSS.n115 4.5005
R12045 VSS.n255 VSS.n115 4.5005
R12046 VSS.n133 VSS.n115 4.5005
R12047 VSS.n256 VSS.n115 4.5005
R12048 VSS.n132 VSS.n115 4.5005
R12049 VSS.n4502 VSS.n115 4.5005
R12050 VSS.n4504 VSS.n115 4.5005
R12051 VSS.n193 VSS.n21 4.5005
R12052 VSS.n195 VSS.n21 4.5005
R12053 VSS.n192 VSS.n21 4.5005
R12054 VSS.n196 VSS.n21 4.5005
R12055 VSS.n191 VSS.n21 4.5005
R12056 VSS.n197 VSS.n21 4.5005
R12057 VSS.n190 VSS.n21 4.5005
R12058 VSS.n198 VSS.n21 4.5005
R12059 VSS.n189 VSS.n21 4.5005
R12060 VSS.n199 VSS.n21 4.5005
R12061 VSS.n188 VSS.n21 4.5005
R12062 VSS.n200 VSS.n21 4.5005
R12063 VSS.n187 VSS.n21 4.5005
R12064 VSS.n201 VSS.n21 4.5005
R12065 VSS.n186 VSS.n21 4.5005
R12066 VSS.n202 VSS.n21 4.5005
R12067 VSS.n185 VSS.n21 4.5005
R12068 VSS.n203 VSS.n21 4.5005
R12069 VSS.n184 VSS.n21 4.5005
R12070 VSS.n204 VSS.n21 4.5005
R12071 VSS.n183 VSS.n21 4.5005
R12072 VSS.n205 VSS.n21 4.5005
R12073 VSS.n182 VSS.n21 4.5005
R12074 VSS.n206 VSS.n21 4.5005
R12075 VSS.n181 VSS.n21 4.5005
R12076 VSS.n207 VSS.n21 4.5005
R12077 VSS.n180 VSS.n21 4.5005
R12078 VSS.n208 VSS.n21 4.5005
R12079 VSS.n179 VSS.n21 4.5005
R12080 VSS.n209 VSS.n21 4.5005
R12081 VSS.n178 VSS.n21 4.5005
R12082 VSS.n210 VSS.n21 4.5005
R12083 VSS.n177 VSS.n21 4.5005
R12084 VSS.n211 VSS.n21 4.5005
R12085 VSS.n176 VSS.n21 4.5005
R12086 VSS.n212 VSS.n21 4.5005
R12087 VSS.n175 VSS.n21 4.5005
R12088 VSS.n213 VSS.n21 4.5005
R12089 VSS.n174 VSS.n21 4.5005
R12090 VSS.n214 VSS.n21 4.5005
R12091 VSS.n173 VSS.n21 4.5005
R12092 VSS.n215 VSS.n21 4.5005
R12093 VSS.n172 VSS.n21 4.5005
R12094 VSS.n216 VSS.n21 4.5005
R12095 VSS.n171 VSS.n21 4.5005
R12096 VSS.n217 VSS.n21 4.5005
R12097 VSS.n170 VSS.n21 4.5005
R12098 VSS.n218 VSS.n21 4.5005
R12099 VSS.n169 VSS.n21 4.5005
R12100 VSS.n219 VSS.n21 4.5005
R12101 VSS.n168 VSS.n21 4.5005
R12102 VSS.n220 VSS.n21 4.5005
R12103 VSS.n167 VSS.n21 4.5005
R12104 VSS.n221 VSS.n21 4.5005
R12105 VSS.n166 VSS.n21 4.5005
R12106 VSS.n222 VSS.n21 4.5005
R12107 VSS.n165 VSS.n21 4.5005
R12108 VSS.n223 VSS.n21 4.5005
R12109 VSS.n164 VSS.n21 4.5005
R12110 VSS.n224 VSS.n21 4.5005
R12111 VSS.n163 VSS.n21 4.5005
R12112 VSS.n225 VSS.n21 4.5005
R12113 VSS.n162 VSS.n21 4.5005
R12114 VSS.n226 VSS.n21 4.5005
R12115 VSS.n161 VSS.n21 4.5005
R12116 VSS.n227 VSS.n21 4.5005
R12117 VSS.n160 VSS.n21 4.5005
R12118 VSS.n228 VSS.n21 4.5005
R12119 VSS.n159 VSS.n21 4.5005
R12120 VSS.n229 VSS.n21 4.5005
R12121 VSS.n158 VSS.n21 4.5005
R12122 VSS.n230 VSS.n21 4.5005
R12123 VSS.n157 VSS.n21 4.5005
R12124 VSS.n231 VSS.n21 4.5005
R12125 VSS.n156 VSS.n21 4.5005
R12126 VSS.n232 VSS.n21 4.5005
R12127 VSS.n155 VSS.n21 4.5005
R12128 VSS.n233 VSS.n21 4.5005
R12129 VSS.n154 VSS.n21 4.5005
R12130 VSS.n234 VSS.n21 4.5005
R12131 VSS.n153 VSS.n21 4.5005
R12132 VSS.n235 VSS.n21 4.5005
R12133 VSS.n4506 VSS.n21 4.5005
R12134 VSS.n236 VSS.n21 4.5005
R12135 VSS.n152 VSS.n21 4.5005
R12136 VSS.n237 VSS.n21 4.5005
R12137 VSS.n151 VSS.n21 4.5005
R12138 VSS.n238 VSS.n21 4.5005
R12139 VSS.n150 VSS.n21 4.5005
R12140 VSS.n239 VSS.n21 4.5005
R12141 VSS.n149 VSS.n21 4.5005
R12142 VSS.n240 VSS.n21 4.5005
R12143 VSS.n148 VSS.n21 4.5005
R12144 VSS.n241 VSS.n21 4.5005
R12145 VSS.n147 VSS.n21 4.5005
R12146 VSS.n242 VSS.n21 4.5005
R12147 VSS.n146 VSS.n21 4.5005
R12148 VSS.n243 VSS.n21 4.5005
R12149 VSS.n145 VSS.n21 4.5005
R12150 VSS.n244 VSS.n21 4.5005
R12151 VSS.n144 VSS.n21 4.5005
R12152 VSS.n245 VSS.n21 4.5005
R12153 VSS.n143 VSS.n21 4.5005
R12154 VSS.n246 VSS.n21 4.5005
R12155 VSS.n142 VSS.n21 4.5005
R12156 VSS.n247 VSS.n21 4.5005
R12157 VSS.n141 VSS.n21 4.5005
R12158 VSS.n248 VSS.n21 4.5005
R12159 VSS.n140 VSS.n21 4.5005
R12160 VSS.n249 VSS.n21 4.5005
R12161 VSS.n139 VSS.n21 4.5005
R12162 VSS.n250 VSS.n21 4.5005
R12163 VSS.n138 VSS.n21 4.5005
R12164 VSS.n251 VSS.n21 4.5005
R12165 VSS.n137 VSS.n21 4.5005
R12166 VSS.n252 VSS.n21 4.5005
R12167 VSS.n136 VSS.n21 4.5005
R12168 VSS.n253 VSS.n21 4.5005
R12169 VSS.n135 VSS.n21 4.5005
R12170 VSS.n254 VSS.n21 4.5005
R12171 VSS.n134 VSS.n21 4.5005
R12172 VSS.n255 VSS.n21 4.5005
R12173 VSS.n133 VSS.n21 4.5005
R12174 VSS.n256 VSS.n21 4.5005
R12175 VSS.n132 VSS.n21 4.5005
R12176 VSS.n4502 VSS.n21 4.5005
R12177 VSS.n4504 VSS.n21 4.5005
R12178 VSS.n193 VSS.n116 4.5005
R12179 VSS.n195 VSS.n116 4.5005
R12180 VSS.n192 VSS.n116 4.5005
R12181 VSS.n196 VSS.n116 4.5005
R12182 VSS.n191 VSS.n116 4.5005
R12183 VSS.n197 VSS.n116 4.5005
R12184 VSS.n190 VSS.n116 4.5005
R12185 VSS.n198 VSS.n116 4.5005
R12186 VSS.n189 VSS.n116 4.5005
R12187 VSS.n199 VSS.n116 4.5005
R12188 VSS.n188 VSS.n116 4.5005
R12189 VSS.n200 VSS.n116 4.5005
R12190 VSS.n187 VSS.n116 4.5005
R12191 VSS.n201 VSS.n116 4.5005
R12192 VSS.n186 VSS.n116 4.5005
R12193 VSS.n202 VSS.n116 4.5005
R12194 VSS.n185 VSS.n116 4.5005
R12195 VSS.n203 VSS.n116 4.5005
R12196 VSS.n184 VSS.n116 4.5005
R12197 VSS.n204 VSS.n116 4.5005
R12198 VSS.n183 VSS.n116 4.5005
R12199 VSS.n205 VSS.n116 4.5005
R12200 VSS.n182 VSS.n116 4.5005
R12201 VSS.n206 VSS.n116 4.5005
R12202 VSS.n181 VSS.n116 4.5005
R12203 VSS.n207 VSS.n116 4.5005
R12204 VSS.n180 VSS.n116 4.5005
R12205 VSS.n208 VSS.n116 4.5005
R12206 VSS.n179 VSS.n116 4.5005
R12207 VSS.n209 VSS.n116 4.5005
R12208 VSS.n178 VSS.n116 4.5005
R12209 VSS.n210 VSS.n116 4.5005
R12210 VSS.n177 VSS.n116 4.5005
R12211 VSS.n211 VSS.n116 4.5005
R12212 VSS.n176 VSS.n116 4.5005
R12213 VSS.n212 VSS.n116 4.5005
R12214 VSS.n175 VSS.n116 4.5005
R12215 VSS.n213 VSS.n116 4.5005
R12216 VSS.n174 VSS.n116 4.5005
R12217 VSS.n214 VSS.n116 4.5005
R12218 VSS.n173 VSS.n116 4.5005
R12219 VSS.n215 VSS.n116 4.5005
R12220 VSS.n172 VSS.n116 4.5005
R12221 VSS.n216 VSS.n116 4.5005
R12222 VSS.n171 VSS.n116 4.5005
R12223 VSS.n217 VSS.n116 4.5005
R12224 VSS.n170 VSS.n116 4.5005
R12225 VSS.n218 VSS.n116 4.5005
R12226 VSS.n169 VSS.n116 4.5005
R12227 VSS.n219 VSS.n116 4.5005
R12228 VSS.n168 VSS.n116 4.5005
R12229 VSS.n220 VSS.n116 4.5005
R12230 VSS.n167 VSS.n116 4.5005
R12231 VSS.n221 VSS.n116 4.5005
R12232 VSS.n166 VSS.n116 4.5005
R12233 VSS.n222 VSS.n116 4.5005
R12234 VSS.n165 VSS.n116 4.5005
R12235 VSS.n223 VSS.n116 4.5005
R12236 VSS.n164 VSS.n116 4.5005
R12237 VSS.n224 VSS.n116 4.5005
R12238 VSS.n163 VSS.n116 4.5005
R12239 VSS.n225 VSS.n116 4.5005
R12240 VSS.n162 VSS.n116 4.5005
R12241 VSS.n226 VSS.n116 4.5005
R12242 VSS.n161 VSS.n116 4.5005
R12243 VSS.n227 VSS.n116 4.5005
R12244 VSS.n160 VSS.n116 4.5005
R12245 VSS.n228 VSS.n116 4.5005
R12246 VSS.n159 VSS.n116 4.5005
R12247 VSS.n229 VSS.n116 4.5005
R12248 VSS.n158 VSS.n116 4.5005
R12249 VSS.n230 VSS.n116 4.5005
R12250 VSS.n157 VSS.n116 4.5005
R12251 VSS.n231 VSS.n116 4.5005
R12252 VSS.n156 VSS.n116 4.5005
R12253 VSS.n232 VSS.n116 4.5005
R12254 VSS.n155 VSS.n116 4.5005
R12255 VSS.n233 VSS.n116 4.5005
R12256 VSS.n154 VSS.n116 4.5005
R12257 VSS.n234 VSS.n116 4.5005
R12258 VSS.n153 VSS.n116 4.5005
R12259 VSS.n235 VSS.n116 4.5005
R12260 VSS.n4506 VSS.n116 4.5005
R12261 VSS.n236 VSS.n116 4.5005
R12262 VSS.n152 VSS.n116 4.5005
R12263 VSS.n237 VSS.n116 4.5005
R12264 VSS.n151 VSS.n116 4.5005
R12265 VSS.n238 VSS.n116 4.5005
R12266 VSS.n150 VSS.n116 4.5005
R12267 VSS.n239 VSS.n116 4.5005
R12268 VSS.n149 VSS.n116 4.5005
R12269 VSS.n240 VSS.n116 4.5005
R12270 VSS.n148 VSS.n116 4.5005
R12271 VSS.n241 VSS.n116 4.5005
R12272 VSS.n147 VSS.n116 4.5005
R12273 VSS.n242 VSS.n116 4.5005
R12274 VSS.n146 VSS.n116 4.5005
R12275 VSS.n243 VSS.n116 4.5005
R12276 VSS.n145 VSS.n116 4.5005
R12277 VSS.n244 VSS.n116 4.5005
R12278 VSS.n144 VSS.n116 4.5005
R12279 VSS.n245 VSS.n116 4.5005
R12280 VSS.n143 VSS.n116 4.5005
R12281 VSS.n246 VSS.n116 4.5005
R12282 VSS.n142 VSS.n116 4.5005
R12283 VSS.n247 VSS.n116 4.5005
R12284 VSS.n141 VSS.n116 4.5005
R12285 VSS.n248 VSS.n116 4.5005
R12286 VSS.n140 VSS.n116 4.5005
R12287 VSS.n249 VSS.n116 4.5005
R12288 VSS.n139 VSS.n116 4.5005
R12289 VSS.n250 VSS.n116 4.5005
R12290 VSS.n138 VSS.n116 4.5005
R12291 VSS.n251 VSS.n116 4.5005
R12292 VSS.n137 VSS.n116 4.5005
R12293 VSS.n252 VSS.n116 4.5005
R12294 VSS.n136 VSS.n116 4.5005
R12295 VSS.n253 VSS.n116 4.5005
R12296 VSS.n135 VSS.n116 4.5005
R12297 VSS.n254 VSS.n116 4.5005
R12298 VSS.n134 VSS.n116 4.5005
R12299 VSS.n255 VSS.n116 4.5005
R12300 VSS.n133 VSS.n116 4.5005
R12301 VSS.n256 VSS.n116 4.5005
R12302 VSS.n132 VSS.n116 4.5005
R12303 VSS.n4502 VSS.n116 4.5005
R12304 VSS.n4504 VSS.n116 4.5005
R12305 VSS.n193 VSS.n20 4.5005
R12306 VSS.n195 VSS.n20 4.5005
R12307 VSS.n192 VSS.n20 4.5005
R12308 VSS.n196 VSS.n20 4.5005
R12309 VSS.n191 VSS.n20 4.5005
R12310 VSS.n197 VSS.n20 4.5005
R12311 VSS.n190 VSS.n20 4.5005
R12312 VSS.n198 VSS.n20 4.5005
R12313 VSS.n189 VSS.n20 4.5005
R12314 VSS.n199 VSS.n20 4.5005
R12315 VSS.n188 VSS.n20 4.5005
R12316 VSS.n200 VSS.n20 4.5005
R12317 VSS.n187 VSS.n20 4.5005
R12318 VSS.n201 VSS.n20 4.5005
R12319 VSS.n186 VSS.n20 4.5005
R12320 VSS.n202 VSS.n20 4.5005
R12321 VSS.n185 VSS.n20 4.5005
R12322 VSS.n203 VSS.n20 4.5005
R12323 VSS.n184 VSS.n20 4.5005
R12324 VSS.n204 VSS.n20 4.5005
R12325 VSS.n183 VSS.n20 4.5005
R12326 VSS.n205 VSS.n20 4.5005
R12327 VSS.n182 VSS.n20 4.5005
R12328 VSS.n206 VSS.n20 4.5005
R12329 VSS.n181 VSS.n20 4.5005
R12330 VSS.n207 VSS.n20 4.5005
R12331 VSS.n180 VSS.n20 4.5005
R12332 VSS.n208 VSS.n20 4.5005
R12333 VSS.n179 VSS.n20 4.5005
R12334 VSS.n209 VSS.n20 4.5005
R12335 VSS.n178 VSS.n20 4.5005
R12336 VSS.n210 VSS.n20 4.5005
R12337 VSS.n177 VSS.n20 4.5005
R12338 VSS.n211 VSS.n20 4.5005
R12339 VSS.n176 VSS.n20 4.5005
R12340 VSS.n212 VSS.n20 4.5005
R12341 VSS.n175 VSS.n20 4.5005
R12342 VSS.n213 VSS.n20 4.5005
R12343 VSS.n174 VSS.n20 4.5005
R12344 VSS.n214 VSS.n20 4.5005
R12345 VSS.n173 VSS.n20 4.5005
R12346 VSS.n215 VSS.n20 4.5005
R12347 VSS.n172 VSS.n20 4.5005
R12348 VSS.n216 VSS.n20 4.5005
R12349 VSS.n171 VSS.n20 4.5005
R12350 VSS.n217 VSS.n20 4.5005
R12351 VSS.n170 VSS.n20 4.5005
R12352 VSS.n218 VSS.n20 4.5005
R12353 VSS.n169 VSS.n20 4.5005
R12354 VSS.n219 VSS.n20 4.5005
R12355 VSS.n168 VSS.n20 4.5005
R12356 VSS.n220 VSS.n20 4.5005
R12357 VSS.n167 VSS.n20 4.5005
R12358 VSS.n221 VSS.n20 4.5005
R12359 VSS.n166 VSS.n20 4.5005
R12360 VSS.n222 VSS.n20 4.5005
R12361 VSS.n165 VSS.n20 4.5005
R12362 VSS.n223 VSS.n20 4.5005
R12363 VSS.n164 VSS.n20 4.5005
R12364 VSS.n224 VSS.n20 4.5005
R12365 VSS.n163 VSS.n20 4.5005
R12366 VSS.n225 VSS.n20 4.5005
R12367 VSS.n162 VSS.n20 4.5005
R12368 VSS.n226 VSS.n20 4.5005
R12369 VSS.n161 VSS.n20 4.5005
R12370 VSS.n227 VSS.n20 4.5005
R12371 VSS.n160 VSS.n20 4.5005
R12372 VSS.n228 VSS.n20 4.5005
R12373 VSS.n159 VSS.n20 4.5005
R12374 VSS.n229 VSS.n20 4.5005
R12375 VSS.n158 VSS.n20 4.5005
R12376 VSS.n230 VSS.n20 4.5005
R12377 VSS.n157 VSS.n20 4.5005
R12378 VSS.n231 VSS.n20 4.5005
R12379 VSS.n156 VSS.n20 4.5005
R12380 VSS.n232 VSS.n20 4.5005
R12381 VSS.n155 VSS.n20 4.5005
R12382 VSS.n233 VSS.n20 4.5005
R12383 VSS.n154 VSS.n20 4.5005
R12384 VSS.n234 VSS.n20 4.5005
R12385 VSS.n153 VSS.n20 4.5005
R12386 VSS.n235 VSS.n20 4.5005
R12387 VSS.n4506 VSS.n20 4.5005
R12388 VSS.n236 VSS.n20 4.5005
R12389 VSS.n152 VSS.n20 4.5005
R12390 VSS.n237 VSS.n20 4.5005
R12391 VSS.n151 VSS.n20 4.5005
R12392 VSS.n238 VSS.n20 4.5005
R12393 VSS.n150 VSS.n20 4.5005
R12394 VSS.n239 VSS.n20 4.5005
R12395 VSS.n149 VSS.n20 4.5005
R12396 VSS.n240 VSS.n20 4.5005
R12397 VSS.n148 VSS.n20 4.5005
R12398 VSS.n241 VSS.n20 4.5005
R12399 VSS.n147 VSS.n20 4.5005
R12400 VSS.n242 VSS.n20 4.5005
R12401 VSS.n146 VSS.n20 4.5005
R12402 VSS.n243 VSS.n20 4.5005
R12403 VSS.n145 VSS.n20 4.5005
R12404 VSS.n244 VSS.n20 4.5005
R12405 VSS.n144 VSS.n20 4.5005
R12406 VSS.n245 VSS.n20 4.5005
R12407 VSS.n143 VSS.n20 4.5005
R12408 VSS.n246 VSS.n20 4.5005
R12409 VSS.n142 VSS.n20 4.5005
R12410 VSS.n247 VSS.n20 4.5005
R12411 VSS.n141 VSS.n20 4.5005
R12412 VSS.n248 VSS.n20 4.5005
R12413 VSS.n140 VSS.n20 4.5005
R12414 VSS.n249 VSS.n20 4.5005
R12415 VSS.n139 VSS.n20 4.5005
R12416 VSS.n250 VSS.n20 4.5005
R12417 VSS.n138 VSS.n20 4.5005
R12418 VSS.n251 VSS.n20 4.5005
R12419 VSS.n137 VSS.n20 4.5005
R12420 VSS.n252 VSS.n20 4.5005
R12421 VSS.n136 VSS.n20 4.5005
R12422 VSS.n253 VSS.n20 4.5005
R12423 VSS.n135 VSS.n20 4.5005
R12424 VSS.n254 VSS.n20 4.5005
R12425 VSS.n134 VSS.n20 4.5005
R12426 VSS.n255 VSS.n20 4.5005
R12427 VSS.n133 VSS.n20 4.5005
R12428 VSS.n256 VSS.n20 4.5005
R12429 VSS.n132 VSS.n20 4.5005
R12430 VSS.n4502 VSS.n20 4.5005
R12431 VSS.n4504 VSS.n20 4.5005
R12432 VSS.n193 VSS.n117 4.5005
R12433 VSS.n195 VSS.n117 4.5005
R12434 VSS.n192 VSS.n117 4.5005
R12435 VSS.n196 VSS.n117 4.5005
R12436 VSS.n191 VSS.n117 4.5005
R12437 VSS.n197 VSS.n117 4.5005
R12438 VSS.n190 VSS.n117 4.5005
R12439 VSS.n198 VSS.n117 4.5005
R12440 VSS.n189 VSS.n117 4.5005
R12441 VSS.n199 VSS.n117 4.5005
R12442 VSS.n188 VSS.n117 4.5005
R12443 VSS.n200 VSS.n117 4.5005
R12444 VSS.n187 VSS.n117 4.5005
R12445 VSS.n201 VSS.n117 4.5005
R12446 VSS.n186 VSS.n117 4.5005
R12447 VSS.n202 VSS.n117 4.5005
R12448 VSS.n185 VSS.n117 4.5005
R12449 VSS.n203 VSS.n117 4.5005
R12450 VSS.n184 VSS.n117 4.5005
R12451 VSS.n204 VSS.n117 4.5005
R12452 VSS.n183 VSS.n117 4.5005
R12453 VSS.n205 VSS.n117 4.5005
R12454 VSS.n182 VSS.n117 4.5005
R12455 VSS.n206 VSS.n117 4.5005
R12456 VSS.n181 VSS.n117 4.5005
R12457 VSS.n207 VSS.n117 4.5005
R12458 VSS.n180 VSS.n117 4.5005
R12459 VSS.n208 VSS.n117 4.5005
R12460 VSS.n179 VSS.n117 4.5005
R12461 VSS.n209 VSS.n117 4.5005
R12462 VSS.n178 VSS.n117 4.5005
R12463 VSS.n210 VSS.n117 4.5005
R12464 VSS.n177 VSS.n117 4.5005
R12465 VSS.n211 VSS.n117 4.5005
R12466 VSS.n176 VSS.n117 4.5005
R12467 VSS.n212 VSS.n117 4.5005
R12468 VSS.n175 VSS.n117 4.5005
R12469 VSS.n213 VSS.n117 4.5005
R12470 VSS.n174 VSS.n117 4.5005
R12471 VSS.n214 VSS.n117 4.5005
R12472 VSS.n173 VSS.n117 4.5005
R12473 VSS.n215 VSS.n117 4.5005
R12474 VSS.n172 VSS.n117 4.5005
R12475 VSS.n216 VSS.n117 4.5005
R12476 VSS.n171 VSS.n117 4.5005
R12477 VSS.n217 VSS.n117 4.5005
R12478 VSS.n170 VSS.n117 4.5005
R12479 VSS.n218 VSS.n117 4.5005
R12480 VSS.n169 VSS.n117 4.5005
R12481 VSS.n219 VSS.n117 4.5005
R12482 VSS.n168 VSS.n117 4.5005
R12483 VSS.n220 VSS.n117 4.5005
R12484 VSS.n167 VSS.n117 4.5005
R12485 VSS.n221 VSS.n117 4.5005
R12486 VSS.n166 VSS.n117 4.5005
R12487 VSS.n222 VSS.n117 4.5005
R12488 VSS.n165 VSS.n117 4.5005
R12489 VSS.n223 VSS.n117 4.5005
R12490 VSS.n164 VSS.n117 4.5005
R12491 VSS.n224 VSS.n117 4.5005
R12492 VSS.n163 VSS.n117 4.5005
R12493 VSS.n225 VSS.n117 4.5005
R12494 VSS.n162 VSS.n117 4.5005
R12495 VSS.n226 VSS.n117 4.5005
R12496 VSS.n161 VSS.n117 4.5005
R12497 VSS.n227 VSS.n117 4.5005
R12498 VSS.n160 VSS.n117 4.5005
R12499 VSS.n228 VSS.n117 4.5005
R12500 VSS.n159 VSS.n117 4.5005
R12501 VSS.n229 VSS.n117 4.5005
R12502 VSS.n158 VSS.n117 4.5005
R12503 VSS.n230 VSS.n117 4.5005
R12504 VSS.n157 VSS.n117 4.5005
R12505 VSS.n231 VSS.n117 4.5005
R12506 VSS.n156 VSS.n117 4.5005
R12507 VSS.n232 VSS.n117 4.5005
R12508 VSS.n155 VSS.n117 4.5005
R12509 VSS.n233 VSS.n117 4.5005
R12510 VSS.n154 VSS.n117 4.5005
R12511 VSS.n234 VSS.n117 4.5005
R12512 VSS.n153 VSS.n117 4.5005
R12513 VSS.n235 VSS.n117 4.5005
R12514 VSS.n4506 VSS.n117 4.5005
R12515 VSS.n236 VSS.n117 4.5005
R12516 VSS.n152 VSS.n117 4.5005
R12517 VSS.n237 VSS.n117 4.5005
R12518 VSS.n151 VSS.n117 4.5005
R12519 VSS.n238 VSS.n117 4.5005
R12520 VSS.n150 VSS.n117 4.5005
R12521 VSS.n239 VSS.n117 4.5005
R12522 VSS.n149 VSS.n117 4.5005
R12523 VSS.n240 VSS.n117 4.5005
R12524 VSS.n148 VSS.n117 4.5005
R12525 VSS.n241 VSS.n117 4.5005
R12526 VSS.n147 VSS.n117 4.5005
R12527 VSS.n242 VSS.n117 4.5005
R12528 VSS.n146 VSS.n117 4.5005
R12529 VSS.n243 VSS.n117 4.5005
R12530 VSS.n145 VSS.n117 4.5005
R12531 VSS.n244 VSS.n117 4.5005
R12532 VSS.n144 VSS.n117 4.5005
R12533 VSS.n245 VSS.n117 4.5005
R12534 VSS.n143 VSS.n117 4.5005
R12535 VSS.n246 VSS.n117 4.5005
R12536 VSS.n142 VSS.n117 4.5005
R12537 VSS.n247 VSS.n117 4.5005
R12538 VSS.n141 VSS.n117 4.5005
R12539 VSS.n248 VSS.n117 4.5005
R12540 VSS.n140 VSS.n117 4.5005
R12541 VSS.n249 VSS.n117 4.5005
R12542 VSS.n139 VSS.n117 4.5005
R12543 VSS.n250 VSS.n117 4.5005
R12544 VSS.n138 VSS.n117 4.5005
R12545 VSS.n251 VSS.n117 4.5005
R12546 VSS.n137 VSS.n117 4.5005
R12547 VSS.n252 VSS.n117 4.5005
R12548 VSS.n136 VSS.n117 4.5005
R12549 VSS.n253 VSS.n117 4.5005
R12550 VSS.n135 VSS.n117 4.5005
R12551 VSS.n254 VSS.n117 4.5005
R12552 VSS.n134 VSS.n117 4.5005
R12553 VSS.n255 VSS.n117 4.5005
R12554 VSS.n133 VSS.n117 4.5005
R12555 VSS.n256 VSS.n117 4.5005
R12556 VSS.n132 VSS.n117 4.5005
R12557 VSS.n4502 VSS.n117 4.5005
R12558 VSS.n4504 VSS.n117 4.5005
R12559 VSS.n193 VSS.n19 4.5005
R12560 VSS.n195 VSS.n19 4.5005
R12561 VSS.n192 VSS.n19 4.5005
R12562 VSS.n196 VSS.n19 4.5005
R12563 VSS.n191 VSS.n19 4.5005
R12564 VSS.n197 VSS.n19 4.5005
R12565 VSS.n190 VSS.n19 4.5005
R12566 VSS.n198 VSS.n19 4.5005
R12567 VSS.n189 VSS.n19 4.5005
R12568 VSS.n199 VSS.n19 4.5005
R12569 VSS.n188 VSS.n19 4.5005
R12570 VSS.n200 VSS.n19 4.5005
R12571 VSS.n187 VSS.n19 4.5005
R12572 VSS.n201 VSS.n19 4.5005
R12573 VSS.n186 VSS.n19 4.5005
R12574 VSS.n202 VSS.n19 4.5005
R12575 VSS.n185 VSS.n19 4.5005
R12576 VSS.n203 VSS.n19 4.5005
R12577 VSS.n184 VSS.n19 4.5005
R12578 VSS.n204 VSS.n19 4.5005
R12579 VSS.n183 VSS.n19 4.5005
R12580 VSS.n205 VSS.n19 4.5005
R12581 VSS.n182 VSS.n19 4.5005
R12582 VSS.n206 VSS.n19 4.5005
R12583 VSS.n181 VSS.n19 4.5005
R12584 VSS.n207 VSS.n19 4.5005
R12585 VSS.n180 VSS.n19 4.5005
R12586 VSS.n208 VSS.n19 4.5005
R12587 VSS.n179 VSS.n19 4.5005
R12588 VSS.n209 VSS.n19 4.5005
R12589 VSS.n178 VSS.n19 4.5005
R12590 VSS.n210 VSS.n19 4.5005
R12591 VSS.n177 VSS.n19 4.5005
R12592 VSS.n211 VSS.n19 4.5005
R12593 VSS.n176 VSS.n19 4.5005
R12594 VSS.n212 VSS.n19 4.5005
R12595 VSS.n175 VSS.n19 4.5005
R12596 VSS.n213 VSS.n19 4.5005
R12597 VSS.n174 VSS.n19 4.5005
R12598 VSS.n214 VSS.n19 4.5005
R12599 VSS.n173 VSS.n19 4.5005
R12600 VSS.n215 VSS.n19 4.5005
R12601 VSS.n172 VSS.n19 4.5005
R12602 VSS.n216 VSS.n19 4.5005
R12603 VSS.n171 VSS.n19 4.5005
R12604 VSS.n217 VSS.n19 4.5005
R12605 VSS.n170 VSS.n19 4.5005
R12606 VSS.n218 VSS.n19 4.5005
R12607 VSS.n169 VSS.n19 4.5005
R12608 VSS.n219 VSS.n19 4.5005
R12609 VSS.n168 VSS.n19 4.5005
R12610 VSS.n220 VSS.n19 4.5005
R12611 VSS.n167 VSS.n19 4.5005
R12612 VSS.n221 VSS.n19 4.5005
R12613 VSS.n166 VSS.n19 4.5005
R12614 VSS.n222 VSS.n19 4.5005
R12615 VSS.n165 VSS.n19 4.5005
R12616 VSS.n223 VSS.n19 4.5005
R12617 VSS.n164 VSS.n19 4.5005
R12618 VSS.n224 VSS.n19 4.5005
R12619 VSS.n163 VSS.n19 4.5005
R12620 VSS.n225 VSS.n19 4.5005
R12621 VSS.n162 VSS.n19 4.5005
R12622 VSS.n226 VSS.n19 4.5005
R12623 VSS.n161 VSS.n19 4.5005
R12624 VSS.n227 VSS.n19 4.5005
R12625 VSS.n160 VSS.n19 4.5005
R12626 VSS.n228 VSS.n19 4.5005
R12627 VSS.n159 VSS.n19 4.5005
R12628 VSS.n229 VSS.n19 4.5005
R12629 VSS.n158 VSS.n19 4.5005
R12630 VSS.n230 VSS.n19 4.5005
R12631 VSS.n157 VSS.n19 4.5005
R12632 VSS.n231 VSS.n19 4.5005
R12633 VSS.n156 VSS.n19 4.5005
R12634 VSS.n232 VSS.n19 4.5005
R12635 VSS.n155 VSS.n19 4.5005
R12636 VSS.n233 VSS.n19 4.5005
R12637 VSS.n154 VSS.n19 4.5005
R12638 VSS.n234 VSS.n19 4.5005
R12639 VSS.n153 VSS.n19 4.5005
R12640 VSS.n235 VSS.n19 4.5005
R12641 VSS.n4506 VSS.n19 4.5005
R12642 VSS.n236 VSS.n19 4.5005
R12643 VSS.n152 VSS.n19 4.5005
R12644 VSS.n237 VSS.n19 4.5005
R12645 VSS.n151 VSS.n19 4.5005
R12646 VSS.n238 VSS.n19 4.5005
R12647 VSS.n150 VSS.n19 4.5005
R12648 VSS.n239 VSS.n19 4.5005
R12649 VSS.n149 VSS.n19 4.5005
R12650 VSS.n240 VSS.n19 4.5005
R12651 VSS.n148 VSS.n19 4.5005
R12652 VSS.n241 VSS.n19 4.5005
R12653 VSS.n147 VSS.n19 4.5005
R12654 VSS.n242 VSS.n19 4.5005
R12655 VSS.n146 VSS.n19 4.5005
R12656 VSS.n243 VSS.n19 4.5005
R12657 VSS.n145 VSS.n19 4.5005
R12658 VSS.n244 VSS.n19 4.5005
R12659 VSS.n144 VSS.n19 4.5005
R12660 VSS.n245 VSS.n19 4.5005
R12661 VSS.n143 VSS.n19 4.5005
R12662 VSS.n246 VSS.n19 4.5005
R12663 VSS.n142 VSS.n19 4.5005
R12664 VSS.n247 VSS.n19 4.5005
R12665 VSS.n141 VSS.n19 4.5005
R12666 VSS.n248 VSS.n19 4.5005
R12667 VSS.n140 VSS.n19 4.5005
R12668 VSS.n249 VSS.n19 4.5005
R12669 VSS.n139 VSS.n19 4.5005
R12670 VSS.n250 VSS.n19 4.5005
R12671 VSS.n138 VSS.n19 4.5005
R12672 VSS.n251 VSS.n19 4.5005
R12673 VSS.n137 VSS.n19 4.5005
R12674 VSS.n252 VSS.n19 4.5005
R12675 VSS.n136 VSS.n19 4.5005
R12676 VSS.n253 VSS.n19 4.5005
R12677 VSS.n135 VSS.n19 4.5005
R12678 VSS.n254 VSS.n19 4.5005
R12679 VSS.n134 VSS.n19 4.5005
R12680 VSS.n255 VSS.n19 4.5005
R12681 VSS.n133 VSS.n19 4.5005
R12682 VSS.n256 VSS.n19 4.5005
R12683 VSS.n132 VSS.n19 4.5005
R12684 VSS.n4502 VSS.n19 4.5005
R12685 VSS.n4504 VSS.n19 4.5005
R12686 VSS.n193 VSS.n118 4.5005
R12687 VSS.n195 VSS.n118 4.5005
R12688 VSS.n192 VSS.n118 4.5005
R12689 VSS.n196 VSS.n118 4.5005
R12690 VSS.n191 VSS.n118 4.5005
R12691 VSS.n197 VSS.n118 4.5005
R12692 VSS.n190 VSS.n118 4.5005
R12693 VSS.n198 VSS.n118 4.5005
R12694 VSS.n189 VSS.n118 4.5005
R12695 VSS.n199 VSS.n118 4.5005
R12696 VSS.n188 VSS.n118 4.5005
R12697 VSS.n200 VSS.n118 4.5005
R12698 VSS.n187 VSS.n118 4.5005
R12699 VSS.n201 VSS.n118 4.5005
R12700 VSS.n186 VSS.n118 4.5005
R12701 VSS.n202 VSS.n118 4.5005
R12702 VSS.n185 VSS.n118 4.5005
R12703 VSS.n203 VSS.n118 4.5005
R12704 VSS.n184 VSS.n118 4.5005
R12705 VSS.n204 VSS.n118 4.5005
R12706 VSS.n183 VSS.n118 4.5005
R12707 VSS.n205 VSS.n118 4.5005
R12708 VSS.n182 VSS.n118 4.5005
R12709 VSS.n206 VSS.n118 4.5005
R12710 VSS.n181 VSS.n118 4.5005
R12711 VSS.n207 VSS.n118 4.5005
R12712 VSS.n180 VSS.n118 4.5005
R12713 VSS.n208 VSS.n118 4.5005
R12714 VSS.n179 VSS.n118 4.5005
R12715 VSS.n209 VSS.n118 4.5005
R12716 VSS.n178 VSS.n118 4.5005
R12717 VSS.n210 VSS.n118 4.5005
R12718 VSS.n177 VSS.n118 4.5005
R12719 VSS.n211 VSS.n118 4.5005
R12720 VSS.n176 VSS.n118 4.5005
R12721 VSS.n212 VSS.n118 4.5005
R12722 VSS.n175 VSS.n118 4.5005
R12723 VSS.n213 VSS.n118 4.5005
R12724 VSS.n174 VSS.n118 4.5005
R12725 VSS.n214 VSS.n118 4.5005
R12726 VSS.n173 VSS.n118 4.5005
R12727 VSS.n215 VSS.n118 4.5005
R12728 VSS.n172 VSS.n118 4.5005
R12729 VSS.n216 VSS.n118 4.5005
R12730 VSS.n171 VSS.n118 4.5005
R12731 VSS.n217 VSS.n118 4.5005
R12732 VSS.n170 VSS.n118 4.5005
R12733 VSS.n218 VSS.n118 4.5005
R12734 VSS.n169 VSS.n118 4.5005
R12735 VSS.n219 VSS.n118 4.5005
R12736 VSS.n168 VSS.n118 4.5005
R12737 VSS.n220 VSS.n118 4.5005
R12738 VSS.n167 VSS.n118 4.5005
R12739 VSS.n221 VSS.n118 4.5005
R12740 VSS.n166 VSS.n118 4.5005
R12741 VSS.n222 VSS.n118 4.5005
R12742 VSS.n165 VSS.n118 4.5005
R12743 VSS.n223 VSS.n118 4.5005
R12744 VSS.n164 VSS.n118 4.5005
R12745 VSS.n224 VSS.n118 4.5005
R12746 VSS.n163 VSS.n118 4.5005
R12747 VSS.n225 VSS.n118 4.5005
R12748 VSS.n162 VSS.n118 4.5005
R12749 VSS.n226 VSS.n118 4.5005
R12750 VSS.n161 VSS.n118 4.5005
R12751 VSS.n227 VSS.n118 4.5005
R12752 VSS.n160 VSS.n118 4.5005
R12753 VSS.n228 VSS.n118 4.5005
R12754 VSS.n159 VSS.n118 4.5005
R12755 VSS.n229 VSS.n118 4.5005
R12756 VSS.n158 VSS.n118 4.5005
R12757 VSS.n230 VSS.n118 4.5005
R12758 VSS.n157 VSS.n118 4.5005
R12759 VSS.n231 VSS.n118 4.5005
R12760 VSS.n156 VSS.n118 4.5005
R12761 VSS.n232 VSS.n118 4.5005
R12762 VSS.n155 VSS.n118 4.5005
R12763 VSS.n233 VSS.n118 4.5005
R12764 VSS.n154 VSS.n118 4.5005
R12765 VSS.n234 VSS.n118 4.5005
R12766 VSS.n153 VSS.n118 4.5005
R12767 VSS.n235 VSS.n118 4.5005
R12768 VSS.n4506 VSS.n118 4.5005
R12769 VSS.n236 VSS.n118 4.5005
R12770 VSS.n152 VSS.n118 4.5005
R12771 VSS.n237 VSS.n118 4.5005
R12772 VSS.n151 VSS.n118 4.5005
R12773 VSS.n238 VSS.n118 4.5005
R12774 VSS.n150 VSS.n118 4.5005
R12775 VSS.n239 VSS.n118 4.5005
R12776 VSS.n149 VSS.n118 4.5005
R12777 VSS.n240 VSS.n118 4.5005
R12778 VSS.n148 VSS.n118 4.5005
R12779 VSS.n241 VSS.n118 4.5005
R12780 VSS.n147 VSS.n118 4.5005
R12781 VSS.n242 VSS.n118 4.5005
R12782 VSS.n146 VSS.n118 4.5005
R12783 VSS.n243 VSS.n118 4.5005
R12784 VSS.n145 VSS.n118 4.5005
R12785 VSS.n244 VSS.n118 4.5005
R12786 VSS.n144 VSS.n118 4.5005
R12787 VSS.n245 VSS.n118 4.5005
R12788 VSS.n143 VSS.n118 4.5005
R12789 VSS.n246 VSS.n118 4.5005
R12790 VSS.n142 VSS.n118 4.5005
R12791 VSS.n247 VSS.n118 4.5005
R12792 VSS.n141 VSS.n118 4.5005
R12793 VSS.n248 VSS.n118 4.5005
R12794 VSS.n140 VSS.n118 4.5005
R12795 VSS.n249 VSS.n118 4.5005
R12796 VSS.n139 VSS.n118 4.5005
R12797 VSS.n250 VSS.n118 4.5005
R12798 VSS.n138 VSS.n118 4.5005
R12799 VSS.n251 VSS.n118 4.5005
R12800 VSS.n137 VSS.n118 4.5005
R12801 VSS.n252 VSS.n118 4.5005
R12802 VSS.n136 VSS.n118 4.5005
R12803 VSS.n253 VSS.n118 4.5005
R12804 VSS.n135 VSS.n118 4.5005
R12805 VSS.n254 VSS.n118 4.5005
R12806 VSS.n134 VSS.n118 4.5005
R12807 VSS.n255 VSS.n118 4.5005
R12808 VSS.n133 VSS.n118 4.5005
R12809 VSS.n256 VSS.n118 4.5005
R12810 VSS.n132 VSS.n118 4.5005
R12811 VSS.n4502 VSS.n118 4.5005
R12812 VSS.n4504 VSS.n118 4.5005
R12813 VSS.n193 VSS.n18 4.5005
R12814 VSS.n195 VSS.n18 4.5005
R12815 VSS.n192 VSS.n18 4.5005
R12816 VSS.n196 VSS.n18 4.5005
R12817 VSS.n191 VSS.n18 4.5005
R12818 VSS.n197 VSS.n18 4.5005
R12819 VSS.n190 VSS.n18 4.5005
R12820 VSS.n198 VSS.n18 4.5005
R12821 VSS.n189 VSS.n18 4.5005
R12822 VSS.n199 VSS.n18 4.5005
R12823 VSS.n188 VSS.n18 4.5005
R12824 VSS.n200 VSS.n18 4.5005
R12825 VSS.n187 VSS.n18 4.5005
R12826 VSS.n201 VSS.n18 4.5005
R12827 VSS.n186 VSS.n18 4.5005
R12828 VSS.n202 VSS.n18 4.5005
R12829 VSS.n185 VSS.n18 4.5005
R12830 VSS.n203 VSS.n18 4.5005
R12831 VSS.n184 VSS.n18 4.5005
R12832 VSS.n204 VSS.n18 4.5005
R12833 VSS.n183 VSS.n18 4.5005
R12834 VSS.n205 VSS.n18 4.5005
R12835 VSS.n182 VSS.n18 4.5005
R12836 VSS.n206 VSS.n18 4.5005
R12837 VSS.n181 VSS.n18 4.5005
R12838 VSS.n207 VSS.n18 4.5005
R12839 VSS.n180 VSS.n18 4.5005
R12840 VSS.n208 VSS.n18 4.5005
R12841 VSS.n179 VSS.n18 4.5005
R12842 VSS.n209 VSS.n18 4.5005
R12843 VSS.n178 VSS.n18 4.5005
R12844 VSS.n210 VSS.n18 4.5005
R12845 VSS.n177 VSS.n18 4.5005
R12846 VSS.n211 VSS.n18 4.5005
R12847 VSS.n176 VSS.n18 4.5005
R12848 VSS.n212 VSS.n18 4.5005
R12849 VSS.n175 VSS.n18 4.5005
R12850 VSS.n213 VSS.n18 4.5005
R12851 VSS.n174 VSS.n18 4.5005
R12852 VSS.n214 VSS.n18 4.5005
R12853 VSS.n173 VSS.n18 4.5005
R12854 VSS.n215 VSS.n18 4.5005
R12855 VSS.n172 VSS.n18 4.5005
R12856 VSS.n216 VSS.n18 4.5005
R12857 VSS.n171 VSS.n18 4.5005
R12858 VSS.n217 VSS.n18 4.5005
R12859 VSS.n170 VSS.n18 4.5005
R12860 VSS.n218 VSS.n18 4.5005
R12861 VSS.n169 VSS.n18 4.5005
R12862 VSS.n219 VSS.n18 4.5005
R12863 VSS.n168 VSS.n18 4.5005
R12864 VSS.n220 VSS.n18 4.5005
R12865 VSS.n167 VSS.n18 4.5005
R12866 VSS.n221 VSS.n18 4.5005
R12867 VSS.n166 VSS.n18 4.5005
R12868 VSS.n222 VSS.n18 4.5005
R12869 VSS.n165 VSS.n18 4.5005
R12870 VSS.n223 VSS.n18 4.5005
R12871 VSS.n164 VSS.n18 4.5005
R12872 VSS.n224 VSS.n18 4.5005
R12873 VSS.n163 VSS.n18 4.5005
R12874 VSS.n225 VSS.n18 4.5005
R12875 VSS.n162 VSS.n18 4.5005
R12876 VSS.n226 VSS.n18 4.5005
R12877 VSS.n161 VSS.n18 4.5005
R12878 VSS.n227 VSS.n18 4.5005
R12879 VSS.n160 VSS.n18 4.5005
R12880 VSS.n228 VSS.n18 4.5005
R12881 VSS.n159 VSS.n18 4.5005
R12882 VSS.n229 VSS.n18 4.5005
R12883 VSS.n158 VSS.n18 4.5005
R12884 VSS.n230 VSS.n18 4.5005
R12885 VSS.n157 VSS.n18 4.5005
R12886 VSS.n231 VSS.n18 4.5005
R12887 VSS.n156 VSS.n18 4.5005
R12888 VSS.n232 VSS.n18 4.5005
R12889 VSS.n155 VSS.n18 4.5005
R12890 VSS.n233 VSS.n18 4.5005
R12891 VSS.n154 VSS.n18 4.5005
R12892 VSS.n234 VSS.n18 4.5005
R12893 VSS.n153 VSS.n18 4.5005
R12894 VSS.n235 VSS.n18 4.5005
R12895 VSS.n4506 VSS.n18 4.5005
R12896 VSS.n236 VSS.n18 4.5005
R12897 VSS.n152 VSS.n18 4.5005
R12898 VSS.n237 VSS.n18 4.5005
R12899 VSS.n151 VSS.n18 4.5005
R12900 VSS.n238 VSS.n18 4.5005
R12901 VSS.n150 VSS.n18 4.5005
R12902 VSS.n239 VSS.n18 4.5005
R12903 VSS.n149 VSS.n18 4.5005
R12904 VSS.n240 VSS.n18 4.5005
R12905 VSS.n148 VSS.n18 4.5005
R12906 VSS.n241 VSS.n18 4.5005
R12907 VSS.n147 VSS.n18 4.5005
R12908 VSS.n242 VSS.n18 4.5005
R12909 VSS.n146 VSS.n18 4.5005
R12910 VSS.n243 VSS.n18 4.5005
R12911 VSS.n145 VSS.n18 4.5005
R12912 VSS.n244 VSS.n18 4.5005
R12913 VSS.n144 VSS.n18 4.5005
R12914 VSS.n245 VSS.n18 4.5005
R12915 VSS.n143 VSS.n18 4.5005
R12916 VSS.n246 VSS.n18 4.5005
R12917 VSS.n142 VSS.n18 4.5005
R12918 VSS.n247 VSS.n18 4.5005
R12919 VSS.n141 VSS.n18 4.5005
R12920 VSS.n248 VSS.n18 4.5005
R12921 VSS.n140 VSS.n18 4.5005
R12922 VSS.n249 VSS.n18 4.5005
R12923 VSS.n139 VSS.n18 4.5005
R12924 VSS.n250 VSS.n18 4.5005
R12925 VSS.n138 VSS.n18 4.5005
R12926 VSS.n251 VSS.n18 4.5005
R12927 VSS.n137 VSS.n18 4.5005
R12928 VSS.n252 VSS.n18 4.5005
R12929 VSS.n136 VSS.n18 4.5005
R12930 VSS.n253 VSS.n18 4.5005
R12931 VSS.n135 VSS.n18 4.5005
R12932 VSS.n254 VSS.n18 4.5005
R12933 VSS.n134 VSS.n18 4.5005
R12934 VSS.n255 VSS.n18 4.5005
R12935 VSS.n133 VSS.n18 4.5005
R12936 VSS.n256 VSS.n18 4.5005
R12937 VSS.n132 VSS.n18 4.5005
R12938 VSS.n4502 VSS.n18 4.5005
R12939 VSS.n4504 VSS.n18 4.5005
R12940 VSS.n193 VSS.n119 4.5005
R12941 VSS.n195 VSS.n119 4.5005
R12942 VSS.n192 VSS.n119 4.5005
R12943 VSS.n196 VSS.n119 4.5005
R12944 VSS.n191 VSS.n119 4.5005
R12945 VSS.n197 VSS.n119 4.5005
R12946 VSS.n190 VSS.n119 4.5005
R12947 VSS.n198 VSS.n119 4.5005
R12948 VSS.n189 VSS.n119 4.5005
R12949 VSS.n199 VSS.n119 4.5005
R12950 VSS.n188 VSS.n119 4.5005
R12951 VSS.n200 VSS.n119 4.5005
R12952 VSS.n187 VSS.n119 4.5005
R12953 VSS.n201 VSS.n119 4.5005
R12954 VSS.n186 VSS.n119 4.5005
R12955 VSS.n202 VSS.n119 4.5005
R12956 VSS.n185 VSS.n119 4.5005
R12957 VSS.n203 VSS.n119 4.5005
R12958 VSS.n184 VSS.n119 4.5005
R12959 VSS.n204 VSS.n119 4.5005
R12960 VSS.n183 VSS.n119 4.5005
R12961 VSS.n205 VSS.n119 4.5005
R12962 VSS.n182 VSS.n119 4.5005
R12963 VSS.n206 VSS.n119 4.5005
R12964 VSS.n181 VSS.n119 4.5005
R12965 VSS.n207 VSS.n119 4.5005
R12966 VSS.n180 VSS.n119 4.5005
R12967 VSS.n208 VSS.n119 4.5005
R12968 VSS.n179 VSS.n119 4.5005
R12969 VSS.n209 VSS.n119 4.5005
R12970 VSS.n178 VSS.n119 4.5005
R12971 VSS.n210 VSS.n119 4.5005
R12972 VSS.n177 VSS.n119 4.5005
R12973 VSS.n211 VSS.n119 4.5005
R12974 VSS.n176 VSS.n119 4.5005
R12975 VSS.n212 VSS.n119 4.5005
R12976 VSS.n175 VSS.n119 4.5005
R12977 VSS.n213 VSS.n119 4.5005
R12978 VSS.n174 VSS.n119 4.5005
R12979 VSS.n214 VSS.n119 4.5005
R12980 VSS.n173 VSS.n119 4.5005
R12981 VSS.n215 VSS.n119 4.5005
R12982 VSS.n172 VSS.n119 4.5005
R12983 VSS.n216 VSS.n119 4.5005
R12984 VSS.n171 VSS.n119 4.5005
R12985 VSS.n217 VSS.n119 4.5005
R12986 VSS.n170 VSS.n119 4.5005
R12987 VSS.n218 VSS.n119 4.5005
R12988 VSS.n169 VSS.n119 4.5005
R12989 VSS.n219 VSS.n119 4.5005
R12990 VSS.n168 VSS.n119 4.5005
R12991 VSS.n220 VSS.n119 4.5005
R12992 VSS.n167 VSS.n119 4.5005
R12993 VSS.n221 VSS.n119 4.5005
R12994 VSS.n166 VSS.n119 4.5005
R12995 VSS.n222 VSS.n119 4.5005
R12996 VSS.n165 VSS.n119 4.5005
R12997 VSS.n223 VSS.n119 4.5005
R12998 VSS.n164 VSS.n119 4.5005
R12999 VSS.n224 VSS.n119 4.5005
R13000 VSS.n163 VSS.n119 4.5005
R13001 VSS.n225 VSS.n119 4.5005
R13002 VSS.n162 VSS.n119 4.5005
R13003 VSS.n226 VSS.n119 4.5005
R13004 VSS.n161 VSS.n119 4.5005
R13005 VSS.n227 VSS.n119 4.5005
R13006 VSS.n160 VSS.n119 4.5005
R13007 VSS.n228 VSS.n119 4.5005
R13008 VSS.n159 VSS.n119 4.5005
R13009 VSS.n229 VSS.n119 4.5005
R13010 VSS.n158 VSS.n119 4.5005
R13011 VSS.n230 VSS.n119 4.5005
R13012 VSS.n157 VSS.n119 4.5005
R13013 VSS.n231 VSS.n119 4.5005
R13014 VSS.n156 VSS.n119 4.5005
R13015 VSS.n232 VSS.n119 4.5005
R13016 VSS.n155 VSS.n119 4.5005
R13017 VSS.n233 VSS.n119 4.5005
R13018 VSS.n154 VSS.n119 4.5005
R13019 VSS.n234 VSS.n119 4.5005
R13020 VSS.n153 VSS.n119 4.5005
R13021 VSS.n235 VSS.n119 4.5005
R13022 VSS.n4506 VSS.n119 4.5005
R13023 VSS.n236 VSS.n119 4.5005
R13024 VSS.n152 VSS.n119 4.5005
R13025 VSS.n237 VSS.n119 4.5005
R13026 VSS.n151 VSS.n119 4.5005
R13027 VSS.n238 VSS.n119 4.5005
R13028 VSS.n150 VSS.n119 4.5005
R13029 VSS.n239 VSS.n119 4.5005
R13030 VSS.n149 VSS.n119 4.5005
R13031 VSS.n240 VSS.n119 4.5005
R13032 VSS.n148 VSS.n119 4.5005
R13033 VSS.n241 VSS.n119 4.5005
R13034 VSS.n147 VSS.n119 4.5005
R13035 VSS.n242 VSS.n119 4.5005
R13036 VSS.n146 VSS.n119 4.5005
R13037 VSS.n243 VSS.n119 4.5005
R13038 VSS.n145 VSS.n119 4.5005
R13039 VSS.n244 VSS.n119 4.5005
R13040 VSS.n144 VSS.n119 4.5005
R13041 VSS.n245 VSS.n119 4.5005
R13042 VSS.n143 VSS.n119 4.5005
R13043 VSS.n246 VSS.n119 4.5005
R13044 VSS.n142 VSS.n119 4.5005
R13045 VSS.n247 VSS.n119 4.5005
R13046 VSS.n141 VSS.n119 4.5005
R13047 VSS.n248 VSS.n119 4.5005
R13048 VSS.n140 VSS.n119 4.5005
R13049 VSS.n249 VSS.n119 4.5005
R13050 VSS.n139 VSS.n119 4.5005
R13051 VSS.n250 VSS.n119 4.5005
R13052 VSS.n138 VSS.n119 4.5005
R13053 VSS.n251 VSS.n119 4.5005
R13054 VSS.n137 VSS.n119 4.5005
R13055 VSS.n252 VSS.n119 4.5005
R13056 VSS.n136 VSS.n119 4.5005
R13057 VSS.n253 VSS.n119 4.5005
R13058 VSS.n135 VSS.n119 4.5005
R13059 VSS.n254 VSS.n119 4.5005
R13060 VSS.n134 VSS.n119 4.5005
R13061 VSS.n255 VSS.n119 4.5005
R13062 VSS.n133 VSS.n119 4.5005
R13063 VSS.n256 VSS.n119 4.5005
R13064 VSS.n132 VSS.n119 4.5005
R13065 VSS.n4502 VSS.n119 4.5005
R13066 VSS.n4504 VSS.n119 4.5005
R13067 VSS.n193 VSS.n17 4.5005
R13068 VSS.n195 VSS.n17 4.5005
R13069 VSS.n192 VSS.n17 4.5005
R13070 VSS.n196 VSS.n17 4.5005
R13071 VSS.n191 VSS.n17 4.5005
R13072 VSS.n197 VSS.n17 4.5005
R13073 VSS.n190 VSS.n17 4.5005
R13074 VSS.n198 VSS.n17 4.5005
R13075 VSS.n189 VSS.n17 4.5005
R13076 VSS.n199 VSS.n17 4.5005
R13077 VSS.n188 VSS.n17 4.5005
R13078 VSS.n200 VSS.n17 4.5005
R13079 VSS.n187 VSS.n17 4.5005
R13080 VSS.n201 VSS.n17 4.5005
R13081 VSS.n186 VSS.n17 4.5005
R13082 VSS.n202 VSS.n17 4.5005
R13083 VSS.n185 VSS.n17 4.5005
R13084 VSS.n203 VSS.n17 4.5005
R13085 VSS.n184 VSS.n17 4.5005
R13086 VSS.n204 VSS.n17 4.5005
R13087 VSS.n183 VSS.n17 4.5005
R13088 VSS.n205 VSS.n17 4.5005
R13089 VSS.n182 VSS.n17 4.5005
R13090 VSS.n206 VSS.n17 4.5005
R13091 VSS.n181 VSS.n17 4.5005
R13092 VSS.n207 VSS.n17 4.5005
R13093 VSS.n180 VSS.n17 4.5005
R13094 VSS.n208 VSS.n17 4.5005
R13095 VSS.n179 VSS.n17 4.5005
R13096 VSS.n209 VSS.n17 4.5005
R13097 VSS.n178 VSS.n17 4.5005
R13098 VSS.n210 VSS.n17 4.5005
R13099 VSS.n177 VSS.n17 4.5005
R13100 VSS.n211 VSS.n17 4.5005
R13101 VSS.n176 VSS.n17 4.5005
R13102 VSS.n212 VSS.n17 4.5005
R13103 VSS.n175 VSS.n17 4.5005
R13104 VSS.n213 VSS.n17 4.5005
R13105 VSS.n174 VSS.n17 4.5005
R13106 VSS.n214 VSS.n17 4.5005
R13107 VSS.n173 VSS.n17 4.5005
R13108 VSS.n215 VSS.n17 4.5005
R13109 VSS.n172 VSS.n17 4.5005
R13110 VSS.n216 VSS.n17 4.5005
R13111 VSS.n171 VSS.n17 4.5005
R13112 VSS.n217 VSS.n17 4.5005
R13113 VSS.n170 VSS.n17 4.5005
R13114 VSS.n218 VSS.n17 4.5005
R13115 VSS.n169 VSS.n17 4.5005
R13116 VSS.n219 VSS.n17 4.5005
R13117 VSS.n168 VSS.n17 4.5005
R13118 VSS.n220 VSS.n17 4.5005
R13119 VSS.n167 VSS.n17 4.5005
R13120 VSS.n221 VSS.n17 4.5005
R13121 VSS.n166 VSS.n17 4.5005
R13122 VSS.n222 VSS.n17 4.5005
R13123 VSS.n165 VSS.n17 4.5005
R13124 VSS.n223 VSS.n17 4.5005
R13125 VSS.n164 VSS.n17 4.5005
R13126 VSS.n224 VSS.n17 4.5005
R13127 VSS.n163 VSS.n17 4.5005
R13128 VSS.n225 VSS.n17 4.5005
R13129 VSS.n162 VSS.n17 4.5005
R13130 VSS.n226 VSS.n17 4.5005
R13131 VSS.n161 VSS.n17 4.5005
R13132 VSS.n227 VSS.n17 4.5005
R13133 VSS.n160 VSS.n17 4.5005
R13134 VSS.n228 VSS.n17 4.5005
R13135 VSS.n159 VSS.n17 4.5005
R13136 VSS.n229 VSS.n17 4.5005
R13137 VSS.n158 VSS.n17 4.5005
R13138 VSS.n230 VSS.n17 4.5005
R13139 VSS.n157 VSS.n17 4.5005
R13140 VSS.n231 VSS.n17 4.5005
R13141 VSS.n156 VSS.n17 4.5005
R13142 VSS.n232 VSS.n17 4.5005
R13143 VSS.n155 VSS.n17 4.5005
R13144 VSS.n233 VSS.n17 4.5005
R13145 VSS.n154 VSS.n17 4.5005
R13146 VSS.n234 VSS.n17 4.5005
R13147 VSS.n153 VSS.n17 4.5005
R13148 VSS.n235 VSS.n17 4.5005
R13149 VSS.n4506 VSS.n17 4.5005
R13150 VSS.n236 VSS.n17 4.5005
R13151 VSS.n152 VSS.n17 4.5005
R13152 VSS.n237 VSS.n17 4.5005
R13153 VSS.n151 VSS.n17 4.5005
R13154 VSS.n238 VSS.n17 4.5005
R13155 VSS.n150 VSS.n17 4.5005
R13156 VSS.n239 VSS.n17 4.5005
R13157 VSS.n149 VSS.n17 4.5005
R13158 VSS.n240 VSS.n17 4.5005
R13159 VSS.n148 VSS.n17 4.5005
R13160 VSS.n241 VSS.n17 4.5005
R13161 VSS.n147 VSS.n17 4.5005
R13162 VSS.n242 VSS.n17 4.5005
R13163 VSS.n146 VSS.n17 4.5005
R13164 VSS.n243 VSS.n17 4.5005
R13165 VSS.n145 VSS.n17 4.5005
R13166 VSS.n244 VSS.n17 4.5005
R13167 VSS.n144 VSS.n17 4.5005
R13168 VSS.n245 VSS.n17 4.5005
R13169 VSS.n143 VSS.n17 4.5005
R13170 VSS.n246 VSS.n17 4.5005
R13171 VSS.n142 VSS.n17 4.5005
R13172 VSS.n247 VSS.n17 4.5005
R13173 VSS.n141 VSS.n17 4.5005
R13174 VSS.n248 VSS.n17 4.5005
R13175 VSS.n140 VSS.n17 4.5005
R13176 VSS.n249 VSS.n17 4.5005
R13177 VSS.n139 VSS.n17 4.5005
R13178 VSS.n250 VSS.n17 4.5005
R13179 VSS.n138 VSS.n17 4.5005
R13180 VSS.n251 VSS.n17 4.5005
R13181 VSS.n137 VSS.n17 4.5005
R13182 VSS.n252 VSS.n17 4.5005
R13183 VSS.n136 VSS.n17 4.5005
R13184 VSS.n253 VSS.n17 4.5005
R13185 VSS.n135 VSS.n17 4.5005
R13186 VSS.n254 VSS.n17 4.5005
R13187 VSS.n134 VSS.n17 4.5005
R13188 VSS.n255 VSS.n17 4.5005
R13189 VSS.n133 VSS.n17 4.5005
R13190 VSS.n256 VSS.n17 4.5005
R13191 VSS.n132 VSS.n17 4.5005
R13192 VSS.n4502 VSS.n17 4.5005
R13193 VSS.n4504 VSS.n17 4.5005
R13194 VSS.n193 VSS.n120 4.5005
R13195 VSS.n195 VSS.n120 4.5005
R13196 VSS.n192 VSS.n120 4.5005
R13197 VSS.n196 VSS.n120 4.5005
R13198 VSS.n191 VSS.n120 4.5005
R13199 VSS.n197 VSS.n120 4.5005
R13200 VSS.n190 VSS.n120 4.5005
R13201 VSS.n198 VSS.n120 4.5005
R13202 VSS.n189 VSS.n120 4.5005
R13203 VSS.n199 VSS.n120 4.5005
R13204 VSS.n188 VSS.n120 4.5005
R13205 VSS.n200 VSS.n120 4.5005
R13206 VSS.n187 VSS.n120 4.5005
R13207 VSS.n201 VSS.n120 4.5005
R13208 VSS.n186 VSS.n120 4.5005
R13209 VSS.n202 VSS.n120 4.5005
R13210 VSS.n185 VSS.n120 4.5005
R13211 VSS.n203 VSS.n120 4.5005
R13212 VSS.n184 VSS.n120 4.5005
R13213 VSS.n204 VSS.n120 4.5005
R13214 VSS.n183 VSS.n120 4.5005
R13215 VSS.n205 VSS.n120 4.5005
R13216 VSS.n182 VSS.n120 4.5005
R13217 VSS.n206 VSS.n120 4.5005
R13218 VSS.n181 VSS.n120 4.5005
R13219 VSS.n207 VSS.n120 4.5005
R13220 VSS.n180 VSS.n120 4.5005
R13221 VSS.n208 VSS.n120 4.5005
R13222 VSS.n179 VSS.n120 4.5005
R13223 VSS.n209 VSS.n120 4.5005
R13224 VSS.n178 VSS.n120 4.5005
R13225 VSS.n210 VSS.n120 4.5005
R13226 VSS.n177 VSS.n120 4.5005
R13227 VSS.n211 VSS.n120 4.5005
R13228 VSS.n176 VSS.n120 4.5005
R13229 VSS.n212 VSS.n120 4.5005
R13230 VSS.n175 VSS.n120 4.5005
R13231 VSS.n213 VSS.n120 4.5005
R13232 VSS.n174 VSS.n120 4.5005
R13233 VSS.n214 VSS.n120 4.5005
R13234 VSS.n173 VSS.n120 4.5005
R13235 VSS.n215 VSS.n120 4.5005
R13236 VSS.n172 VSS.n120 4.5005
R13237 VSS.n216 VSS.n120 4.5005
R13238 VSS.n171 VSS.n120 4.5005
R13239 VSS.n217 VSS.n120 4.5005
R13240 VSS.n170 VSS.n120 4.5005
R13241 VSS.n218 VSS.n120 4.5005
R13242 VSS.n169 VSS.n120 4.5005
R13243 VSS.n219 VSS.n120 4.5005
R13244 VSS.n168 VSS.n120 4.5005
R13245 VSS.n220 VSS.n120 4.5005
R13246 VSS.n167 VSS.n120 4.5005
R13247 VSS.n221 VSS.n120 4.5005
R13248 VSS.n166 VSS.n120 4.5005
R13249 VSS.n222 VSS.n120 4.5005
R13250 VSS.n165 VSS.n120 4.5005
R13251 VSS.n223 VSS.n120 4.5005
R13252 VSS.n164 VSS.n120 4.5005
R13253 VSS.n224 VSS.n120 4.5005
R13254 VSS.n163 VSS.n120 4.5005
R13255 VSS.n225 VSS.n120 4.5005
R13256 VSS.n162 VSS.n120 4.5005
R13257 VSS.n226 VSS.n120 4.5005
R13258 VSS.n161 VSS.n120 4.5005
R13259 VSS.n227 VSS.n120 4.5005
R13260 VSS.n160 VSS.n120 4.5005
R13261 VSS.n228 VSS.n120 4.5005
R13262 VSS.n159 VSS.n120 4.5005
R13263 VSS.n229 VSS.n120 4.5005
R13264 VSS.n158 VSS.n120 4.5005
R13265 VSS.n230 VSS.n120 4.5005
R13266 VSS.n157 VSS.n120 4.5005
R13267 VSS.n231 VSS.n120 4.5005
R13268 VSS.n156 VSS.n120 4.5005
R13269 VSS.n232 VSS.n120 4.5005
R13270 VSS.n155 VSS.n120 4.5005
R13271 VSS.n233 VSS.n120 4.5005
R13272 VSS.n154 VSS.n120 4.5005
R13273 VSS.n234 VSS.n120 4.5005
R13274 VSS.n153 VSS.n120 4.5005
R13275 VSS.n235 VSS.n120 4.5005
R13276 VSS.n4506 VSS.n120 4.5005
R13277 VSS.n236 VSS.n120 4.5005
R13278 VSS.n152 VSS.n120 4.5005
R13279 VSS.n237 VSS.n120 4.5005
R13280 VSS.n151 VSS.n120 4.5005
R13281 VSS.n238 VSS.n120 4.5005
R13282 VSS.n150 VSS.n120 4.5005
R13283 VSS.n239 VSS.n120 4.5005
R13284 VSS.n149 VSS.n120 4.5005
R13285 VSS.n240 VSS.n120 4.5005
R13286 VSS.n148 VSS.n120 4.5005
R13287 VSS.n241 VSS.n120 4.5005
R13288 VSS.n147 VSS.n120 4.5005
R13289 VSS.n242 VSS.n120 4.5005
R13290 VSS.n146 VSS.n120 4.5005
R13291 VSS.n243 VSS.n120 4.5005
R13292 VSS.n145 VSS.n120 4.5005
R13293 VSS.n244 VSS.n120 4.5005
R13294 VSS.n144 VSS.n120 4.5005
R13295 VSS.n245 VSS.n120 4.5005
R13296 VSS.n143 VSS.n120 4.5005
R13297 VSS.n246 VSS.n120 4.5005
R13298 VSS.n142 VSS.n120 4.5005
R13299 VSS.n247 VSS.n120 4.5005
R13300 VSS.n141 VSS.n120 4.5005
R13301 VSS.n248 VSS.n120 4.5005
R13302 VSS.n140 VSS.n120 4.5005
R13303 VSS.n249 VSS.n120 4.5005
R13304 VSS.n139 VSS.n120 4.5005
R13305 VSS.n250 VSS.n120 4.5005
R13306 VSS.n138 VSS.n120 4.5005
R13307 VSS.n251 VSS.n120 4.5005
R13308 VSS.n137 VSS.n120 4.5005
R13309 VSS.n252 VSS.n120 4.5005
R13310 VSS.n136 VSS.n120 4.5005
R13311 VSS.n253 VSS.n120 4.5005
R13312 VSS.n135 VSS.n120 4.5005
R13313 VSS.n254 VSS.n120 4.5005
R13314 VSS.n134 VSS.n120 4.5005
R13315 VSS.n255 VSS.n120 4.5005
R13316 VSS.n133 VSS.n120 4.5005
R13317 VSS.n256 VSS.n120 4.5005
R13318 VSS.n132 VSS.n120 4.5005
R13319 VSS.n4502 VSS.n120 4.5005
R13320 VSS.n4504 VSS.n120 4.5005
R13321 VSS.n193 VSS.n16 4.5005
R13322 VSS.n195 VSS.n16 4.5005
R13323 VSS.n192 VSS.n16 4.5005
R13324 VSS.n196 VSS.n16 4.5005
R13325 VSS.n191 VSS.n16 4.5005
R13326 VSS.n197 VSS.n16 4.5005
R13327 VSS.n190 VSS.n16 4.5005
R13328 VSS.n198 VSS.n16 4.5005
R13329 VSS.n189 VSS.n16 4.5005
R13330 VSS.n199 VSS.n16 4.5005
R13331 VSS.n188 VSS.n16 4.5005
R13332 VSS.n200 VSS.n16 4.5005
R13333 VSS.n187 VSS.n16 4.5005
R13334 VSS.n201 VSS.n16 4.5005
R13335 VSS.n186 VSS.n16 4.5005
R13336 VSS.n202 VSS.n16 4.5005
R13337 VSS.n185 VSS.n16 4.5005
R13338 VSS.n203 VSS.n16 4.5005
R13339 VSS.n184 VSS.n16 4.5005
R13340 VSS.n204 VSS.n16 4.5005
R13341 VSS.n183 VSS.n16 4.5005
R13342 VSS.n205 VSS.n16 4.5005
R13343 VSS.n182 VSS.n16 4.5005
R13344 VSS.n206 VSS.n16 4.5005
R13345 VSS.n181 VSS.n16 4.5005
R13346 VSS.n207 VSS.n16 4.5005
R13347 VSS.n180 VSS.n16 4.5005
R13348 VSS.n208 VSS.n16 4.5005
R13349 VSS.n179 VSS.n16 4.5005
R13350 VSS.n209 VSS.n16 4.5005
R13351 VSS.n178 VSS.n16 4.5005
R13352 VSS.n210 VSS.n16 4.5005
R13353 VSS.n177 VSS.n16 4.5005
R13354 VSS.n211 VSS.n16 4.5005
R13355 VSS.n176 VSS.n16 4.5005
R13356 VSS.n212 VSS.n16 4.5005
R13357 VSS.n175 VSS.n16 4.5005
R13358 VSS.n213 VSS.n16 4.5005
R13359 VSS.n174 VSS.n16 4.5005
R13360 VSS.n214 VSS.n16 4.5005
R13361 VSS.n173 VSS.n16 4.5005
R13362 VSS.n215 VSS.n16 4.5005
R13363 VSS.n172 VSS.n16 4.5005
R13364 VSS.n216 VSS.n16 4.5005
R13365 VSS.n171 VSS.n16 4.5005
R13366 VSS.n217 VSS.n16 4.5005
R13367 VSS.n170 VSS.n16 4.5005
R13368 VSS.n218 VSS.n16 4.5005
R13369 VSS.n169 VSS.n16 4.5005
R13370 VSS.n219 VSS.n16 4.5005
R13371 VSS.n168 VSS.n16 4.5005
R13372 VSS.n220 VSS.n16 4.5005
R13373 VSS.n167 VSS.n16 4.5005
R13374 VSS.n221 VSS.n16 4.5005
R13375 VSS.n166 VSS.n16 4.5005
R13376 VSS.n222 VSS.n16 4.5005
R13377 VSS.n165 VSS.n16 4.5005
R13378 VSS.n223 VSS.n16 4.5005
R13379 VSS.n164 VSS.n16 4.5005
R13380 VSS.n224 VSS.n16 4.5005
R13381 VSS.n163 VSS.n16 4.5005
R13382 VSS.n225 VSS.n16 4.5005
R13383 VSS.n162 VSS.n16 4.5005
R13384 VSS.n226 VSS.n16 4.5005
R13385 VSS.n161 VSS.n16 4.5005
R13386 VSS.n227 VSS.n16 4.5005
R13387 VSS.n160 VSS.n16 4.5005
R13388 VSS.n228 VSS.n16 4.5005
R13389 VSS.n159 VSS.n16 4.5005
R13390 VSS.n229 VSS.n16 4.5005
R13391 VSS.n158 VSS.n16 4.5005
R13392 VSS.n230 VSS.n16 4.5005
R13393 VSS.n157 VSS.n16 4.5005
R13394 VSS.n231 VSS.n16 4.5005
R13395 VSS.n156 VSS.n16 4.5005
R13396 VSS.n232 VSS.n16 4.5005
R13397 VSS.n155 VSS.n16 4.5005
R13398 VSS.n233 VSS.n16 4.5005
R13399 VSS.n154 VSS.n16 4.5005
R13400 VSS.n234 VSS.n16 4.5005
R13401 VSS.n153 VSS.n16 4.5005
R13402 VSS.n235 VSS.n16 4.5005
R13403 VSS.n4506 VSS.n16 4.5005
R13404 VSS.n236 VSS.n16 4.5005
R13405 VSS.n152 VSS.n16 4.5005
R13406 VSS.n237 VSS.n16 4.5005
R13407 VSS.n151 VSS.n16 4.5005
R13408 VSS.n238 VSS.n16 4.5005
R13409 VSS.n150 VSS.n16 4.5005
R13410 VSS.n239 VSS.n16 4.5005
R13411 VSS.n149 VSS.n16 4.5005
R13412 VSS.n240 VSS.n16 4.5005
R13413 VSS.n148 VSS.n16 4.5005
R13414 VSS.n241 VSS.n16 4.5005
R13415 VSS.n147 VSS.n16 4.5005
R13416 VSS.n242 VSS.n16 4.5005
R13417 VSS.n146 VSS.n16 4.5005
R13418 VSS.n243 VSS.n16 4.5005
R13419 VSS.n145 VSS.n16 4.5005
R13420 VSS.n244 VSS.n16 4.5005
R13421 VSS.n144 VSS.n16 4.5005
R13422 VSS.n245 VSS.n16 4.5005
R13423 VSS.n143 VSS.n16 4.5005
R13424 VSS.n246 VSS.n16 4.5005
R13425 VSS.n142 VSS.n16 4.5005
R13426 VSS.n247 VSS.n16 4.5005
R13427 VSS.n141 VSS.n16 4.5005
R13428 VSS.n248 VSS.n16 4.5005
R13429 VSS.n140 VSS.n16 4.5005
R13430 VSS.n249 VSS.n16 4.5005
R13431 VSS.n139 VSS.n16 4.5005
R13432 VSS.n250 VSS.n16 4.5005
R13433 VSS.n138 VSS.n16 4.5005
R13434 VSS.n251 VSS.n16 4.5005
R13435 VSS.n137 VSS.n16 4.5005
R13436 VSS.n252 VSS.n16 4.5005
R13437 VSS.n136 VSS.n16 4.5005
R13438 VSS.n253 VSS.n16 4.5005
R13439 VSS.n135 VSS.n16 4.5005
R13440 VSS.n254 VSS.n16 4.5005
R13441 VSS.n134 VSS.n16 4.5005
R13442 VSS.n255 VSS.n16 4.5005
R13443 VSS.n133 VSS.n16 4.5005
R13444 VSS.n256 VSS.n16 4.5005
R13445 VSS.n132 VSS.n16 4.5005
R13446 VSS.n4502 VSS.n16 4.5005
R13447 VSS.n4504 VSS.n16 4.5005
R13448 VSS.n193 VSS.n121 4.5005
R13449 VSS.n195 VSS.n121 4.5005
R13450 VSS.n192 VSS.n121 4.5005
R13451 VSS.n196 VSS.n121 4.5005
R13452 VSS.n191 VSS.n121 4.5005
R13453 VSS.n197 VSS.n121 4.5005
R13454 VSS.n190 VSS.n121 4.5005
R13455 VSS.n198 VSS.n121 4.5005
R13456 VSS.n189 VSS.n121 4.5005
R13457 VSS.n199 VSS.n121 4.5005
R13458 VSS.n188 VSS.n121 4.5005
R13459 VSS.n200 VSS.n121 4.5005
R13460 VSS.n187 VSS.n121 4.5005
R13461 VSS.n201 VSS.n121 4.5005
R13462 VSS.n186 VSS.n121 4.5005
R13463 VSS.n202 VSS.n121 4.5005
R13464 VSS.n185 VSS.n121 4.5005
R13465 VSS.n203 VSS.n121 4.5005
R13466 VSS.n184 VSS.n121 4.5005
R13467 VSS.n204 VSS.n121 4.5005
R13468 VSS.n183 VSS.n121 4.5005
R13469 VSS.n205 VSS.n121 4.5005
R13470 VSS.n182 VSS.n121 4.5005
R13471 VSS.n206 VSS.n121 4.5005
R13472 VSS.n181 VSS.n121 4.5005
R13473 VSS.n207 VSS.n121 4.5005
R13474 VSS.n180 VSS.n121 4.5005
R13475 VSS.n208 VSS.n121 4.5005
R13476 VSS.n179 VSS.n121 4.5005
R13477 VSS.n209 VSS.n121 4.5005
R13478 VSS.n178 VSS.n121 4.5005
R13479 VSS.n210 VSS.n121 4.5005
R13480 VSS.n177 VSS.n121 4.5005
R13481 VSS.n211 VSS.n121 4.5005
R13482 VSS.n176 VSS.n121 4.5005
R13483 VSS.n212 VSS.n121 4.5005
R13484 VSS.n175 VSS.n121 4.5005
R13485 VSS.n213 VSS.n121 4.5005
R13486 VSS.n174 VSS.n121 4.5005
R13487 VSS.n214 VSS.n121 4.5005
R13488 VSS.n173 VSS.n121 4.5005
R13489 VSS.n215 VSS.n121 4.5005
R13490 VSS.n172 VSS.n121 4.5005
R13491 VSS.n216 VSS.n121 4.5005
R13492 VSS.n171 VSS.n121 4.5005
R13493 VSS.n217 VSS.n121 4.5005
R13494 VSS.n170 VSS.n121 4.5005
R13495 VSS.n218 VSS.n121 4.5005
R13496 VSS.n169 VSS.n121 4.5005
R13497 VSS.n219 VSS.n121 4.5005
R13498 VSS.n168 VSS.n121 4.5005
R13499 VSS.n220 VSS.n121 4.5005
R13500 VSS.n167 VSS.n121 4.5005
R13501 VSS.n221 VSS.n121 4.5005
R13502 VSS.n166 VSS.n121 4.5005
R13503 VSS.n222 VSS.n121 4.5005
R13504 VSS.n165 VSS.n121 4.5005
R13505 VSS.n223 VSS.n121 4.5005
R13506 VSS.n164 VSS.n121 4.5005
R13507 VSS.n224 VSS.n121 4.5005
R13508 VSS.n163 VSS.n121 4.5005
R13509 VSS.n225 VSS.n121 4.5005
R13510 VSS.n162 VSS.n121 4.5005
R13511 VSS.n226 VSS.n121 4.5005
R13512 VSS.n161 VSS.n121 4.5005
R13513 VSS.n227 VSS.n121 4.5005
R13514 VSS.n160 VSS.n121 4.5005
R13515 VSS.n228 VSS.n121 4.5005
R13516 VSS.n159 VSS.n121 4.5005
R13517 VSS.n229 VSS.n121 4.5005
R13518 VSS.n158 VSS.n121 4.5005
R13519 VSS.n230 VSS.n121 4.5005
R13520 VSS.n157 VSS.n121 4.5005
R13521 VSS.n231 VSS.n121 4.5005
R13522 VSS.n156 VSS.n121 4.5005
R13523 VSS.n232 VSS.n121 4.5005
R13524 VSS.n155 VSS.n121 4.5005
R13525 VSS.n233 VSS.n121 4.5005
R13526 VSS.n154 VSS.n121 4.5005
R13527 VSS.n234 VSS.n121 4.5005
R13528 VSS.n153 VSS.n121 4.5005
R13529 VSS.n235 VSS.n121 4.5005
R13530 VSS.n4506 VSS.n121 4.5005
R13531 VSS.n236 VSS.n121 4.5005
R13532 VSS.n152 VSS.n121 4.5005
R13533 VSS.n237 VSS.n121 4.5005
R13534 VSS.n151 VSS.n121 4.5005
R13535 VSS.n238 VSS.n121 4.5005
R13536 VSS.n150 VSS.n121 4.5005
R13537 VSS.n239 VSS.n121 4.5005
R13538 VSS.n149 VSS.n121 4.5005
R13539 VSS.n240 VSS.n121 4.5005
R13540 VSS.n148 VSS.n121 4.5005
R13541 VSS.n241 VSS.n121 4.5005
R13542 VSS.n147 VSS.n121 4.5005
R13543 VSS.n242 VSS.n121 4.5005
R13544 VSS.n146 VSS.n121 4.5005
R13545 VSS.n243 VSS.n121 4.5005
R13546 VSS.n145 VSS.n121 4.5005
R13547 VSS.n244 VSS.n121 4.5005
R13548 VSS.n144 VSS.n121 4.5005
R13549 VSS.n245 VSS.n121 4.5005
R13550 VSS.n143 VSS.n121 4.5005
R13551 VSS.n246 VSS.n121 4.5005
R13552 VSS.n142 VSS.n121 4.5005
R13553 VSS.n247 VSS.n121 4.5005
R13554 VSS.n141 VSS.n121 4.5005
R13555 VSS.n248 VSS.n121 4.5005
R13556 VSS.n140 VSS.n121 4.5005
R13557 VSS.n249 VSS.n121 4.5005
R13558 VSS.n139 VSS.n121 4.5005
R13559 VSS.n250 VSS.n121 4.5005
R13560 VSS.n138 VSS.n121 4.5005
R13561 VSS.n251 VSS.n121 4.5005
R13562 VSS.n137 VSS.n121 4.5005
R13563 VSS.n252 VSS.n121 4.5005
R13564 VSS.n136 VSS.n121 4.5005
R13565 VSS.n253 VSS.n121 4.5005
R13566 VSS.n135 VSS.n121 4.5005
R13567 VSS.n254 VSS.n121 4.5005
R13568 VSS.n134 VSS.n121 4.5005
R13569 VSS.n255 VSS.n121 4.5005
R13570 VSS.n133 VSS.n121 4.5005
R13571 VSS.n256 VSS.n121 4.5005
R13572 VSS.n132 VSS.n121 4.5005
R13573 VSS.n4502 VSS.n121 4.5005
R13574 VSS.n4504 VSS.n121 4.5005
R13575 VSS.n193 VSS.n15 4.5005
R13576 VSS.n195 VSS.n15 4.5005
R13577 VSS.n192 VSS.n15 4.5005
R13578 VSS.n196 VSS.n15 4.5005
R13579 VSS.n191 VSS.n15 4.5005
R13580 VSS.n197 VSS.n15 4.5005
R13581 VSS.n190 VSS.n15 4.5005
R13582 VSS.n198 VSS.n15 4.5005
R13583 VSS.n189 VSS.n15 4.5005
R13584 VSS.n199 VSS.n15 4.5005
R13585 VSS.n188 VSS.n15 4.5005
R13586 VSS.n200 VSS.n15 4.5005
R13587 VSS.n187 VSS.n15 4.5005
R13588 VSS.n201 VSS.n15 4.5005
R13589 VSS.n186 VSS.n15 4.5005
R13590 VSS.n202 VSS.n15 4.5005
R13591 VSS.n185 VSS.n15 4.5005
R13592 VSS.n203 VSS.n15 4.5005
R13593 VSS.n184 VSS.n15 4.5005
R13594 VSS.n204 VSS.n15 4.5005
R13595 VSS.n183 VSS.n15 4.5005
R13596 VSS.n205 VSS.n15 4.5005
R13597 VSS.n182 VSS.n15 4.5005
R13598 VSS.n206 VSS.n15 4.5005
R13599 VSS.n181 VSS.n15 4.5005
R13600 VSS.n207 VSS.n15 4.5005
R13601 VSS.n180 VSS.n15 4.5005
R13602 VSS.n208 VSS.n15 4.5005
R13603 VSS.n179 VSS.n15 4.5005
R13604 VSS.n209 VSS.n15 4.5005
R13605 VSS.n178 VSS.n15 4.5005
R13606 VSS.n210 VSS.n15 4.5005
R13607 VSS.n177 VSS.n15 4.5005
R13608 VSS.n211 VSS.n15 4.5005
R13609 VSS.n176 VSS.n15 4.5005
R13610 VSS.n212 VSS.n15 4.5005
R13611 VSS.n175 VSS.n15 4.5005
R13612 VSS.n213 VSS.n15 4.5005
R13613 VSS.n174 VSS.n15 4.5005
R13614 VSS.n214 VSS.n15 4.5005
R13615 VSS.n173 VSS.n15 4.5005
R13616 VSS.n215 VSS.n15 4.5005
R13617 VSS.n172 VSS.n15 4.5005
R13618 VSS.n216 VSS.n15 4.5005
R13619 VSS.n171 VSS.n15 4.5005
R13620 VSS.n217 VSS.n15 4.5005
R13621 VSS.n170 VSS.n15 4.5005
R13622 VSS.n218 VSS.n15 4.5005
R13623 VSS.n169 VSS.n15 4.5005
R13624 VSS.n219 VSS.n15 4.5005
R13625 VSS.n168 VSS.n15 4.5005
R13626 VSS.n220 VSS.n15 4.5005
R13627 VSS.n167 VSS.n15 4.5005
R13628 VSS.n221 VSS.n15 4.5005
R13629 VSS.n166 VSS.n15 4.5005
R13630 VSS.n222 VSS.n15 4.5005
R13631 VSS.n165 VSS.n15 4.5005
R13632 VSS.n223 VSS.n15 4.5005
R13633 VSS.n164 VSS.n15 4.5005
R13634 VSS.n224 VSS.n15 4.5005
R13635 VSS.n163 VSS.n15 4.5005
R13636 VSS.n225 VSS.n15 4.5005
R13637 VSS.n162 VSS.n15 4.5005
R13638 VSS.n226 VSS.n15 4.5005
R13639 VSS.n161 VSS.n15 4.5005
R13640 VSS.n227 VSS.n15 4.5005
R13641 VSS.n160 VSS.n15 4.5005
R13642 VSS.n228 VSS.n15 4.5005
R13643 VSS.n159 VSS.n15 4.5005
R13644 VSS.n229 VSS.n15 4.5005
R13645 VSS.n158 VSS.n15 4.5005
R13646 VSS.n230 VSS.n15 4.5005
R13647 VSS.n157 VSS.n15 4.5005
R13648 VSS.n231 VSS.n15 4.5005
R13649 VSS.n156 VSS.n15 4.5005
R13650 VSS.n232 VSS.n15 4.5005
R13651 VSS.n155 VSS.n15 4.5005
R13652 VSS.n233 VSS.n15 4.5005
R13653 VSS.n154 VSS.n15 4.5005
R13654 VSS.n234 VSS.n15 4.5005
R13655 VSS.n153 VSS.n15 4.5005
R13656 VSS.n235 VSS.n15 4.5005
R13657 VSS.n4506 VSS.n15 4.5005
R13658 VSS.n236 VSS.n15 4.5005
R13659 VSS.n152 VSS.n15 4.5005
R13660 VSS.n237 VSS.n15 4.5005
R13661 VSS.n151 VSS.n15 4.5005
R13662 VSS.n238 VSS.n15 4.5005
R13663 VSS.n150 VSS.n15 4.5005
R13664 VSS.n239 VSS.n15 4.5005
R13665 VSS.n149 VSS.n15 4.5005
R13666 VSS.n240 VSS.n15 4.5005
R13667 VSS.n148 VSS.n15 4.5005
R13668 VSS.n241 VSS.n15 4.5005
R13669 VSS.n147 VSS.n15 4.5005
R13670 VSS.n242 VSS.n15 4.5005
R13671 VSS.n146 VSS.n15 4.5005
R13672 VSS.n243 VSS.n15 4.5005
R13673 VSS.n145 VSS.n15 4.5005
R13674 VSS.n244 VSS.n15 4.5005
R13675 VSS.n144 VSS.n15 4.5005
R13676 VSS.n245 VSS.n15 4.5005
R13677 VSS.n143 VSS.n15 4.5005
R13678 VSS.n246 VSS.n15 4.5005
R13679 VSS.n142 VSS.n15 4.5005
R13680 VSS.n247 VSS.n15 4.5005
R13681 VSS.n141 VSS.n15 4.5005
R13682 VSS.n248 VSS.n15 4.5005
R13683 VSS.n140 VSS.n15 4.5005
R13684 VSS.n249 VSS.n15 4.5005
R13685 VSS.n139 VSS.n15 4.5005
R13686 VSS.n250 VSS.n15 4.5005
R13687 VSS.n138 VSS.n15 4.5005
R13688 VSS.n251 VSS.n15 4.5005
R13689 VSS.n137 VSS.n15 4.5005
R13690 VSS.n252 VSS.n15 4.5005
R13691 VSS.n136 VSS.n15 4.5005
R13692 VSS.n253 VSS.n15 4.5005
R13693 VSS.n135 VSS.n15 4.5005
R13694 VSS.n254 VSS.n15 4.5005
R13695 VSS.n134 VSS.n15 4.5005
R13696 VSS.n255 VSS.n15 4.5005
R13697 VSS.n133 VSS.n15 4.5005
R13698 VSS.n256 VSS.n15 4.5005
R13699 VSS.n132 VSS.n15 4.5005
R13700 VSS.n4502 VSS.n15 4.5005
R13701 VSS.n4504 VSS.n15 4.5005
R13702 VSS.n193 VSS.n122 4.5005
R13703 VSS.n195 VSS.n122 4.5005
R13704 VSS.n192 VSS.n122 4.5005
R13705 VSS.n196 VSS.n122 4.5005
R13706 VSS.n191 VSS.n122 4.5005
R13707 VSS.n197 VSS.n122 4.5005
R13708 VSS.n190 VSS.n122 4.5005
R13709 VSS.n198 VSS.n122 4.5005
R13710 VSS.n189 VSS.n122 4.5005
R13711 VSS.n199 VSS.n122 4.5005
R13712 VSS.n188 VSS.n122 4.5005
R13713 VSS.n200 VSS.n122 4.5005
R13714 VSS.n187 VSS.n122 4.5005
R13715 VSS.n201 VSS.n122 4.5005
R13716 VSS.n186 VSS.n122 4.5005
R13717 VSS.n202 VSS.n122 4.5005
R13718 VSS.n185 VSS.n122 4.5005
R13719 VSS.n203 VSS.n122 4.5005
R13720 VSS.n184 VSS.n122 4.5005
R13721 VSS.n204 VSS.n122 4.5005
R13722 VSS.n183 VSS.n122 4.5005
R13723 VSS.n205 VSS.n122 4.5005
R13724 VSS.n182 VSS.n122 4.5005
R13725 VSS.n206 VSS.n122 4.5005
R13726 VSS.n181 VSS.n122 4.5005
R13727 VSS.n207 VSS.n122 4.5005
R13728 VSS.n180 VSS.n122 4.5005
R13729 VSS.n208 VSS.n122 4.5005
R13730 VSS.n179 VSS.n122 4.5005
R13731 VSS.n209 VSS.n122 4.5005
R13732 VSS.n178 VSS.n122 4.5005
R13733 VSS.n210 VSS.n122 4.5005
R13734 VSS.n177 VSS.n122 4.5005
R13735 VSS.n211 VSS.n122 4.5005
R13736 VSS.n176 VSS.n122 4.5005
R13737 VSS.n212 VSS.n122 4.5005
R13738 VSS.n175 VSS.n122 4.5005
R13739 VSS.n213 VSS.n122 4.5005
R13740 VSS.n174 VSS.n122 4.5005
R13741 VSS.n214 VSS.n122 4.5005
R13742 VSS.n173 VSS.n122 4.5005
R13743 VSS.n215 VSS.n122 4.5005
R13744 VSS.n172 VSS.n122 4.5005
R13745 VSS.n216 VSS.n122 4.5005
R13746 VSS.n171 VSS.n122 4.5005
R13747 VSS.n217 VSS.n122 4.5005
R13748 VSS.n170 VSS.n122 4.5005
R13749 VSS.n218 VSS.n122 4.5005
R13750 VSS.n169 VSS.n122 4.5005
R13751 VSS.n219 VSS.n122 4.5005
R13752 VSS.n168 VSS.n122 4.5005
R13753 VSS.n220 VSS.n122 4.5005
R13754 VSS.n167 VSS.n122 4.5005
R13755 VSS.n221 VSS.n122 4.5005
R13756 VSS.n166 VSS.n122 4.5005
R13757 VSS.n222 VSS.n122 4.5005
R13758 VSS.n165 VSS.n122 4.5005
R13759 VSS.n223 VSS.n122 4.5005
R13760 VSS.n164 VSS.n122 4.5005
R13761 VSS.n224 VSS.n122 4.5005
R13762 VSS.n163 VSS.n122 4.5005
R13763 VSS.n225 VSS.n122 4.5005
R13764 VSS.n162 VSS.n122 4.5005
R13765 VSS.n226 VSS.n122 4.5005
R13766 VSS.n161 VSS.n122 4.5005
R13767 VSS.n227 VSS.n122 4.5005
R13768 VSS.n160 VSS.n122 4.5005
R13769 VSS.n228 VSS.n122 4.5005
R13770 VSS.n159 VSS.n122 4.5005
R13771 VSS.n229 VSS.n122 4.5005
R13772 VSS.n158 VSS.n122 4.5005
R13773 VSS.n230 VSS.n122 4.5005
R13774 VSS.n157 VSS.n122 4.5005
R13775 VSS.n231 VSS.n122 4.5005
R13776 VSS.n156 VSS.n122 4.5005
R13777 VSS.n232 VSS.n122 4.5005
R13778 VSS.n155 VSS.n122 4.5005
R13779 VSS.n233 VSS.n122 4.5005
R13780 VSS.n154 VSS.n122 4.5005
R13781 VSS.n234 VSS.n122 4.5005
R13782 VSS.n153 VSS.n122 4.5005
R13783 VSS.n235 VSS.n122 4.5005
R13784 VSS.n4506 VSS.n122 4.5005
R13785 VSS.n236 VSS.n122 4.5005
R13786 VSS.n152 VSS.n122 4.5005
R13787 VSS.n237 VSS.n122 4.5005
R13788 VSS.n151 VSS.n122 4.5005
R13789 VSS.n238 VSS.n122 4.5005
R13790 VSS.n150 VSS.n122 4.5005
R13791 VSS.n239 VSS.n122 4.5005
R13792 VSS.n149 VSS.n122 4.5005
R13793 VSS.n240 VSS.n122 4.5005
R13794 VSS.n148 VSS.n122 4.5005
R13795 VSS.n241 VSS.n122 4.5005
R13796 VSS.n147 VSS.n122 4.5005
R13797 VSS.n242 VSS.n122 4.5005
R13798 VSS.n146 VSS.n122 4.5005
R13799 VSS.n243 VSS.n122 4.5005
R13800 VSS.n145 VSS.n122 4.5005
R13801 VSS.n244 VSS.n122 4.5005
R13802 VSS.n144 VSS.n122 4.5005
R13803 VSS.n245 VSS.n122 4.5005
R13804 VSS.n143 VSS.n122 4.5005
R13805 VSS.n246 VSS.n122 4.5005
R13806 VSS.n142 VSS.n122 4.5005
R13807 VSS.n247 VSS.n122 4.5005
R13808 VSS.n141 VSS.n122 4.5005
R13809 VSS.n248 VSS.n122 4.5005
R13810 VSS.n140 VSS.n122 4.5005
R13811 VSS.n249 VSS.n122 4.5005
R13812 VSS.n139 VSS.n122 4.5005
R13813 VSS.n250 VSS.n122 4.5005
R13814 VSS.n138 VSS.n122 4.5005
R13815 VSS.n251 VSS.n122 4.5005
R13816 VSS.n137 VSS.n122 4.5005
R13817 VSS.n252 VSS.n122 4.5005
R13818 VSS.n136 VSS.n122 4.5005
R13819 VSS.n253 VSS.n122 4.5005
R13820 VSS.n135 VSS.n122 4.5005
R13821 VSS.n254 VSS.n122 4.5005
R13822 VSS.n134 VSS.n122 4.5005
R13823 VSS.n255 VSS.n122 4.5005
R13824 VSS.n133 VSS.n122 4.5005
R13825 VSS.n256 VSS.n122 4.5005
R13826 VSS.n132 VSS.n122 4.5005
R13827 VSS.n4502 VSS.n122 4.5005
R13828 VSS.n4504 VSS.n122 4.5005
R13829 VSS.n193 VSS.n14 4.5005
R13830 VSS.n195 VSS.n14 4.5005
R13831 VSS.n192 VSS.n14 4.5005
R13832 VSS.n196 VSS.n14 4.5005
R13833 VSS.n191 VSS.n14 4.5005
R13834 VSS.n197 VSS.n14 4.5005
R13835 VSS.n190 VSS.n14 4.5005
R13836 VSS.n198 VSS.n14 4.5005
R13837 VSS.n189 VSS.n14 4.5005
R13838 VSS.n199 VSS.n14 4.5005
R13839 VSS.n188 VSS.n14 4.5005
R13840 VSS.n200 VSS.n14 4.5005
R13841 VSS.n187 VSS.n14 4.5005
R13842 VSS.n201 VSS.n14 4.5005
R13843 VSS.n186 VSS.n14 4.5005
R13844 VSS.n202 VSS.n14 4.5005
R13845 VSS.n185 VSS.n14 4.5005
R13846 VSS.n203 VSS.n14 4.5005
R13847 VSS.n184 VSS.n14 4.5005
R13848 VSS.n204 VSS.n14 4.5005
R13849 VSS.n183 VSS.n14 4.5005
R13850 VSS.n205 VSS.n14 4.5005
R13851 VSS.n182 VSS.n14 4.5005
R13852 VSS.n206 VSS.n14 4.5005
R13853 VSS.n181 VSS.n14 4.5005
R13854 VSS.n207 VSS.n14 4.5005
R13855 VSS.n180 VSS.n14 4.5005
R13856 VSS.n208 VSS.n14 4.5005
R13857 VSS.n179 VSS.n14 4.5005
R13858 VSS.n209 VSS.n14 4.5005
R13859 VSS.n178 VSS.n14 4.5005
R13860 VSS.n210 VSS.n14 4.5005
R13861 VSS.n177 VSS.n14 4.5005
R13862 VSS.n211 VSS.n14 4.5005
R13863 VSS.n176 VSS.n14 4.5005
R13864 VSS.n212 VSS.n14 4.5005
R13865 VSS.n175 VSS.n14 4.5005
R13866 VSS.n213 VSS.n14 4.5005
R13867 VSS.n174 VSS.n14 4.5005
R13868 VSS.n214 VSS.n14 4.5005
R13869 VSS.n173 VSS.n14 4.5005
R13870 VSS.n215 VSS.n14 4.5005
R13871 VSS.n172 VSS.n14 4.5005
R13872 VSS.n216 VSS.n14 4.5005
R13873 VSS.n171 VSS.n14 4.5005
R13874 VSS.n217 VSS.n14 4.5005
R13875 VSS.n170 VSS.n14 4.5005
R13876 VSS.n218 VSS.n14 4.5005
R13877 VSS.n169 VSS.n14 4.5005
R13878 VSS.n219 VSS.n14 4.5005
R13879 VSS.n168 VSS.n14 4.5005
R13880 VSS.n220 VSS.n14 4.5005
R13881 VSS.n167 VSS.n14 4.5005
R13882 VSS.n221 VSS.n14 4.5005
R13883 VSS.n166 VSS.n14 4.5005
R13884 VSS.n222 VSS.n14 4.5005
R13885 VSS.n165 VSS.n14 4.5005
R13886 VSS.n223 VSS.n14 4.5005
R13887 VSS.n164 VSS.n14 4.5005
R13888 VSS.n224 VSS.n14 4.5005
R13889 VSS.n163 VSS.n14 4.5005
R13890 VSS.n225 VSS.n14 4.5005
R13891 VSS.n162 VSS.n14 4.5005
R13892 VSS.n226 VSS.n14 4.5005
R13893 VSS.n161 VSS.n14 4.5005
R13894 VSS.n227 VSS.n14 4.5005
R13895 VSS.n160 VSS.n14 4.5005
R13896 VSS.n228 VSS.n14 4.5005
R13897 VSS.n159 VSS.n14 4.5005
R13898 VSS.n229 VSS.n14 4.5005
R13899 VSS.n158 VSS.n14 4.5005
R13900 VSS.n230 VSS.n14 4.5005
R13901 VSS.n157 VSS.n14 4.5005
R13902 VSS.n231 VSS.n14 4.5005
R13903 VSS.n156 VSS.n14 4.5005
R13904 VSS.n232 VSS.n14 4.5005
R13905 VSS.n155 VSS.n14 4.5005
R13906 VSS.n233 VSS.n14 4.5005
R13907 VSS.n154 VSS.n14 4.5005
R13908 VSS.n234 VSS.n14 4.5005
R13909 VSS.n153 VSS.n14 4.5005
R13910 VSS.n235 VSS.n14 4.5005
R13911 VSS.n4506 VSS.n14 4.5005
R13912 VSS.n236 VSS.n14 4.5005
R13913 VSS.n152 VSS.n14 4.5005
R13914 VSS.n237 VSS.n14 4.5005
R13915 VSS.n151 VSS.n14 4.5005
R13916 VSS.n238 VSS.n14 4.5005
R13917 VSS.n150 VSS.n14 4.5005
R13918 VSS.n239 VSS.n14 4.5005
R13919 VSS.n149 VSS.n14 4.5005
R13920 VSS.n240 VSS.n14 4.5005
R13921 VSS.n148 VSS.n14 4.5005
R13922 VSS.n241 VSS.n14 4.5005
R13923 VSS.n147 VSS.n14 4.5005
R13924 VSS.n242 VSS.n14 4.5005
R13925 VSS.n146 VSS.n14 4.5005
R13926 VSS.n243 VSS.n14 4.5005
R13927 VSS.n145 VSS.n14 4.5005
R13928 VSS.n244 VSS.n14 4.5005
R13929 VSS.n144 VSS.n14 4.5005
R13930 VSS.n245 VSS.n14 4.5005
R13931 VSS.n143 VSS.n14 4.5005
R13932 VSS.n246 VSS.n14 4.5005
R13933 VSS.n142 VSS.n14 4.5005
R13934 VSS.n247 VSS.n14 4.5005
R13935 VSS.n141 VSS.n14 4.5005
R13936 VSS.n248 VSS.n14 4.5005
R13937 VSS.n140 VSS.n14 4.5005
R13938 VSS.n249 VSS.n14 4.5005
R13939 VSS.n139 VSS.n14 4.5005
R13940 VSS.n250 VSS.n14 4.5005
R13941 VSS.n138 VSS.n14 4.5005
R13942 VSS.n251 VSS.n14 4.5005
R13943 VSS.n137 VSS.n14 4.5005
R13944 VSS.n252 VSS.n14 4.5005
R13945 VSS.n136 VSS.n14 4.5005
R13946 VSS.n253 VSS.n14 4.5005
R13947 VSS.n135 VSS.n14 4.5005
R13948 VSS.n254 VSS.n14 4.5005
R13949 VSS.n134 VSS.n14 4.5005
R13950 VSS.n255 VSS.n14 4.5005
R13951 VSS.n133 VSS.n14 4.5005
R13952 VSS.n256 VSS.n14 4.5005
R13953 VSS.n132 VSS.n14 4.5005
R13954 VSS.n4502 VSS.n14 4.5005
R13955 VSS.n4504 VSS.n14 4.5005
R13956 VSS.n193 VSS.n123 4.5005
R13957 VSS.n195 VSS.n123 4.5005
R13958 VSS.n192 VSS.n123 4.5005
R13959 VSS.n196 VSS.n123 4.5005
R13960 VSS.n191 VSS.n123 4.5005
R13961 VSS.n197 VSS.n123 4.5005
R13962 VSS.n190 VSS.n123 4.5005
R13963 VSS.n198 VSS.n123 4.5005
R13964 VSS.n189 VSS.n123 4.5005
R13965 VSS.n199 VSS.n123 4.5005
R13966 VSS.n188 VSS.n123 4.5005
R13967 VSS.n200 VSS.n123 4.5005
R13968 VSS.n187 VSS.n123 4.5005
R13969 VSS.n201 VSS.n123 4.5005
R13970 VSS.n186 VSS.n123 4.5005
R13971 VSS.n202 VSS.n123 4.5005
R13972 VSS.n185 VSS.n123 4.5005
R13973 VSS.n203 VSS.n123 4.5005
R13974 VSS.n184 VSS.n123 4.5005
R13975 VSS.n204 VSS.n123 4.5005
R13976 VSS.n183 VSS.n123 4.5005
R13977 VSS.n205 VSS.n123 4.5005
R13978 VSS.n182 VSS.n123 4.5005
R13979 VSS.n206 VSS.n123 4.5005
R13980 VSS.n181 VSS.n123 4.5005
R13981 VSS.n207 VSS.n123 4.5005
R13982 VSS.n180 VSS.n123 4.5005
R13983 VSS.n208 VSS.n123 4.5005
R13984 VSS.n179 VSS.n123 4.5005
R13985 VSS.n209 VSS.n123 4.5005
R13986 VSS.n178 VSS.n123 4.5005
R13987 VSS.n210 VSS.n123 4.5005
R13988 VSS.n177 VSS.n123 4.5005
R13989 VSS.n211 VSS.n123 4.5005
R13990 VSS.n176 VSS.n123 4.5005
R13991 VSS.n212 VSS.n123 4.5005
R13992 VSS.n175 VSS.n123 4.5005
R13993 VSS.n213 VSS.n123 4.5005
R13994 VSS.n174 VSS.n123 4.5005
R13995 VSS.n214 VSS.n123 4.5005
R13996 VSS.n173 VSS.n123 4.5005
R13997 VSS.n215 VSS.n123 4.5005
R13998 VSS.n172 VSS.n123 4.5005
R13999 VSS.n216 VSS.n123 4.5005
R14000 VSS.n171 VSS.n123 4.5005
R14001 VSS.n217 VSS.n123 4.5005
R14002 VSS.n170 VSS.n123 4.5005
R14003 VSS.n218 VSS.n123 4.5005
R14004 VSS.n169 VSS.n123 4.5005
R14005 VSS.n219 VSS.n123 4.5005
R14006 VSS.n168 VSS.n123 4.5005
R14007 VSS.n220 VSS.n123 4.5005
R14008 VSS.n167 VSS.n123 4.5005
R14009 VSS.n221 VSS.n123 4.5005
R14010 VSS.n166 VSS.n123 4.5005
R14011 VSS.n222 VSS.n123 4.5005
R14012 VSS.n165 VSS.n123 4.5005
R14013 VSS.n223 VSS.n123 4.5005
R14014 VSS.n164 VSS.n123 4.5005
R14015 VSS.n224 VSS.n123 4.5005
R14016 VSS.n163 VSS.n123 4.5005
R14017 VSS.n225 VSS.n123 4.5005
R14018 VSS.n162 VSS.n123 4.5005
R14019 VSS.n226 VSS.n123 4.5005
R14020 VSS.n161 VSS.n123 4.5005
R14021 VSS.n227 VSS.n123 4.5005
R14022 VSS.n160 VSS.n123 4.5005
R14023 VSS.n228 VSS.n123 4.5005
R14024 VSS.n159 VSS.n123 4.5005
R14025 VSS.n229 VSS.n123 4.5005
R14026 VSS.n158 VSS.n123 4.5005
R14027 VSS.n230 VSS.n123 4.5005
R14028 VSS.n157 VSS.n123 4.5005
R14029 VSS.n231 VSS.n123 4.5005
R14030 VSS.n156 VSS.n123 4.5005
R14031 VSS.n232 VSS.n123 4.5005
R14032 VSS.n155 VSS.n123 4.5005
R14033 VSS.n233 VSS.n123 4.5005
R14034 VSS.n154 VSS.n123 4.5005
R14035 VSS.n234 VSS.n123 4.5005
R14036 VSS.n153 VSS.n123 4.5005
R14037 VSS.n235 VSS.n123 4.5005
R14038 VSS.n4506 VSS.n123 4.5005
R14039 VSS.n236 VSS.n123 4.5005
R14040 VSS.n152 VSS.n123 4.5005
R14041 VSS.n237 VSS.n123 4.5005
R14042 VSS.n151 VSS.n123 4.5005
R14043 VSS.n238 VSS.n123 4.5005
R14044 VSS.n150 VSS.n123 4.5005
R14045 VSS.n239 VSS.n123 4.5005
R14046 VSS.n149 VSS.n123 4.5005
R14047 VSS.n240 VSS.n123 4.5005
R14048 VSS.n148 VSS.n123 4.5005
R14049 VSS.n241 VSS.n123 4.5005
R14050 VSS.n147 VSS.n123 4.5005
R14051 VSS.n242 VSS.n123 4.5005
R14052 VSS.n146 VSS.n123 4.5005
R14053 VSS.n243 VSS.n123 4.5005
R14054 VSS.n145 VSS.n123 4.5005
R14055 VSS.n244 VSS.n123 4.5005
R14056 VSS.n144 VSS.n123 4.5005
R14057 VSS.n245 VSS.n123 4.5005
R14058 VSS.n143 VSS.n123 4.5005
R14059 VSS.n246 VSS.n123 4.5005
R14060 VSS.n142 VSS.n123 4.5005
R14061 VSS.n247 VSS.n123 4.5005
R14062 VSS.n141 VSS.n123 4.5005
R14063 VSS.n248 VSS.n123 4.5005
R14064 VSS.n140 VSS.n123 4.5005
R14065 VSS.n249 VSS.n123 4.5005
R14066 VSS.n139 VSS.n123 4.5005
R14067 VSS.n250 VSS.n123 4.5005
R14068 VSS.n138 VSS.n123 4.5005
R14069 VSS.n251 VSS.n123 4.5005
R14070 VSS.n137 VSS.n123 4.5005
R14071 VSS.n252 VSS.n123 4.5005
R14072 VSS.n136 VSS.n123 4.5005
R14073 VSS.n253 VSS.n123 4.5005
R14074 VSS.n135 VSS.n123 4.5005
R14075 VSS.n254 VSS.n123 4.5005
R14076 VSS.n134 VSS.n123 4.5005
R14077 VSS.n255 VSS.n123 4.5005
R14078 VSS.n133 VSS.n123 4.5005
R14079 VSS.n256 VSS.n123 4.5005
R14080 VSS.n132 VSS.n123 4.5005
R14081 VSS.n4502 VSS.n123 4.5005
R14082 VSS.n4504 VSS.n123 4.5005
R14083 VSS.n193 VSS.n13 4.5005
R14084 VSS.n195 VSS.n13 4.5005
R14085 VSS.n192 VSS.n13 4.5005
R14086 VSS.n196 VSS.n13 4.5005
R14087 VSS.n191 VSS.n13 4.5005
R14088 VSS.n197 VSS.n13 4.5005
R14089 VSS.n190 VSS.n13 4.5005
R14090 VSS.n198 VSS.n13 4.5005
R14091 VSS.n189 VSS.n13 4.5005
R14092 VSS.n199 VSS.n13 4.5005
R14093 VSS.n188 VSS.n13 4.5005
R14094 VSS.n200 VSS.n13 4.5005
R14095 VSS.n187 VSS.n13 4.5005
R14096 VSS.n201 VSS.n13 4.5005
R14097 VSS.n186 VSS.n13 4.5005
R14098 VSS.n202 VSS.n13 4.5005
R14099 VSS.n185 VSS.n13 4.5005
R14100 VSS.n203 VSS.n13 4.5005
R14101 VSS.n184 VSS.n13 4.5005
R14102 VSS.n204 VSS.n13 4.5005
R14103 VSS.n183 VSS.n13 4.5005
R14104 VSS.n205 VSS.n13 4.5005
R14105 VSS.n182 VSS.n13 4.5005
R14106 VSS.n206 VSS.n13 4.5005
R14107 VSS.n181 VSS.n13 4.5005
R14108 VSS.n207 VSS.n13 4.5005
R14109 VSS.n180 VSS.n13 4.5005
R14110 VSS.n208 VSS.n13 4.5005
R14111 VSS.n179 VSS.n13 4.5005
R14112 VSS.n209 VSS.n13 4.5005
R14113 VSS.n178 VSS.n13 4.5005
R14114 VSS.n210 VSS.n13 4.5005
R14115 VSS.n177 VSS.n13 4.5005
R14116 VSS.n211 VSS.n13 4.5005
R14117 VSS.n176 VSS.n13 4.5005
R14118 VSS.n212 VSS.n13 4.5005
R14119 VSS.n175 VSS.n13 4.5005
R14120 VSS.n213 VSS.n13 4.5005
R14121 VSS.n174 VSS.n13 4.5005
R14122 VSS.n214 VSS.n13 4.5005
R14123 VSS.n173 VSS.n13 4.5005
R14124 VSS.n215 VSS.n13 4.5005
R14125 VSS.n172 VSS.n13 4.5005
R14126 VSS.n216 VSS.n13 4.5005
R14127 VSS.n171 VSS.n13 4.5005
R14128 VSS.n217 VSS.n13 4.5005
R14129 VSS.n170 VSS.n13 4.5005
R14130 VSS.n218 VSS.n13 4.5005
R14131 VSS.n169 VSS.n13 4.5005
R14132 VSS.n219 VSS.n13 4.5005
R14133 VSS.n168 VSS.n13 4.5005
R14134 VSS.n220 VSS.n13 4.5005
R14135 VSS.n167 VSS.n13 4.5005
R14136 VSS.n221 VSS.n13 4.5005
R14137 VSS.n166 VSS.n13 4.5005
R14138 VSS.n222 VSS.n13 4.5005
R14139 VSS.n165 VSS.n13 4.5005
R14140 VSS.n223 VSS.n13 4.5005
R14141 VSS.n164 VSS.n13 4.5005
R14142 VSS.n224 VSS.n13 4.5005
R14143 VSS.n163 VSS.n13 4.5005
R14144 VSS.n225 VSS.n13 4.5005
R14145 VSS.n162 VSS.n13 4.5005
R14146 VSS.n226 VSS.n13 4.5005
R14147 VSS.n161 VSS.n13 4.5005
R14148 VSS.n227 VSS.n13 4.5005
R14149 VSS.n160 VSS.n13 4.5005
R14150 VSS.n228 VSS.n13 4.5005
R14151 VSS.n159 VSS.n13 4.5005
R14152 VSS.n229 VSS.n13 4.5005
R14153 VSS.n158 VSS.n13 4.5005
R14154 VSS.n230 VSS.n13 4.5005
R14155 VSS.n157 VSS.n13 4.5005
R14156 VSS.n231 VSS.n13 4.5005
R14157 VSS.n156 VSS.n13 4.5005
R14158 VSS.n232 VSS.n13 4.5005
R14159 VSS.n155 VSS.n13 4.5005
R14160 VSS.n233 VSS.n13 4.5005
R14161 VSS.n154 VSS.n13 4.5005
R14162 VSS.n234 VSS.n13 4.5005
R14163 VSS.n153 VSS.n13 4.5005
R14164 VSS.n235 VSS.n13 4.5005
R14165 VSS.n4506 VSS.n13 4.5005
R14166 VSS.n236 VSS.n13 4.5005
R14167 VSS.n152 VSS.n13 4.5005
R14168 VSS.n237 VSS.n13 4.5005
R14169 VSS.n151 VSS.n13 4.5005
R14170 VSS.n238 VSS.n13 4.5005
R14171 VSS.n150 VSS.n13 4.5005
R14172 VSS.n239 VSS.n13 4.5005
R14173 VSS.n149 VSS.n13 4.5005
R14174 VSS.n240 VSS.n13 4.5005
R14175 VSS.n148 VSS.n13 4.5005
R14176 VSS.n241 VSS.n13 4.5005
R14177 VSS.n147 VSS.n13 4.5005
R14178 VSS.n242 VSS.n13 4.5005
R14179 VSS.n146 VSS.n13 4.5005
R14180 VSS.n243 VSS.n13 4.5005
R14181 VSS.n145 VSS.n13 4.5005
R14182 VSS.n244 VSS.n13 4.5005
R14183 VSS.n144 VSS.n13 4.5005
R14184 VSS.n245 VSS.n13 4.5005
R14185 VSS.n143 VSS.n13 4.5005
R14186 VSS.n246 VSS.n13 4.5005
R14187 VSS.n142 VSS.n13 4.5005
R14188 VSS.n247 VSS.n13 4.5005
R14189 VSS.n141 VSS.n13 4.5005
R14190 VSS.n248 VSS.n13 4.5005
R14191 VSS.n140 VSS.n13 4.5005
R14192 VSS.n249 VSS.n13 4.5005
R14193 VSS.n139 VSS.n13 4.5005
R14194 VSS.n250 VSS.n13 4.5005
R14195 VSS.n138 VSS.n13 4.5005
R14196 VSS.n251 VSS.n13 4.5005
R14197 VSS.n137 VSS.n13 4.5005
R14198 VSS.n252 VSS.n13 4.5005
R14199 VSS.n136 VSS.n13 4.5005
R14200 VSS.n253 VSS.n13 4.5005
R14201 VSS.n135 VSS.n13 4.5005
R14202 VSS.n254 VSS.n13 4.5005
R14203 VSS.n134 VSS.n13 4.5005
R14204 VSS.n255 VSS.n13 4.5005
R14205 VSS.n133 VSS.n13 4.5005
R14206 VSS.n256 VSS.n13 4.5005
R14207 VSS.n132 VSS.n13 4.5005
R14208 VSS.n4502 VSS.n13 4.5005
R14209 VSS.n4504 VSS.n13 4.5005
R14210 VSS.n193 VSS.n124 4.5005
R14211 VSS.n195 VSS.n124 4.5005
R14212 VSS.n192 VSS.n124 4.5005
R14213 VSS.n196 VSS.n124 4.5005
R14214 VSS.n191 VSS.n124 4.5005
R14215 VSS.n197 VSS.n124 4.5005
R14216 VSS.n190 VSS.n124 4.5005
R14217 VSS.n198 VSS.n124 4.5005
R14218 VSS.n189 VSS.n124 4.5005
R14219 VSS.n199 VSS.n124 4.5005
R14220 VSS.n188 VSS.n124 4.5005
R14221 VSS.n200 VSS.n124 4.5005
R14222 VSS.n187 VSS.n124 4.5005
R14223 VSS.n201 VSS.n124 4.5005
R14224 VSS.n186 VSS.n124 4.5005
R14225 VSS.n202 VSS.n124 4.5005
R14226 VSS.n185 VSS.n124 4.5005
R14227 VSS.n203 VSS.n124 4.5005
R14228 VSS.n184 VSS.n124 4.5005
R14229 VSS.n204 VSS.n124 4.5005
R14230 VSS.n183 VSS.n124 4.5005
R14231 VSS.n205 VSS.n124 4.5005
R14232 VSS.n182 VSS.n124 4.5005
R14233 VSS.n206 VSS.n124 4.5005
R14234 VSS.n181 VSS.n124 4.5005
R14235 VSS.n207 VSS.n124 4.5005
R14236 VSS.n180 VSS.n124 4.5005
R14237 VSS.n208 VSS.n124 4.5005
R14238 VSS.n179 VSS.n124 4.5005
R14239 VSS.n209 VSS.n124 4.5005
R14240 VSS.n178 VSS.n124 4.5005
R14241 VSS.n210 VSS.n124 4.5005
R14242 VSS.n177 VSS.n124 4.5005
R14243 VSS.n211 VSS.n124 4.5005
R14244 VSS.n176 VSS.n124 4.5005
R14245 VSS.n212 VSS.n124 4.5005
R14246 VSS.n175 VSS.n124 4.5005
R14247 VSS.n213 VSS.n124 4.5005
R14248 VSS.n174 VSS.n124 4.5005
R14249 VSS.n214 VSS.n124 4.5005
R14250 VSS.n173 VSS.n124 4.5005
R14251 VSS.n215 VSS.n124 4.5005
R14252 VSS.n172 VSS.n124 4.5005
R14253 VSS.n216 VSS.n124 4.5005
R14254 VSS.n171 VSS.n124 4.5005
R14255 VSS.n217 VSS.n124 4.5005
R14256 VSS.n170 VSS.n124 4.5005
R14257 VSS.n218 VSS.n124 4.5005
R14258 VSS.n169 VSS.n124 4.5005
R14259 VSS.n219 VSS.n124 4.5005
R14260 VSS.n168 VSS.n124 4.5005
R14261 VSS.n220 VSS.n124 4.5005
R14262 VSS.n167 VSS.n124 4.5005
R14263 VSS.n221 VSS.n124 4.5005
R14264 VSS.n166 VSS.n124 4.5005
R14265 VSS.n222 VSS.n124 4.5005
R14266 VSS.n165 VSS.n124 4.5005
R14267 VSS.n223 VSS.n124 4.5005
R14268 VSS.n164 VSS.n124 4.5005
R14269 VSS.n224 VSS.n124 4.5005
R14270 VSS.n163 VSS.n124 4.5005
R14271 VSS.n225 VSS.n124 4.5005
R14272 VSS.n162 VSS.n124 4.5005
R14273 VSS.n226 VSS.n124 4.5005
R14274 VSS.n161 VSS.n124 4.5005
R14275 VSS.n227 VSS.n124 4.5005
R14276 VSS.n160 VSS.n124 4.5005
R14277 VSS.n228 VSS.n124 4.5005
R14278 VSS.n159 VSS.n124 4.5005
R14279 VSS.n229 VSS.n124 4.5005
R14280 VSS.n158 VSS.n124 4.5005
R14281 VSS.n230 VSS.n124 4.5005
R14282 VSS.n157 VSS.n124 4.5005
R14283 VSS.n231 VSS.n124 4.5005
R14284 VSS.n156 VSS.n124 4.5005
R14285 VSS.n232 VSS.n124 4.5005
R14286 VSS.n155 VSS.n124 4.5005
R14287 VSS.n233 VSS.n124 4.5005
R14288 VSS.n154 VSS.n124 4.5005
R14289 VSS.n234 VSS.n124 4.5005
R14290 VSS.n153 VSS.n124 4.5005
R14291 VSS.n235 VSS.n124 4.5005
R14292 VSS.n4506 VSS.n124 4.5005
R14293 VSS.n236 VSS.n124 4.5005
R14294 VSS.n152 VSS.n124 4.5005
R14295 VSS.n237 VSS.n124 4.5005
R14296 VSS.n151 VSS.n124 4.5005
R14297 VSS.n238 VSS.n124 4.5005
R14298 VSS.n150 VSS.n124 4.5005
R14299 VSS.n239 VSS.n124 4.5005
R14300 VSS.n149 VSS.n124 4.5005
R14301 VSS.n240 VSS.n124 4.5005
R14302 VSS.n148 VSS.n124 4.5005
R14303 VSS.n241 VSS.n124 4.5005
R14304 VSS.n147 VSS.n124 4.5005
R14305 VSS.n242 VSS.n124 4.5005
R14306 VSS.n146 VSS.n124 4.5005
R14307 VSS.n243 VSS.n124 4.5005
R14308 VSS.n145 VSS.n124 4.5005
R14309 VSS.n244 VSS.n124 4.5005
R14310 VSS.n144 VSS.n124 4.5005
R14311 VSS.n245 VSS.n124 4.5005
R14312 VSS.n143 VSS.n124 4.5005
R14313 VSS.n246 VSS.n124 4.5005
R14314 VSS.n142 VSS.n124 4.5005
R14315 VSS.n247 VSS.n124 4.5005
R14316 VSS.n141 VSS.n124 4.5005
R14317 VSS.n248 VSS.n124 4.5005
R14318 VSS.n140 VSS.n124 4.5005
R14319 VSS.n249 VSS.n124 4.5005
R14320 VSS.n139 VSS.n124 4.5005
R14321 VSS.n250 VSS.n124 4.5005
R14322 VSS.n138 VSS.n124 4.5005
R14323 VSS.n251 VSS.n124 4.5005
R14324 VSS.n137 VSS.n124 4.5005
R14325 VSS.n252 VSS.n124 4.5005
R14326 VSS.n136 VSS.n124 4.5005
R14327 VSS.n253 VSS.n124 4.5005
R14328 VSS.n135 VSS.n124 4.5005
R14329 VSS.n254 VSS.n124 4.5005
R14330 VSS.n134 VSS.n124 4.5005
R14331 VSS.n255 VSS.n124 4.5005
R14332 VSS.n133 VSS.n124 4.5005
R14333 VSS.n256 VSS.n124 4.5005
R14334 VSS.n132 VSS.n124 4.5005
R14335 VSS.n4502 VSS.n124 4.5005
R14336 VSS.n4504 VSS.n124 4.5005
R14337 VSS.n193 VSS.n12 4.5005
R14338 VSS.n195 VSS.n12 4.5005
R14339 VSS.n192 VSS.n12 4.5005
R14340 VSS.n196 VSS.n12 4.5005
R14341 VSS.n191 VSS.n12 4.5005
R14342 VSS.n197 VSS.n12 4.5005
R14343 VSS.n190 VSS.n12 4.5005
R14344 VSS.n198 VSS.n12 4.5005
R14345 VSS.n189 VSS.n12 4.5005
R14346 VSS.n199 VSS.n12 4.5005
R14347 VSS.n188 VSS.n12 4.5005
R14348 VSS.n200 VSS.n12 4.5005
R14349 VSS.n187 VSS.n12 4.5005
R14350 VSS.n201 VSS.n12 4.5005
R14351 VSS.n186 VSS.n12 4.5005
R14352 VSS.n202 VSS.n12 4.5005
R14353 VSS.n185 VSS.n12 4.5005
R14354 VSS.n203 VSS.n12 4.5005
R14355 VSS.n184 VSS.n12 4.5005
R14356 VSS.n204 VSS.n12 4.5005
R14357 VSS.n183 VSS.n12 4.5005
R14358 VSS.n205 VSS.n12 4.5005
R14359 VSS.n182 VSS.n12 4.5005
R14360 VSS.n206 VSS.n12 4.5005
R14361 VSS.n181 VSS.n12 4.5005
R14362 VSS.n207 VSS.n12 4.5005
R14363 VSS.n180 VSS.n12 4.5005
R14364 VSS.n208 VSS.n12 4.5005
R14365 VSS.n179 VSS.n12 4.5005
R14366 VSS.n209 VSS.n12 4.5005
R14367 VSS.n178 VSS.n12 4.5005
R14368 VSS.n210 VSS.n12 4.5005
R14369 VSS.n177 VSS.n12 4.5005
R14370 VSS.n211 VSS.n12 4.5005
R14371 VSS.n176 VSS.n12 4.5005
R14372 VSS.n212 VSS.n12 4.5005
R14373 VSS.n175 VSS.n12 4.5005
R14374 VSS.n213 VSS.n12 4.5005
R14375 VSS.n174 VSS.n12 4.5005
R14376 VSS.n214 VSS.n12 4.5005
R14377 VSS.n173 VSS.n12 4.5005
R14378 VSS.n215 VSS.n12 4.5005
R14379 VSS.n172 VSS.n12 4.5005
R14380 VSS.n216 VSS.n12 4.5005
R14381 VSS.n171 VSS.n12 4.5005
R14382 VSS.n217 VSS.n12 4.5005
R14383 VSS.n170 VSS.n12 4.5005
R14384 VSS.n218 VSS.n12 4.5005
R14385 VSS.n169 VSS.n12 4.5005
R14386 VSS.n219 VSS.n12 4.5005
R14387 VSS.n168 VSS.n12 4.5005
R14388 VSS.n220 VSS.n12 4.5005
R14389 VSS.n167 VSS.n12 4.5005
R14390 VSS.n221 VSS.n12 4.5005
R14391 VSS.n166 VSS.n12 4.5005
R14392 VSS.n222 VSS.n12 4.5005
R14393 VSS.n165 VSS.n12 4.5005
R14394 VSS.n223 VSS.n12 4.5005
R14395 VSS.n164 VSS.n12 4.5005
R14396 VSS.n224 VSS.n12 4.5005
R14397 VSS.n163 VSS.n12 4.5005
R14398 VSS.n225 VSS.n12 4.5005
R14399 VSS.n162 VSS.n12 4.5005
R14400 VSS.n226 VSS.n12 4.5005
R14401 VSS.n161 VSS.n12 4.5005
R14402 VSS.n227 VSS.n12 4.5005
R14403 VSS.n160 VSS.n12 4.5005
R14404 VSS.n228 VSS.n12 4.5005
R14405 VSS.n159 VSS.n12 4.5005
R14406 VSS.n229 VSS.n12 4.5005
R14407 VSS.n158 VSS.n12 4.5005
R14408 VSS.n230 VSS.n12 4.5005
R14409 VSS.n157 VSS.n12 4.5005
R14410 VSS.n231 VSS.n12 4.5005
R14411 VSS.n156 VSS.n12 4.5005
R14412 VSS.n232 VSS.n12 4.5005
R14413 VSS.n155 VSS.n12 4.5005
R14414 VSS.n233 VSS.n12 4.5005
R14415 VSS.n154 VSS.n12 4.5005
R14416 VSS.n234 VSS.n12 4.5005
R14417 VSS.n153 VSS.n12 4.5005
R14418 VSS.n235 VSS.n12 4.5005
R14419 VSS.n4506 VSS.n12 4.5005
R14420 VSS.n236 VSS.n12 4.5005
R14421 VSS.n152 VSS.n12 4.5005
R14422 VSS.n237 VSS.n12 4.5005
R14423 VSS.n151 VSS.n12 4.5005
R14424 VSS.n238 VSS.n12 4.5005
R14425 VSS.n150 VSS.n12 4.5005
R14426 VSS.n239 VSS.n12 4.5005
R14427 VSS.n149 VSS.n12 4.5005
R14428 VSS.n240 VSS.n12 4.5005
R14429 VSS.n148 VSS.n12 4.5005
R14430 VSS.n241 VSS.n12 4.5005
R14431 VSS.n147 VSS.n12 4.5005
R14432 VSS.n242 VSS.n12 4.5005
R14433 VSS.n146 VSS.n12 4.5005
R14434 VSS.n243 VSS.n12 4.5005
R14435 VSS.n145 VSS.n12 4.5005
R14436 VSS.n244 VSS.n12 4.5005
R14437 VSS.n144 VSS.n12 4.5005
R14438 VSS.n245 VSS.n12 4.5005
R14439 VSS.n143 VSS.n12 4.5005
R14440 VSS.n246 VSS.n12 4.5005
R14441 VSS.n142 VSS.n12 4.5005
R14442 VSS.n247 VSS.n12 4.5005
R14443 VSS.n141 VSS.n12 4.5005
R14444 VSS.n248 VSS.n12 4.5005
R14445 VSS.n140 VSS.n12 4.5005
R14446 VSS.n249 VSS.n12 4.5005
R14447 VSS.n139 VSS.n12 4.5005
R14448 VSS.n250 VSS.n12 4.5005
R14449 VSS.n138 VSS.n12 4.5005
R14450 VSS.n251 VSS.n12 4.5005
R14451 VSS.n137 VSS.n12 4.5005
R14452 VSS.n252 VSS.n12 4.5005
R14453 VSS.n136 VSS.n12 4.5005
R14454 VSS.n253 VSS.n12 4.5005
R14455 VSS.n135 VSS.n12 4.5005
R14456 VSS.n254 VSS.n12 4.5005
R14457 VSS.n134 VSS.n12 4.5005
R14458 VSS.n255 VSS.n12 4.5005
R14459 VSS.n133 VSS.n12 4.5005
R14460 VSS.n256 VSS.n12 4.5005
R14461 VSS.n132 VSS.n12 4.5005
R14462 VSS.n4502 VSS.n12 4.5005
R14463 VSS.n4504 VSS.n12 4.5005
R14464 VSS.n193 VSS.n125 4.5005
R14465 VSS.n195 VSS.n125 4.5005
R14466 VSS.n192 VSS.n125 4.5005
R14467 VSS.n196 VSS.n125 4.5005
R14468 VSS.n191 VSS.n125 4.5005
R14469 VSS.n197 VSS.n125 4.5005
R14470 VSS.n190 VSS.n125 4.5005
R14471 VSS.n198 VSS.n125 4.5005
R14472 VSS.n189 VSS.n125 4.5005
R14473 VSS.n199 VSS.n125 4.5005
R14474 VSS.n188 VSS.n125 4.5005
R14475 VSS.n200 VSS.n125 4.5005
R14476 VSS.n187 VSS.n125 4.5005
R14477 VSS.n201 VSS.n125 4.5005
R14478 VSS.n186 VSS.n125 4.5005
R14479 VSS.n202 VSS.n125 4.5005
R14480 VSS.n185 VSS.n125 4.5005
R14481 VSS.n203 VSS.n125 4.5005
R14482 VSS.n184 VSS.n125 4.5005
R14483 VSS.n204 VSS.n125 4.5005
R14484 VSS.n183 VSS.n125 4.5005
R14485 VSS.n205 VSS.n125 4.5005
R14486 VSS.n182 VSS.n125 4.5005
R14487 VSS.n206 VSS.n125 4.5005
R14488 VSS.n181 VSS.n125 4.5005
R14489 VSS.n207 VSS.n125 4.5005
R14490 VSS.n180 VSS.n125 4.5005
R14491 VSS.n208 VSS.n125 4.5005
R14492 VSS.n179 VSS.n125 4.5005
R14493 VSS.n209 VSS.n125 4.5005
R14494 VSS.n178 VSS.n125 4.5005
R14495 VSS.n210 VSS.n125 4.5005
R14496 VSS.n177 VSS.n125 4.5005
R14497 VSS.n211 VSS.n125 4.5005
R14498 VSS.n176 VSS.n125 4.5005
R14499 VSS.n212 VSS.n125 4.5005
R14500 VSS.n175 VSS.n125 4.5005
R14501 VSS.n213 VSS.n125 4.5005
R14502 VSS.n174 VSS.n125 4.5005
R14503 VSS.n214 VSS.n125 4.5005
R14504 VSS.n173 VSS.n125 4.5005
R14505 VSS.n215 VSS.n125 4.5005
R14506 VSS.n172 VSS.n125 4.5005
R14507 VSS.n216 VSS.n125 4.5005
R14508 VSS.n171 VSS.n125 4.5005
R14509 VSS.n217 VSS.n125 4.5005
R14510 VSS.n170 VSS.n125 4.5005
R14511 VSS.n218 VSS.n125 4.5005
R14512 VSS.n169 VSS.n125 4.5005
R14513 VSS.n219 VSS.n125 4.5005
R14514 VSS.n168 VSS.n125 4.5005
R14515 VSS.n220 VSS.n125 4.5005
R14516 VSS.n167 VSS.n125 4.5005
R14517 VSS.n221 VSS.n125 4.5005
R14518 VSS.n166 VSS.n125 4.5005
R14519 VSS.n222 VSS.n125 4.5005
R14520 VSS.n165 VSS.n125 4.5005
R14521 VSS.n223 VSS.n125 4.5005
R14522 VSS.n164 VSS.n125 4.5005
R14523 VSS.n224 VSS.n125 4.5005
R14524 VSS.n163 VSS.n125 4.5005
R14525 VSS.n225 VSS.n125 4.5005
R14526 VSS.n162 VSS.n125 4.5005
R14527 VSS.n226 VSS.n125 4.5005
R14528 VSS.n161 VSS.n125 4.5005
R14529 VSS.n227 VSS.n125 4.5005
R14530 VSS.n160 VSS.n125 4.5005
R14531 VSS.n228 VSS.n125 4.5005
R14532 VSS.n159 VSS.n125 4.5005
R14533 VSS.n229 VSS.n125 4.5005
R14534 VSS.n158 VSS.n125 4.5005
R14535 VSS.n230 VSS.n125 4.5005
R14536 VSS.n157 VSS.n125 4.5005
R14537 VSS.n231 VSS.n125 4.5005
R14538 VSS.n156 VSS.n125 4.5005
R14539 VSS.n232 VSS.n125 4.5005
R14540 VSS.n155 VSS.n125 4.5005
R14541 VSS.n233 VSS.n125 4.5005
R14542 VSS.n154 VSS.n125 4.5005
R14543 VSS.n234 VSS.n125 4.5005
R14544 VSS.n153 VSS.n125 4.5005
R14545 VSS.n235 VSS.n125 4.5005
R14546 VSS.n4506 VSS.n125 4.5005
R14547 VSS.n236 VSS.n125 4.5005
R14548 VSS.n152 VSS.n125 4.5005
R14549 VSS.n237 VSS.n125 4.5005
R14550 VSS.n151 VSS.n125 4.5005
R14551 VSS.n238 VSS.n125 4.5005
R14552 VSS.n150 VSS.n125 4.5005
R14553 VSS.n239 VSS.n125 4.5005
R14554 VSS.n149 VSS.n125 4.5005
R14555 VSS.n240 VSS.n125 4.5005
R14556 VSS.n148 VSS.n125 4.5005
R14557 VSS.n241 VSS.n125 4.5005
R14558 VSS.n147 VSS.n125 4.5005
R14559 VSS.n242 VSS.n125 4.5005
R14560 VSS.n146 VSS.n125 4.5005
R14561 VSS.n243 VSS.n125 4.5005
R14562 VSS.n145 VSS.n125 4.5005
R14563 VSS.n244 VSS.n125 4.5005
R14564 VSS.n144 VSS.n125 4.5005
R14565 VSS.n245 VSS.n125 4.5005
R14566 VSS.n143 VSS.n125 4.5005
R14567 VSS.n246 VSS.n125 4.5005
R14568 VSS.n142 VSS.n125 4.5005
R14569 VSS.n247 VSS.n125 4.5005
R14570 VSS.n141 VSS.n125 4.5005
R14571 VSS.n248 VSS.n125 4.5005
R14572 VSS.n140 VSS.n125 4.5005
R14573 VSS.n249 VSS.n125 4.5005
R14574 VSS.n139 VSS.n125 4.5005
R14575 VSS.n250 VSS.n125 4.5005
R14576 VSS.n138 VSS.n125 4.5005
R14577 VSS.n251 VSS.n125 4.5005
R14578 VSS.n137 VSS.n125 4.5005
R14579 VSS.n252 VSS.n125 4.5005
R14580 VSS.n136 VSS.n125 4.5005
R14581 VSS.n253 VSS.n125 4.5005
R14582 VSS.n135 VSS.n125 4.5005
R14583 VSS.n254 VSS.n125 4.5005
R14584 VSS.n134 VSS.n125 4.5005
R14585 VSS.n255 VSS.n125 4.5005
R14586 VSS.n133 VSS.n125 4.5005
R14587 VSS.n256 VSS.n125 4.5005
R14588 VSS.n132 VSS.n125 4.5005
R14589 VSS.n4502 VSS.n125 4.5005
R14590 VSS.n4504 VSS.n125 4.5005
R14591 VSS.n193 VSS.n11 4.5005
R14592 VSS.n195 VSS.n11 4.5005
R14593 VSS.n192 VSS.n11 4.5005
R14594 VSS.n196 VSS.n11 4.5005
R14595 VSS.n191 VSS.n11 4.5005
R14596 VSS.n197 VSS.n11 4.5005
R14597 VSS.n190 VSS.n11 4.5005
R14598 VSS.n198 VSS.n11 4.5005
R14599 VSS.n189 VSS.n11 4.5005
R14600 VSS.n199 VSS.n11 4.5005
R14601 VSS.n188 VSS.n11 4.5005
R14602 VSS.n200 VSS.n11 4.5005
R14603 VSS.n187 VSS.n11 4.5005
R14604 VSS.n201 VSS.n11 4.5005
R14605 VSS.n186 VSS.n11 4.5005
R14606 VSS.n202 VSS.n11 4.5005
R14607 VSS.n185 VSS.n11 4.5005
R14608 VSS.n203 VSS.n11 4.5005
R14609 VSS.n184 VSS.n11 4.5005
R14610 VSS.n204 VSS.n11 4.5005
R14611 VSS.n183 VSS.n11 4.5005
R14612 VSS.n205 VSS.n11 4.5005
R14613 VSS.n182 VSS.n11 4.5005
R14614 VSS.n206 VSS.n11 4.5005
R14615 VSS.n181 VSS.n11 4.5005
R14616 VSS.n207 VSS.n11 4.5005
R14617 VSS.n180 VSS.n11 4.5005
R14618 VSS.n208 VSS.n11 4.5005
R14619 VSS.n179 VSS.n11 4.5005
R14620 VSS.n209 VSS.n11 4.5005
R14621 VSS.n178 VSS.n11 4.5005
R14622 VSS.n210 VSS.n11 4.5005
R14623 VSS.n177 VSS.n11 4.5005
R14624 VSS.n211 VSS.n11 4.5005
R14625 VSS.n176 VSS.n11 4.5005
R14626 VSS.n212 VSS.n11 4.5005
R14627 VSS.n175 VSS.n11 4.5005
R14628 VSS.n213 VSS.n11 4.5005
R14629 VSS.n174 VSS.n11 4.5005
R14630 VSS.n214 VSS.n11 4.5005
R14631 VSS.n173 VSS.n11 4.5005
R14632 VSS.n215 VSS.n11 4.5005
R14633 VSS.n172 VSS.n11 4.5005
R14634 VSS.n216 VSS.n11 4.5005
R14635 VSS.n171 VSS.n11 4.5005
R14636 VSS.n217 VSS.n11 4.5005
R14637 VSS.n170 VSS.n11 4.5005
R14638 VSS.n218 VSS.n11 4.5005
R14639 VSS.n169 VSS.n11 4.5005
R14640 VSS.n219 VSS.n11 4.5005
R14641 VSS.n168 VSS.n11 4.5005
R14642 VSS.n220 VSS.n11 4.5005
R14643 VSS.n167 VSS.n11 4.5005
R14644 VSS.n221 VSS.n11 4.5005
R14645 VSS.n166 VSS.n11 4.5005
R14646 VSS.n222 VSS.n11 4.5005
R14647 VSS.n165 VSS.n11 4.5005
R14648 VSS.n223 VSS.n11 4.5005
R14649 VSS.n164 VSS.n11 4.5005
R14650 VSS.n224 VSS.n11 4.5005
R14651 VSS.n163 VSS.n11 4.5005
R14652 VSS.n225 VSS.n11 4.5005
R14653 VSS.n162 VSS.n11 4.5005
R14654 VSS.n226 VSS.n11 4.5005
R14655 VSS.n161 VSS.n11 4.5005
R14656 VSS.n227 VSS.n11 4.5005
R14657 VSS.n160 VSS.n11 4.5005
R14658 VSS.n228 VSS.n11 4.5005
R14659 VSS.n159 VSS.n11 4.5005
R14660 VSS.n229 VSS.n11 4.5005
R14661 VSS.n158 VSS.n11 4.5005
R14662 VSS.n230 VSS.n11 4.5005
R14663 VSS.n157 VSS.n11 4.5005
R14664 VSS.n231 VSS.n11 4.5005
R14665 VSS.n156 VSS.n11 4.5005
R14666 VSS.n232 VSS.n11 4.5005
R14667 VSS.n155 VSS.n11 4.5005
R14668 VSS.n233 VSS.n11 4.5005
R14669 VSS.n154 VSS.n11 4.5005
R14670 VSS.n234 VSS.n11 4.5005
R14671 VSS.n153 VSS.n11 4.5005
R14672 VSS.n235 VSS.n11 4.5005
R14673 VSS.n4506 VSS.n11 4.5005
R14674 VSS.n236 VSS.n11 4.5005
R14675 VSS.n152 VSS.n11 4.5005
R14676 VSS.n237 VSS.n11 4.5005
R14677 VSS.n151 VSS.n11 4.5005
R14678 VSS.n238 VSS.n11 4.5005
R14679 VSS.n150 VSS.n11 4.5005
R14680 VSS.n239 VSS.n11 4.5005
R14681 VSS.n149 VSS.n11 4.5005
R14682 VSS.n240 VSS.n11 4.5005
R14683 VSS.n148 VSS.n11 4.5005
R14684 VSS.n241 VSS.n11 4.5005
R14685 VSS.n147 VSS.n11 4.5005
R14686 VSS.n242 VSS.n11 4.5005
R14687 VSS.n146 VSS.n11 4.5005
R14688 VSS.n243 VSS.n11 4.5005
R14689 VSS.n145 VSS.n11 4.5005
R14690 VSS.n244 VSS.n11 4.5005
R14691 VSS.n144 VSS.n11 4.5005
R14692 VSS.n245 VSS.n11 4.5005
R14693 VSS.n143 VSS.n11 4.5005
R14694 VSS.n246 VSS.n11 4.5005
R14695 VSS.n142 VSS.n11 4.5005
R14696 VSS.n247 VSS.n11 4.5005
R14697 VSS.n141 VSS.n11 4.5005
R14698 VSS.n248 VSS.n11 4.5005
R14699 VSS.n140 VSS.n11 4.5005
R14700 VSS.n249 VSS.n11 4.5005
R14701 VSS.n139 VSS.n11 4.5005
R14702 VSS.n250 VSS.n11 4.5005
R14703 VSS.n138 VSS.n11 4.5005
R14704 VSS.n251 VSS.n11 4.5005
R14705 VSS.n137 VSS.n11 4.5005
R14706 VSS.n252 VSS.n11 4.5005
R14707 VSS.n136 VSS.n11 4.5005
R14708 VSS.n253 VSS.n11 4.5005
R14709 VSS.n135 VSS.n11 4.5005
R14710 VSS.n254 VSS.n11 4.5005
R14711 VSS.n134 VSS.n11 4.5005
R14712 VSS.n255 VSS.n11 4.5005
R14713 VSS.n133 VSS.n11 4.5005
R14714 VSS.n256 VSS.n11 4.5005
R14715 VSS.n132 VSS.n11 4.5005
R14716 VSS.n4502 VSS.n11 4.5005
R14717 VSS.n4504 VSS.n11 4.5005
R14718 VSS.n193 VSS.n126 4.5005
R14719 VSS.n195 VSS.n126 4.5005
R14720 VSS.n192 VSS.n126 4.5005
R14721 VSS.n196 VSS.n126 4.5005
R14722 VSS.n191 VSS.n126 4.5005
R14723 VSS.n197 VSS.n126 4.5005
R14724 VSS.n190 VSS.n126 4.5005
R14725 VSS.n198 VSS.n126 4.5005
R14726 VSS.n189 VSS.n126 4.5005
R14727 VSS.n199 VSS.n126 4.5005
R14728 VSS.n188 VSS.n126 4.5005
R14729 VSS.n200 VSS.n126 4.5005
R14730 VSS.n187 VSS.n126 4.5005
R14731 VSS.n201 VSS.n126 4.5005
R14732 VSS.n186 VSS.n126 4.5005
R14733 VSS.n202 VSS.n126 4.5005
R14734 VSS.n185 VSS.n126 4.5005
R14735 VSS.n203 VSS.n126 4.5005
R14736 VSS.n184 VSS.n126 4.5005
R14737 VSS.n204 VSS.n126 4.5005
R14738 VSS.n183 VSS.n126 4.5005
R14739 VSS.n205 VSS.n126 4.5005
R14740 VSS.n182 VSS.n126 4.5005
R14741 VSS.n206 VSS.n126 4.5005
R14742 VSS.n181 VSS.n126 4.5005
R14743 VSS.n207 VSS.n126 4.5005
R14744 VSS.n180 VSS.n126 4.5005
R14745 VSS.n208 VSS.n126 4.5005
R14746 VSS.n179 VSS.n126 4.5005
R14747 VSS.n209 VSS.n126 4.5005
R14748 VSS.n178 VSS.n126 4.5005
R14749 VSS.n210 VSS.n126 4.5005
R14750 VSS.n177 VSS.n126 4.5005
R14751 VSS.n211 VSS.n126 4.5005
R14752 VSS.n176 VSS.n126 4.5005
R14753 VSS.n212 VSS.n126 4.5005
R14754 VSS.n175 VSS.n126 4.5005
R14755 VSS.n213 VSS.n126 4.5005
R14756 VSS.n174 VSS.n126 4.5005
R14757 VSS.n214 VSS.n126 4.5005
R14758 VSS.n173 VSS.n126 4.5005
R14759 VSS.n215 VSS.n126 4.5005
R14760 VSS.n172 VSS.n126 4.5005
R14761 VSS.n216 VSS.n126 4.5005
R14762 VSS.n171 VSS.n126 4.5005
R14763 VSS.n217 VSS.n126 4.5005
R14764 VSS.n170 VSS.n126 4.5005
R14765 VSS.n218 VSS.n126 4.5005
R14766 VSS.n169 VSS.n126 4.5005
R14767 VSS.n219 VSS.n126 4.5005
R14768 VSS.n168 VSS.n126 4.5005
R14769 VSS.n220 VSS.n126 4.5005
R14770 VSS.n167 VSS.n126 4.5005
R14771 VSS.n221 VSS.n126 4.5005
R14772 VSS.n166 VSS.n126 4.5005
R14773 VSS.n222 VSS.n126 4.5005
R14774 VSS.n165 VSS.n126 4.5005
R14775 VSS.n223 VSS.n126 4.5005
R14776 VSS.n164 VSS.n126 4.5005
R14777 VSS.n224 VSS.n126 4.5005
R14778 VSS.n163 VSS.n126 4.5005
R14779 VSS.n225 VSS.n126 4.5005
R14780 VSS.n162 VSS.n126 4.5005
R14781 VSS.n226 VSS.n126 4.5005
R14782 VSS.n161 VSS.n126 4.5005
R14783 VSS.n227 VSS.n126 4.5005
R14784 VSS.n160 VSS.n126 4.5005
R14785 VSS.n228 VSS.n126 4.5005
R14786 VSS.n159 VSS.n126 4.5005
R14787 VSS.n229 VSS.n126 4.5005
R14788 VSS.n158 VSS.n126 4.5005
R14789 VSS.n230 VSS.n126 4.5005
R14790 VSS.n157 VSS.n126 4.5005
R14791 VSS.n231 VSS.n126 4.5005
R14792 VSS.n156 VSS.n126 4.5005
R14793 VSS.n232 VSS.n126 4.5005
R14794 VSS.n155 VSS.n126 4.5005
R14795 VSS.n233 VSS.n126 4.5005
R14796 VSS.n154 VSS.n126 4.5005
R14797 VSS.n234 VSS.n126 4.5005
R14798 VSS.n153 VSS.n126 4.5005
R14799 VSS.n235 VSS.n126 4.5005
R14800 VSS.n4506 VSS.n126 4.5005
R14801 VSS.n236 VSS.n126 4.5005
R14802 VSS.n152 VSS.n126 4.5005
R14803 VSS.n237 VSS.n126 4.5005
R14804 VSS.n151 VSS.n126 4.5005
R14805 VSS.n238 VSS.n126 4.5005
R14806 VSS.n150 VSS.n126 4.5005
R14807 VSS.n239 VSS.n126 4.5005
R14808 VSS.n149 VSS.n126 4.5005
R14809 VSS.n240 VSS.n126 4.5005
R14810 VSS.n148 VSS.n126 4.5005
R14811 VSS.n241 VSS.n126 4.5005
R14812 VSS.n147 VSS.n126 4.5005
R14813 VSS.n242 VSS.n126 4.5005
R14814 VSS.n146 VSS.n126 4.5005
R14815 VSS.n243 VSS.n126 4.5005
R14816 VSS.n145 VSS.n126 4.5005
R14817 VSS.n244 VSS.n126 4.5005
R14818 VSS.n144 VSS.n126 4.5005
R14819 VSS.n245 VSS.n126 4.5005
R14820 VSS.n143 VSS.n126 4.5005
R14821 VSS.n246 VSS.n126 4.5005
R14822 VSS.n142 VSS.n126 4.5005
R14823 VSS.n247 VSS.n126 4.5005
R14824 VSS.n141 VSS.n126 4.5005
R14825 VSS.n248 VSS.n126 4.5005
R14826 VSS.n140 VSS.n126 4.5005
R14827 VSS.n249 VSS.n126 4.5005
R14828 VSS.n139 VSS.n126 4.5005
R14829 VSS.n250 VSS.n126 4.5005
R14830 VSS.n138 VSS.n126 4.5005
R14831 VSS.n251 VSS.n126 4.5005
R14832 VSS.n137 VSS.n126 4.5005
R14833 VSS.n252 VSS.n126 4.5005
R14834 VSS.n136 VSS.n126 4.5005
R14835 VSS.n253 VSS.n126 4.5005
R14836 VSS.n135 VSS.n126 4.5005
R14837 VSS.n254 VSS.n126 4.5005
R14838 VSS.n134 VSS.n126 4.5005
R14839 VSS.n255 VSS.n126 4.5005
R14840 VSS.n133 VSS.n126 4.5005
R14841 VSS.n256 VSS.n126 4.5005
R14842 VSS.n132 VSS.n126 4.5005
R14843 VSS.n4502 VSS.n126 4.5005
R14844 VSS.n4504 VSS.n126 4.5005
R14845 VSS.n193 VSS.n10 4.5005
R14846 VSS.n195 VSS.n10 4.5005
R14847 VSS.n192 VSS.n10 4.5005
R14848 VSS.n196 VSS.n10 4.5005
R14849 VSS.n191 VSS.n10 4.5005
R14850 VSS.n197 VSS.n10 4.5005
R14851 VSS.n190 VSS.n10 4.5005
R14852 VSS.n198 VSS.n10 4.5005
R14853 VSS.n189 VSS.n10 4.5005
R14854 VSS.n199 VSS.n10 4.5005
R14855 VSS.n188 VSS.n10 4.5005
R14856 VSS.n200 VSS.n10 4.5005
R14857 VSS.n187 VSS.n10 4.5005
R14858 VSS.n201 VSS.n10 4.5005
R14859 VSS.n186 VSS.n10 4.5005
R14860 VSS.n202 VSS.n10 4.5005
R14861 VSS.n185 VSS.n10 4.5005
R14862 VSS.n203 VSS.n10 4.5005
R14863 VSS.n184 VSS.n10 4.5005
R14864 VSS.n204 VSS.n10 4.5005
R14865 VSS.n183 VSS.n10 4.5005
R14866 VSS.n205 VSS.n10 4.5005
R14867 VSS.n182 VSS.n10 4.5005
R14868 VSS.n206 VSS.n10 4.5005
R14869 VSS.n181 VSS.n10 4.5005
R14870 VSS.n207 VSS.n10 4.5005
R14871 VSS.n180 VSS.n10 4.5005
R14872 VSS.n208 VSS.n10 4.5005
R14873 VSS.n179 VSS.n10 4.5005
R14874 VSS.n209 VSS.n10 4.5005
R14875 VSS.n178 VSS.n10 4.5005
R14876 VSS.n210 VSS.n10 4.5005
R14877 VSS.n177 VSS.n10 4.5005
R14878 VSS.n211 VSS.n10 4.5005
R14879 VSS.n176 VSS.n10 4.5005
R14880 VSS.n212 VSS.n10 4.5005
R14881 VSS.n175 VSS.n10 4.5005
R14882 VSS.n213 VSS.n10 4.5005
R14883 VSS.n174 VSS.n10 4.5005
R14884 VSS.n214 VSS.n10 4.5005
R14885 VSS.n173 VSS.n10 4.5005
R14886 VSS.n215 VSS.n10 4.5005
R14887 VSS.n172 VSS.n10 4.5005
R14888 VSS.n216 VSS.n10 4.5005
R14889 VSS.n171 VSS.n10 4.5005
R14890 VSS.n217 VSS.n10 4.5005
R14891 VSS.n170 VSS.n10 4.5005
R14892 VSS.n218 VSS.n10 4.5005
R14893 VSS.n169 VSS.n10 4.5005
R14894 VSS.n219 VSS.n10 4.5005
R14895 VSS.n168 VSS.n10 4.5005
R14896 VSS.n220 VSS.n10 4.5005
R14897 VSS.n167 VSS.n10 4.5005
R14898 VSS.n221 VSS.n10 4.5005
R14899 VSS.n166 VSS.n10 4.5005
R14900 VSS.n222 VSS.n10 4.5005
R14901 VSS.n165 VSS.n10 4.5005
R14902 VSS.n223 VSS.n10 4.5005
R14903 VSS.n164 VSS.n10 4.5005
R14904 VSS.n224 VSS.n10 4.5005
R14905 VSS.n163 VSS.n10 4.5005
R14906 VSS.n225 VSS.n10 4.5005
R14907 VSS.n162 VSS.n10 4.5005
R14908 VSS.n226 VSS.n10 4.5005
R14909 VSS.n161 VSS.n10 4.5005
R14910 VSS.n227 VSS.n10 4.5005
R14911 VSS.n160 VSS.n10 4.5005
R14912 VSS.n228 VSS.n10 4.5005
R14913 VSS.n159 VSS.n10 4.5005
R14914 VSS.n229 VSS.n10 4.5005
R14915 VSS.n158 VSS.n10 4.5005
R14916 VSS.n230 VSS.n10 4.5005
R14917 VSS.n157 VSS.n10 4.5005
R14918 VSS.n231 VSS.n10 4.5005
R14919 VSS.n156 VSS.n10 4.5005
R14920 VSS.n232 VSS.n10 4.5005
R14921 VSS.n155 VSS.n10 4.5005
R14922 VSS.n233 VSS.n10 4.5005
R14923 VSS.n154 VSS.n10 4.5005
R14924 VSS.n234 VSS.n10 4.5005
R14925 VSS.n153 VSS.n10 4.5005
R14926 VSS.n235 VSS.n10 4.5005
R14927 VSS.n4506 VSS.n10 4.5005
R14928 VSS.n236 VSS.n10 4.5005
R14929 VSS.n152 VSS.n10 4.5005
R14930 VSS.n237 VSS.n10 4.5005
R14931 VSS.n151 VSS.n10 4.5005
R14932 VSS.n238 VSS.n10 4.5005
R14933 VSS.n150 VSS.n10 4.5005
R14934 VSS.n239 VSS.n10 4.5005
R14935 VSS.n149 VSS.n10 4.5005
R14936 VSS.n240 VSS.n10 4.5005
R14937 VSS.n148 VSS.n10 4.5005
R14938 VSS.n241 VSS.n10 4.5005
R14939 VSS.n147 VSS.n10 4.5005
R14940 VSS.n242 VSS.n10 4.5005
R14941 VSS.n146 VSS.n10 4.5005
R14942 VSS.n243 VSS.n10 4.5005
R14943 VSS.n145 VSS.n10 4.5005
R14944 VSS.n244 VSS.n10 4.5005
R14945 VSS.n144 VSS.n10 4.5005
R14946 VSS.n245 VSS.n10 4.5005
R14947 VSS.n143 VSS.n10 4.5005
R14948 VSS.n246 VSS.n10 4.5005
R14949 VSS.n142 VSS.n10 4.5005
R14950 VSS.n247 VSS.n10 4.5005
R14951 VSS.n141 VSS.n10 4.5005
R14952 VSS.n248 VSS.n10 4.5005
R14953 VSS.n140 VSS.n10 4.5005
R14954 VSS.n249 VSS.n10 4.5005
R14955 VSS.n139 VSS.n10 4.5005
R14956 VSS.n250 VSS.n10 4.5005
R14957 VSS.n138 VSS.n10 4.5005
R14958 VSS.n251 VSS.n10 4.5005
R14959 VSS.n137 VSS.n10 4.5005
R14960 VSS.n252 VSS.n10 4.5005
R14961 VSS.n136 VSS.n10 4.5005
R14962 VSS.n253 VSS.n10 4.5005
R14963 VSS.n135 VSS.n10 4.5005
R14964 VSS.n254 VSS.n10 4.5005
R14965 VSS.n134 VSS.n10 4.5005
R14966 VSS.n255 VSS.n10 4.5005
R14967 VSS.n133 VSS.n10 4.5005
R14968 VSS.n256 VSS.n10 4.5005
R14969 VSS.n132 VSS.n10 4.5005
R14970 VSS.n4502 VSS.n10 4.5005
R14971 VSS.n4504 VSS.n10 4.5005
R14972 VSS.n193 VSS.n127 4.5005
R14973 VSS.n195 VSS.n127 4.5005
R14974 VSS.n192 VSS.n127 4.5005
R14975 VSS.n196 VSS.n127 4.5005
R14976 VSS.n191 VSS.n127 4.5005
R14977 VSS.n197 VSS.n127 4.5005
R14978 VSS.n190 VSS.n127 4.5005
R14979 VSS.n198 VSS.n127 4.5005
R14980 VSS.n189 VSS.n127 4.5005
R14981 VSS.n199 VSS.n127 4.5005
R14982 VSS.n188 VSS.n127 4.5005
R14983 VSS.n200 VSS.n127 4.5005
R14984 VSS.n187 VSS.n127 4.5005
R14985 VSS.n201 VSS.n127 4.5005
R14986 VSS.n186 VSS.n127 4.5005
R14987 VSS.n202 VSS.n127 4.5005
R14988 VSS.n185 VSS.n127 4.5005
R14989 VSS.n203 VSS.n127 4.5005
R14990 VSS.n184 VSS.n127 4.5005
R14991 VSS.n204 VSS.n127 4.5005
R14992 VSS.n183 VSS.n127 4.5005
R14993 VSS.n205 VSS.n127 4.5005
R14994 VSS.n182 VSS.n127 4.5005
R14995 VSS.n206 VSS.n127 4.5005
R14996 VSS.n181 VSS.n127 4.5005
R14997 VSS.n207 VSS.n127 4.5005
R14998 VSS.n180 VSS.n127 4.5005
R14999 VSS.n208 VSS.n127 4.5005
R15000 VSS.n179 VSS.n127 4.5005
R15001 VSS.n209 VSS.n127 4.5005
R15002 VSS.n178 VSS.n127 4.5005
R15003 VSS.n210 VSS.n127 4.5005
R15004 VSS.n177 VSS.n127 4.5005
R15005 VSS.n211 VSS.n127 4.5005
R15006 VSS.n176 VSS.n127 4.5005
R15007 VSS.n212 VSS.n127 4.5005
R15008 VSS.n175 VSS.n127 4.5005
R15009 VSS.n213 VSS.n127 4.5005
R15010 VSS.n174 VSS.n127 4.5005
R15011 VSS.n214 VSS.n127 4.5005
R15012 VSS.n173 VSS.n127 4.5005
R15013 VSS.n215 VSS.n127 4.5005
R15014 VSS.n172 VSS.n127 4.5005
R15015 VSS.n216 VSS.n127 4.5005
R15016 VSS.n171 VSS.n127 4.5005
R15017 VSS.n217 VSS.n127 4.5005
R15018 VSS.n170 VSS.n127 4.5005
R15019 VSS.n218 VSS.n127 4.5005
R15020 VSS.n169 VSS.n127 4.5005
R15021 VSS.n219 VSS.n127 4.5005
R15022 VSS.n168 VSS.n127 4.5005
R15023 VSS.n220 VSS.n127 4.5005
R15024 VSS.n167 VSS.n127 4.5005
R15025 VSS.n221 VSS.n127 4.5005
R15026 VSS.n166 VSS.n127 4.5005
R15027 VSS.n222 VSS.n127 4.5005
R15028 VSS.n165 VSS.n127 4.5005
R15029 VSS.n223 VSS.n127 4.5005
R15030 VSS.n164 VSS.n127 4.5005
R15031 VSS.n224 VSS.n127 4.5005
R15032 VSS.n163 VSS.n127 4.5005
R15033 VSS.n225 VSS.n127 4.5005
R15034 VSS.n162 VSS.n127 4.5005
R15035 VSS.n226 VSS.n127 4.5005
R15036 VSS.n161 VSS.n127 4.5005
R15037 VSS.n227 VSS.n127 4.5005
R15038 VSS.n160 VSS.n127 4.5005
R15039 VSS.n228 VSS.n127 4.5005
R15040 VSS.n159 VSS.n127 4.5005
R15041 VSS.n229 VSS.n127 4.5005
R15042 VSS.n158 VSS.n127 4.5005
R15043 VSS.n230 VSS.n127 4.5005
R15044 VSS.n157 VSS.n127 4.5005
R15045 VSS.n231 VSS.n127 4.5005
R15046 VSS.n156 VSS.n127 4.5005
R15047 VSS.n232 VSS.n127 4.5005
R15048 VSS.n155 VSS.n127 4.5005
R15049 VSS.n233 VSS.n127 4.5005
R15050 VSS.n154 VSS.n127 4.5005
R15051 VSS.n234 VSS.n127 4.5005
R15052 VSS.n153 VSS.n127 4.5005
R15053 VSS.n235 VSS.n127 4.5005
R15054 VSS.n4506 VSS.n127 4.5005
R15055 VSS.n236 VSS.n127 4.5005
R15056 VSS.n152 VSS.n127 4.5005
R15057 VSS.n237 VSS.n127 4.5005
R15058 VSS.n151 VSS.n127 4.5005
R15059 VSS.n238 VSS.n127 4.5005
R15060 VSS.n150 VSS.n127 4.5005
R15061 VSS.n239 VSS.n127 4.5005
R15062 VSS.n149 VSS.n127 4.5005
R15063 VSS.n240 VSS.n127 4.5005
R15064 VSS.n148 VSS.n127 4.5005
R15065 VSS.n241 VSS.n127 4.5005
R15066 VSS.n147 VSS.n127 4.5005
R15067 VSS.n242 VSS.n127 4.5005
R15068 VSS.n146 VSS.n127 4.5005
R15069 VSS.n243 VSS.n127 4.5005
R15070 VSS.n145 VSS.n127 4.5005
R15071 VSS.n244 VSS.n127 4.5005
R15072 VSS.n144 VSS.n127 4.5005
R15073 VSS.n245 VSS.n127 4.5005
R15074 VSS.n143 VSS.n127 4.5005
R15075 VSS.n246 VSS.n127 4.5005
R15076 VSS.n142 VSS.n127 4.5005
R15077 VSS.n247 VSS.n127 4.5005
R15078 VSS.n141 VSS.n127 4.5005
R15079 VSS.n248 VSS.n127 4.5005
R15080 VSS.n140 VSS.n127 4.5005
R15081 VSS.n249 VSS.n127 4.5005
R15082 VSS.n139 VSS.n127 4.5005
R15083 VSS.n250 VSS.n127 4.5005
R15084 VSS.n138 VSS.n127 4.5005
R15085 VSS.n251 VSS.n127 4.5005
R15086 VSS.n137 VSS.n127 4.5005
R15087 VSS.n252 VSS.n127 4.5005
R15088 VSS.n136 VSS.n127 4.5005
R15089 VSS.n253 VSS.n127 4.5005
R15090 VSS.n135 VSS.n127 4.5005
R15091 VSS.n254 VSS.n127 4.5005
R15092 VSS.n134 VSS.n127 4.5005
R15093 VSS.n255 VSS.n127 4.5005
R15094 VSS.n133 VSS.n127 4.5005
R15095 VSS.n256 VSS.n127 4.5005
R15096 VSS.n132 VSS.n127 4.5005
R15097 VSS.n4502 VSS.n127 4.5005
R15098 VSS.n4504 VSS.n127 4.5005
R15099 VSS.n193 VSS.n9 4.5005
R15100 VSS.n195 VSS.n9 4.5005
R15101 VSS.n192 VSS.n9 4.5005
R15102 VSS.n196 VSS.n9 4.5005
R15103 VSS.n191 VSS.n9 4.5005
R15104 VSS.n197 VSS.n9 4.5005
R15105 VSS.n190 VSS.n9 4.5005
R15106 VSS.n198 VSS.n9 4.5005
R15107 VSS.n189 VSS.n9 4.5005
R15108 VSS.n199 VSS.n9 4.5005
R15109 VSS.n188 VSS.n9 4.5005
R15110 VSS.n200 VSS.n9 4.5005
R15111 VSS.n187 VSS.n9 4.5005
R15112 VSS.n201 VSS.n9 4.5005
R15113 VSS.n186 VSS.n9 4.5005
R15114 VSS.n202 VSS.n9 4.5005
R15115 VSS.n185 VSS.n9 4.5005
R15116 VSS.n203 VSS.n9 4.5005
R15117 VSS.n184 VSS.n9 4.5005
R15118 VSS.n204 VSS.n9 4.5005
R15119 VSS.n183 VSS.n9 4.5005
R15120 VSS.n205 VSS.n9 4.5005
R15121 VSS.n182 VSS.n9 4.5005
R15122 VSS.n206 VSS.n9 4.5005
R15123 VSS.n181 VSS.n9 4.5005
R15124 VSS.n207 VSS.n9 4.5005
R15125 VSS.n180 VSS.n9 4.5005
R15126 VSS.n208 VSS.n9 4.5005
R15127 VSS.n179 VSS.n9 4.5005
R15128 VSS.n209 VSS.n9 4.5005
R15129 VSS.n178 VSS.n9 4.5005
R15130 VSS.n210 VSS.n9 4.5005
R15131 VSS.n177 VSS.n9 4.5005
R15132 VSS.n211 VSS.n9 4.5005
R15133 VSS.n176 VSS.n9 4.5005
R15134 VSS.n212 VSS.n9 4.5005
R15135 VSS.n175 VSS.n9 4.5005
R15136 VSS.n213 VSS.n9 4.5005
R15137 VSS.n174 VSS.n9 4.5005
R15138 VSS.n214 VSS.n9 4.5005
R15139 VSS.n173 VSS.n9 4.5005
R15140 VSS.n215 VSS.n9 4.5005
R15141 VSS.n172 VSS.n9 4.5005
R15142 VSS.n216 VSS.n9 4.5005
R15143 VSS.n171 VSS.n9 4.5005
R15144 VSS.n217 VSS.n9 4.5005
R15145 VSS.n170 VSS.n9 4.5005
R15146 VSS.n218 VSS.n9 4.5005
R15147 VSS.n169 VSS.n9 4.5005
R15148 VSS.n219 VSS.n9 4.5005
R15149 VSS.n168 VSS.n9 4.5005
R15150 VSS.n220 VSS.n9 4.5005
R15151 VSS.n167 VSS.n9 4.5005
R15152 VSS.n221 VSS.n9 4.5005
R15153 VSS.n166 VSS.n9 4.5005
R15154 VSS.n222 VSS.n9 4.5005
R15155 VSS.n165 VSS.n9 4.5005
R15156 VSS.n223 VSS.n9 4.5005
R15157 VSS.n164 VSS.n9 4.5005
R15158 VSS.n224 VSS.n9 4.5005
R15159 VSS.n163 VSS.n9 4.5005
R15160 VSS.n225 VSS.n9 4.5005
R15161 VSS.n162 VSS.n9 4.5005
R15162 VSS.n226 VSS.n9 4.5005
R15163 VSS.n161 VSS.n9 4.5005
R15164 VSS.n227 VSS.n9 4.5005
R15165 VSS.n160 VSS.n9 4.5005
R15166 VSS.n228 VSS.n9 4.5005
R15167 VSS.n159 VSS.n9 4.5005
R15168 VSS.n229 VSS.n9 4.5005
R15169 VSS.n158 VSS.n9 4.5005
R15170 VSS.n230 VSS.n9 4.5005
R15171 VSS.n157 VSS.n9 4.5005
R15172 VSS.n231 VSS.n9 4.5005
R15173 VSS.n156 VSS.n9 4.5005
R15174 VSS.n232 VSS.n9 4.5005
R15175 VSS.n155 VSS.n9 4.5005
R15176 VSS.n233 VSS.n9 4.5005
R15177 VSS.n154 VSS.n9 4.5005
R15178 VSS.n234 VSS.n9 4.5005
R15179 VSS.n153 VSS.n9 4.5005
R15180 VSS.n235 VSS.n9 4.5005
R15181 VSS.n4506 VSS.n9 4.5005
R15182 VSS.n236 VSS.n9 4.5005
R15183 VSS.n152 VSS.n9 4.5005
R15184 VSS.n237 VSS.n9 4.5005
R15185 VSS.n151 VSS.n9 4.5005
R15186 VSS.n238 VSS.n9 4.5005
R15187 VSS.n150 VSS.n9 4.5005
R15188 VSS.n239 VSS.n9 4.5005
R15189 VSS.n149 VSS.n9 4.5005
R15190 VSS.n240 VSS.n9 4.5005
R15191 VSS.n148 VSS.n9 4.5005
R15192 VSS.n241 VSS.n9 4.5005
R15193 VSS.n147 VSS.n9 4.5005
R15194 VSS.n242 VSS.n9 4.5005
R15195 VSS.n146 VSS.n9 4.5005
R15196 VSS.n243 VSS.n9 4.5005
R15197 VSS.n145 VSS.n9 4.5005
R15198 VSS.n244 VSS.n9 4.5005
R15199 VSS.n144 VSS.n9 4.5005
R15200 VSS.n245 VSS.n9 4.5005
R15201 VSS.n143 VSS.n9 4.5005
R15202 VSS.n246 VSS.n9 4.5005
R15203 VSS.n142 VSS.n9 4.5005
R15204 VSS.n247 VSS.n9 4.5005
R15205 VSS.n141 VSS.n9 4.5005
R15206 VSS.n248 VSS.n9 4.5005
R15207 VSS.n140 VSS.n9 4.5005
R15208 VSS.n249 VSS.n9 4.5005
R15209 VSS.n139 VSS.n9 4.5005
R15210 VSS.n250 VSS.n9 4.5005
R15211 VSS.n138 VSS.n9 4.5005
R15212 VSS.n251 VSS.n9 4.5005
R15213 VSS.n137 VSS.n9 4.5005
R15214 VSS.n252 VSS.n9 4.5005
R15215 VSS.n136 VSS.n9 4.5005
R15216 VSS.n253 VSS.n9 4.5005
R15217 VSS.n135 VSS.n9 4.5005
R15218 VSS.n254 VSS.n9 4.5005
R15219 VSS.n134 VSS.n9 4.5005
R15220 VSS.n255 VSS.n9 4.5005
R15221 VSS.n133 VSS.n9 4.5005
R15222 VSS.n256 VSS.n9 4.5005
R15223 VSS.n132 VSS.n9 4.5005
R15224 VSS.n4502 VSS.n9 4.5005
R15225 VSS.n4504 VSS.n9 4.5005
R15226 VSS.n193 VSS.n128 4.5005
R15227 VSS.n195 VSS.n128 4.5005
R15228 VSS.n192 VSS.n128 4.5005
R15229 VSS.n196 VSS.n128 4.5005
R15230 VSS.n191 VSS.n128 4.5005
R15231 VSS.n197 VSS.n128 4.5005
R15232 VSS.n190 VSS.n128 4.5005
R15233 VSS.n198 VSS.n128 4.5005
R15234 VSS.n189 VSS.n128 4.5005
R15235 VSS.n199 VSS.n128 4.5005
R15236 VSS.n188 VSS.n128 4.5005
R15237 VSS.n200 VSS.n128 4.5005
R15238 VSS.n187 VSS.n128 4.5005
R15239 VSS.n201 VSS.n128 4.5005
R15240 VSS.n186 VSS.n128 4.5005
R15241 VSS.n202 VSS.n128 4.5005
R15242 VSS.n185 VSS.n128 4.5005
R15243 VSS.n203 VSS.n128 4.5005
R15244 VSS.n184 VSS.n128 4.5005
R15245 VSS.n204 VSS.n128 4.5005
R15246 VSS.n183 VSS.n128 4.5005
R15247 VSS.n205 VSS.n128 4.5005
R15248 VSS.n182 VSS.n128 4.5005
R15249 VSS.n206 VSS.n128 4.5005
R15250 VSS.n181 VSS.n128 4.5005
R15251 VSS.n207 VSS.n128 4.5005
R15252 VSS.n180 VSS.n128 4.5005
R15253 VSS.n208 VSS.n128 4.5005
R15254 VSS.n179 VSS.n128 4.5005
R15255 VSS.n209 VSS.n128 4.5005
R15256 VSS.n178 VSS.n128 4.5005
R15257 VSS.n210 VSS.n128 4.5005
R15258 VSS.n177 VSS.n128 4.5005
R15259 VSS.n211 VSS.n128 4.5005
R15260 VSS.n176 VSS.n128 4.5005
R15261 VSS.n212 VSS.n128 4.5005
R15262 VSS.n175 VSS.n128 4.5005
R15263 VSS.n213 VSS.n128 4.5005
R15264 VSS.n174 VSS.n128 4.5005
R15265 VSS.n214 VSS.n128 4.5005
R15266 VSS.n173 VSS.n128 4.5005
R15267 VSS.n215 VSS.n128 4.5005
R15268 VSS.n172 VSS.n128 4.5005
R15269 VSS.n216 VSS.n128 4.5005
R15270 VSS.n171 VSS.n128 4.5005
R15271 VSS.n217 VSS.n128 4.5005
R15272 VSS.n170 VSS.n128 4.5005
R15273 VSS.n218 VSS.n128 4.5005
R15274 VSS.n169 VSS.n128 4.5005
R15275 VSS.n219 VSS.n128 4.5005
R15276 VSS.n168 VSS.n128 4.5005
R15277 VSS.n220 VSS.n128 4.5005
R15278 VSS.n167 VSS.n128 4.5005
R15279 VSS.n221 VSS.n128 4.5005
R15280 VSS.n166 VSS.n128 4.5005
R15281 VSS.n222 VSS.n128 4.5005
R15282 VSS.n165 VSS.n128 4.5005
R15283 VSS.n223 VSS.n128 4.5005
R15284 VSS.n164 VSS.n128 4.5005
R15285 VSS.n224 VSS.n128 4.5005
R15286 VSS.n163 VSS.n128 4.5005
R15287 VSS.n225 VSS.n128 4.5005
R15288 VSS.n162 VSS.n128 4.5005
R15289 VSS.n226 VSS.n128 4.5005
R15290 VSS.n161 VSS.n128 4.5005
R15291 VSS.n227 VSS.n128 4.5005
R15292 VSS.n160 VSS.n128 4.5005
R15293 VSS.n228 VSS.n128 4.5005
R15294 VSS.n159 VSS.n128 4.5005
R15295 VSS.n229 VSS.n128 4.5005
R15296 VSS.n158 VSS.n128 4.5005
R15297 VSS.n230 VSS.n128 4.5005
R15298 VSS.n157 VSS.n128 4.5005
R15299 VSS.n231 VSS.n128 4.5005
R15300 VSS.n156 VSS.n128 4.5005
R15301 VSS.n232 VSS.n128 4.5005
R15302 VSS.n155 VSS.n128 4.5005
R15303 VSS.n233 VSS.n128 4.5005
R15304 VSS.n154 VSS.n128 4.5005
R15305 VSS.n234 VSS.n128 4.5005
R15306 VSS.n153 VSS.n128 4.5005
R15307 VSS.n235 VSS.n128 4.5005
R15308 VSS.n4506 VSS.n128 4.5005
R15309 VSS.n236 VSS.n128 4.5005
R15310 VSS.n152 VSS.n128 4.5005
R15311 VSS.n237 VSS.n128 4.5005
R15312 VSS.n151 VSS.n128 4.5005
R15313 VSS.n238 VSS.n128 4.5005
R15314 VSS.n150 VSS.n128 4.5005
R15315 VSS.n239 VSS.n128 4.5005
R15316 VSS.n149 VSS.n128 4.5005
R15317 VSS.n240 VSS.n128 4.5005
R15318 VSS.n148 VSS.n128 4.5005
R15319 VSS.n241 VSS.n128 4.5005
R15320 VSS.n147 VSS.n128 4.5005
R15321 VSS.n242 VSS.n128 4.5005
R15322 VSS.n146 VSS.n128 4.5005
R15323 VSS.n243 VSS.n128 4.5005
R15324 VSS.n145 VSS.n128 4.5005
R15325 VSS.n244 VSS.n128 4.5005
R15326 VSS.n144 VSS.n128 4.5005
R15327 VSS.n245 VSS.n128 4.5005
R15328 VSS.n143 VSS.n128 4.5005
R15329 VSS.n246 VSS.n128 4.5005
R15330 VSS.n142 VSS.n128 4.5005
R15331 VSS.n247 VSS.n128 4.5005
R15332 VSS.n141 VSS.n128 4.5005
R15333 VSS.n248 VSS.n128 4.5005
R15334 VSS.n140 VSS.n128 4.5005
R15335 VSS.n249 VSS.n128 4.5005
R15336 VSS.n139 VSS.n128 4.5005
R15337 VSS.n250 VSS.n128 4.5005
R15338 VSS.n138 VSS.n128 4.5005
R15339 VSS.n251 VSS.n128 4.5005
R15340 VSS.n137 VSS.n128 4.5005
R15341 VSS.n252 VSS.n128 4.5005
R15342 VSS.n136 VSS.n128 4.5005
R15343 VSS.n253 VSS.n128 4.5005
R15344 VSS.n135 VSS.n128 4.5005
R15345 VSS.n254 VSS.n128 4.5005
R15346 VSS.n134 VSS.n128 4.5005
R15347 VSS.n255 VSS.n128 4.5005
R15348 VSS.n133 VSS.n128 4.5005
R15349 VSS.n256 VSS.n128 4.5005
R15350 VSS.n132 VSS.n128 4.5005
R15351 VSS.n4502 VSS.n128 4.5005
R15352 VSS.n4504 VSS.n128 4.5005
R15353 VSS.n193 VSS.n8 4.5005
R15354 VSS.n195 VSS.n8 4.5005
R15355 VSS.n192 VSS.n8 4.5005
R15356 VSS.n196 VSS.n8 4.5005
R15357 VSS.n191 VSS.n8 4.5005
R15358 VSS.n197 VSS.n8 4.5005
R15359 VSS.n190 VSS.n8 4.5005
R15360 VSS.n198 VSS.n8 4.5005
R15361 VSS.n189 VSS.n8 4.5005
R15362 VSS.n199 VSS.n8 4.5005
R15363 VSS.n188 VSS.n8 4.5005
R15364 VSS.n200 VSS.n8 4.5005
R15365 VSS.n187 VSS.n8 4.5005
R15366 VSS.n201 VSS.n8 4.5005
R15367 VSS.n186 VSS.n8 4.5005
R15368 VSS.n202 VSS.n8 4.5005
R15369 VSS.n185 VSS.n8 4.5005
R15370 VSS.n203 VSS.n8 4.5005
R15371 VSS.n184 VSS.n8 4.5005
R15372 VSS.n204 VSS.n8 4.5005
R15373 VSS.n183 VSS.n8 4.5005
R15374 VSS.n205 VSS.n8 4.5005
R15375 VSS.n182 VSS.n8 4.5005
R15376 VSS.n206 VSS.n8 4.5005
R15377 VSS.n181 VSS.n8 4.5005
R15378 VSS.n207 VSS.n8 4.5005
R15379 VSS.n180 VSS.n8 4.5005
R15380 VSS.n208 VSS.n8 4.5005
R15381 VSS.n179 VSS.n8 4.5005
R15382 VSS.n209 VSS.n8 4.5005
R15383 VSS.n178 VSS.n8 4.5005
R15384 VSS.n210 VSS.n8 4.5005
R15385 VSS.n177 VSS.n8 4.5005
R15386 VSS.n211 VSS.n8 4.5005
R15387 VSS.n176 VSS.n8 4.5005
R15388 VSS.n212 VSS.n8 4.5005
R15389 VSS.n175 VSS.n8 4.5005
R15390 VSS.n213 VSS.n8 4.5005
R15391 VSS.n174 VSS.n8 4.5005
R15392 VSS.n214 VSS.n8 4.5005
R15393 VSS.n173 VSS.n8 4.5005
R15394 VSS.n215 VSS.n8 4.5005
R15395 VSS.n172 VSS.n8 4.5005
R15396 VSS.n216 VSS.n8 4.5005
R15397 VSS.n171 VSS.n8 4.5005
R15398 VSS.n217 VSS.n8 4.5005
R15399 VSS.n170 VSS.n8 4.5005
R15400 VSS.n218 VSS.n8 4.5005
R15401 VSS.n169 VSS.n8 4.5005
R15402 VSS.n219 VSS.n8 4.5005
R15403 VSS.n168 VSS.n8 4.5005
R15404 VSS.n220 VSS.n8 4.5005
R15405 VSS.n167 VSS.n8 4.5005
R15406 VSS.n221 VSS.n8 4.5005
R15407 VSS.n166 VSS.n8 4.5005
R15408 VSS.n222 VSS.n8 4.5005
R15409 VSS.n165 VSS.n8 4.5005
R15410 VSS.n223 VSS.n8 4.5005
R15411 VSS.n164 VSS.n8 4.5005
R15412 VSS.n224 VSS.n8 4.5005
R15413 VSS.n163 VSS.n8 4.5005
R15414 VSS.n225 VSS.n8 4.5005
R15415 VSS.n162 VSS.n8 4.5005
R15416 VSS.n226 VSS.n8 4.5005
R15417 VSS.n161 VSS.n8 4.5005
R15418 VSS.n227 VSS.n8 4.5005
R15419 VSS.n160 VSS.n8 4.5005
R15420 VSS.n228 VSS.n8 4.5005
R15421 VSS.n159 VSS.n8 4.5005
R15422 VSS.n229 VSS.n8 4.5005
R15423 VSS.n158 VSS.n8 4.5005
R15424 VSS.n230 VSS.n8 4.5005
R15425 VSS.n157 VSS.n8 4.5005
R15426 VSS.n231 VSS.n8 4.5005
R15427 VSS.n156 VSS.n8 4.5005
R15428 VSS.n232 VSS.n8 4.5005
R15429 VSS.n155 VSS.n8 4.5005
R15430 VSS.n233 VSS.n8 4.5005
R15431 VSS.n154 VSS.n8 4.5005
R15432 VSS.n234 VSS.n8 4.5005
R15433 VSS.n153 VSS.n8 4.5005
R15434 VSS.n235 VSS.n8 4.5005
R15435 VSS.n4506 VSS.n8 4.5005
R15436 VSS.n236 VSS.n8 4.5005
R15437 VSS.n152 VSS.n8 4.5005
R15438 VSS.n237 VSS.n8 4.5005
R15439 VSS.n151 VSS.n8 4.5005
R15440 VSS.n238 VSS.n8 4.5005
R15441 VSS.n150 VSS.n8 4.5005
R15442 VSS.n239 VSS.n8 4.5005
R15443 VSS.n149 VSS.n8 4.5005
R15444 VSS.n240 VSS.n8 4.5005
R15445 VSS.n148 VSS.n8 4.5005
R15446 VSS.n241 VSS.n8 4.5005
R15447 VSS.n147 VSS.n8 4.5005
R15448 VSS.n242 VSS.n8 4.5005
R15449 VSS.n146 VSS.n8 4.5005
R15450 VSS.n243 VSS.n8 4.5005
R15451 VSS.n145 VSS.n8 4.5005
R15452 VSS.n244 VSS.n8 4.5005
R15453 VSS.n144 VSS.n8 4.5005
R15454 VSS.n245 VSS.n8 4.5005
R15455 VSS.n143 VSS.n8 4.5005
R15456 VSS.n246 VSS.n8 4.5005
R15457 VSS.n142 VSS.n8 4.5005
R15458 VSS.n247 VSS.n8 4.5005
R15459 VSS.n141 VSS.n8 4.5005
R15460 VSS.n248 VSS.n8 4.5005
R15461 VSS.n140 VSS.n8 4.5005
R15462 VSS.n249 VSS.n8 4.5005
R15463 VSS.n139 VSS.n8 4.5005
R15464 VSS.n250 VSS.n8 4.5005
R15465 VSS.n138 VSS.n8 4.5005
R15466 VSS.n251 VSS.n8 4.5005
R15467 VSS.n137 VSS.n8 4.5005
R15468 VSS.n252 VSS.n8 4.5005
R15469 VSS.n136 VSS.n8 4.5005
R15470 VSS.n253 VSS.n8 4.5005
R15471 VSS.n135 VSS.n8 4.5005
R15472 VSS.n254 VSS.n8 4.5005
R15473 VSS.n134 VSS.n8 4.5005
R15474 VSS.n255 VSS.n8 4.5005
R15475 VSS.n133 VSS.n8 4.5005
R15476 VSS.n256 VSS.n8 4.5005
R15477 VSS.n132 VSS.n8 4.5005
R15478 VSS.n4502 VSS.n8 4.5005
R15479 VSS.n4504 VSS.n8 4.5005
R15480 VSS.n193 VSS.n129 4.5005
R15481 VSS.n195 VSS.n129 4.5005
R15482 VSS.n192 VSS.n129 4.5005
R15483 VSS.n196 VSS.n129 4.5005
R15484 VSS.n191 VSS.n129 4.5005
R15485 VSS.n197 VSS.n129 4.5005
R15486 VSS.n190 VSS.n129 4.5005
R15487 VSS.n198 VSS.n129 4.5005
R15488 VSS.n189 VSS.n129 4.5005
R15489 VSS.n199 VSS.n129 4.5005
R15490 VSS.n188 VSS.n129 4.5005
R15491 VSS.n200 VSS.n129 4.5005
R15492 VSS.n187 VSS.n129 4.5005
R15493 VSS.n201 VSS.n129 4.5005
R15494 VSS.n186 VSS.n129 4.5005
R15495 VSS.n202 VSS.n129 4.5005
R15496 VSS.n185 VSS.n129 4.5005
R15497 VSS.n203 VSS.n129 4.5005
R15498 VSS.n184 VSS.n129 4.5005
R15499 VSS.n204 VSS.n129 4.5005
R15500 VSS.n183 VSS.n129 4.5005
R15501 VSS.n205 VSS.n129 4.5005
R15502 VSS.n182 VSS.n129 4.5005
R15503 VSS.n206 VSS.n129 4.5005
R15504 VSS.n181 VSS.n129 4.5005
R15505 VSS.n207 VSS.n129 4.5005
R15506 VSS.n180 VSS.n129 4.5005
R15507 VSS.n208 VSS.n129 4.5005
R15508 VSS.n179 VSS.n129 4.5005
R15509 VSS.n209 VSS.n129 4.5005
R15510 VSS.n178 VSS.n129 4.5005
R15511 VSS.n210 VSS.n129 4.5005
R15512 VSS.n177 VSS.n129 4.5005
R15513 VSS.n211 VSS.n129 4.5005
R15514 VSS.n176 VSS.n129 4.5005
R15515 VSS.n212 VSS.n129 4.5005
R15516 VSS.n175 VSS.n129 4.5005
R15517 VSS.n213 VSS.n129 4.5005
R15518 VSS.n174 VSS.n129 4.5005
R15519 VSS.n214 VSS.n129 4.5005
R15520 VSS.n173 VSS.n129 4.5005
R15521 VSS.n215 VSS.n129 4.5005
R15522 VSS.n172 VSS.n129 4.5005
R15523 VSS.n216 VSS.n129 4.5005
R15524 VSS.n171 VSS.n129 4.5005
R15525 VSS.n217 VSS.n129 4.5005
R15526 VSS.n170 VSS.n129 4.5005
R15527 VSS.n218 VSS.n129 4.5005
R15528 VSS.n169 VSS.n129 4.5005
R15529 VSS.n219 VSS.n129 4.5005
R15530 VSS.n168 VSS.n129 4.5005
R15531 VSS.n220 VSS.n129 4.5005
R15532 VSS.n167 VSS.n129 4.5005
R15533 VSS.n221 VSS.n129 4.5005
R15534 VSS.n166 VSS.n129 4.5005
R15535 VSS.n222 VSS.n129 4.5005
R15536 VSS.n165 VSS.n129 4.5005
R15537 VSS.n223 VSS.n129 4.5005
R15538 VSS.n164 VSS.n129 4.5005
R15539 VSS.n224 VSS.n129 4.5005
R15540 VSS.n163 VSS.n129 4.5005
R15541 VSS.n225 VSS.n129 4.5005
R15542 VSS.n162 VSS.n129 4.5005
R15543 VSS.n226 VSS.n129 4.5005
R15544 VSS.n161 VSS.n129 4.5005
R15545 VSS.n227 VSS.n129 4.5005
R15546 VSS.n160 VSS.n129 4.5005
R15547 VSS.n228 VSS.n129 4.5005
R15548 VSS.n159 VSS.n129 4.5005
R15549 VSS.n229 VSS.n129 4.5005
R15550 VSS.n158 VSS.n129 4.5005
R15551 VSS.n230 VSS.n129 4.5005
R15552 VSS.n157 VSS.n129 4.5005
R15553 VSS.n231 VSS.n129 4.5005
R15554 VSS.n156 VSS.n129 4.5005
R15555 VSS.n232 VSS.n129 4.5005
R15556 VSS.n155 VSS.n129 4.5005
R15557 VSS.n233 VSS.n129 4.5005
R15558 VSS.n154 VSS.n129 4.5005
R15559 VSS.n234 VSS.n129 4.5005
R15560 VSS.n153 VSS.n129 4.5005
R15561 VSS.n235 VSS.n129 4.5005
R15562 VSS.n4506 VSS.n129 4.5005
R15563 VSS.n236 VSS.n129 4.5005
R15564 VSS.n152 VSS.n129 4.5005
R15565 VSS.n237 VSS.n129 4.5005
R15566 VSS.n151 VSS.n129 4.5005
R15567 VSS.n238 VSS.n129 4.5005
R15568 VSS.n150 VSS.n129 4.5005
R15569 VSS.n239 VSS.n129 4.5005
R15570 VSS.n149 VSS.n129 4.5005
R15571 VSS.n240 VSS.n129 4.5005
R15572 VSS.n148 VSS.n129 4.5005
R15573 VSS.n241 VSS.n129 4.5005
R15574 VSS.n147 VSS.n129 4.5005
R15575 VSS.n242 VSS.n129 4.5005
R15576 VSS.n146 VSS.n129 4.5005
R15577 VSS.n243 VSS.n129 4.5005
R15578 VSS.n145 VSS.n129 4.5005
R15579 VSS.n244 VSS.n129 4.5005
R15580 VSS.n144 VSS.n129 4.5005
R15581 VSS.n245 VSS.n129 4.5005
R15582 VSS.n143 VSS.n129 4.5005
R15583 VSS.n246 VSS.n129 4.5005
R15584 VSS.n142 VSS.n129 4.5005
R15585 VSS.n247 VSS.n129 4.5005
R15586 VSS.n141 VSS.n129 4.5005
R15587 VSS.n248 VSS.n129 4.5005
R15588 VSS.n140 VSS.n129 4.5005
R15589 VSS.n249 VSS.n129 4.5005
R15590 VSS.n139 VSS.n129 4.5005
R15591 VSS.n250 VSS.n129 4.5005
R15592 VSS.n138 VSS.n129 4.5005
R15593 VSS.n251 VSS.n129 4.5005
R15594 VSS.n137 VSS.n129 4.5005
R15595 VSS.n252 VSS.n129 4.5005
R15596 VSS.n136 VSS.n129 4.5005
R15597 VSS.n253 VSS.n129 4.5005
R15598 VSS.n135 VSS.n129 4.5005
R15599 VSS.n254 VSS.n129 4.5005
R15600 VSS.n134 VSS.n129 4.5005
R15601 VSS.n255 VSS.n129 4.5005
R15602 VSS.n133 VSS.n129 4.5005
R15603 VSS.n256 VSS.n129 4.5005
R15604 VSS.n132 VSS.n129 4.5005
R15605 VSS.n4502 VSS.n129 4.5005
R15606 VSS.n4504 VSS.n129 4.5005
R15607 VSS.n193 VSS.n7 4.5005
R15608 VSS.n195 VSS.n7 4.5005
R15609 VSS.n192 VSS.n7 4.5005
R15610 VSS.n196 VSS.n7 4.5005
R15611 VSS.n191 VSS.n7 4.5005
R15612 VSS.n197 VSS.n7 4.5005
R15613 VSS.n190 VSS.n7 4.5005
R15614 VSS.n198 VSS.n7 4.5005
R15615 VSS.n189 VSS.n7 4.5005
R15616 VSS.n199 VSS.n7 4.5005
R15617 VSS.n188 VSS.n7 4.5005
R15618 VSS.n200 VSS.n7 4.5005
R15619 VSS.n187 VSS.n7 4.5005
R15620 VSS.n201 VSS.n7 4.5005
R15621 VSS.n186 VSS.n7 4.5005
R15622 VSS.n202 VSS.n7 4.5005
R15623 VSS.n185 VSS.n7 4.5005
R15624 VSS.n203 VSS.n7 4.5005
R15625 VSS.n184 VSS.n7 4.5005
R15626 VSS.n204 VSS.n7 4.5005
R15627 VSS.n183 VSS.n7 4.5005
R15628 VSS.n205 VSS.n7 4.5005
R15629 VSS.n182 VSS.n7 4.5005
R15630 VSS.n206 VSS.n7 4.5005
R15631 VSS.n181 VSS.n7 4.5005
R15632 VSS.n207 VSS.n7 4.5005
R15633 VSS.n180 VSS.n7 4.5005
R15634 VSS.n208 VSS.n7 4.5005
R15635 VSS.n179 VSS.n7 4.5005
R15636 VSS.n209 VSS.n7 4.5005
R15637 VSS.n178 VSS.n7 4.5005
R15638 VSS.n210 VSS.n7 4.5005
R15639 VSS.n177 VSS.n7 4.5005
R15640 VSS.n211 VSS.n7 4.5005
R15641 VSS.n176 VSS.n7 4.5005
R15642 VSS.n212 VSS.n7 4.5005
R15643 VSS.n175 VSS.n7 4.5005
R15644 VSS.n213 VSS.n7 4.5005
R15645 VSS.n174 VSS.n7 4.5005
R15646 VSS.n214 VSS.n7 4.5005
R15647 VSS.n173 VSS.n7 4.5005
R15648 VSS.n215 VSS.n7 4.5005
R15649 VSS.n172 VSS.n7 4.5005
R15650 VSS.n216 VSS.n7 4.5005
R15651 VSS.n171 VSS.n7 4.5005
R15652 VSS.n217 VSS.n7 4.5005
R15653 VSS.n170 VSS.n7 4.5005
R15654 VSS.n218 VSS.n7 4.5005
R15655 VSS.n169 VSS.n7 4.5005
R15656 VSS.n219 VSS.n7 4.5005
R15657 VSS.n168 VSS.n7 4.5005
R15658 VSS.n220 VSS.n7 4.5005
R15659 VSS.n167 VSS.n7 4.5005
R15660 VSS.n221 VSS.n7 4.5005
R15661 VSS.n166 VSS.n7 4.5005
R15662 VSS.n222 VSS.n7 4.5005
R15663 VSS.n165 VSS.n7 4.5005
R15664 VSS.n223 VSS.n7 4.5005
R15665 VSS.n164 VSS.n7 4.5005
R15666 VSS.n224 VSS.n7 4.5005
R15667 VSS.n163 VSS.n7 4.5005
R15668 VSS.n225 VSS.n7 4.5005
R15669 VSS.n162 VSS.n7 4.5005
R15670 VSS.n226 VSS.n7 4.5005
R15671 VSS.n161 VSS.n7 4.5005
R15672 VSS.n227 VSS.n7 4.5005
R15673 VSS.n160 VSS.n7 4.5005
R15674 VSS.n228 VSS.n7 4.5005
R15675 VSS.n159 VSS.n7 4.5005
R15676 VSS.n229 VSS.n7 4.5005
R15677 VSS.n158 VSS.n7 4.5005
R15678 VSS.n230 VSS.n7 4.5005
R15679 VSS.n157 VSS.n7 4.5005
R15680 VSS.n231 VSS.n7 4.5005
R15681 VSS.n156 VSS.n7 4.5005
R15682 VSS.n232 VSS.n7 4.5005
R15683 VSS.n155 VSS.n7 4.5005
R15684 VSS.n233 VSS.n7 4.5005
R15685 VSS.n154 VSS.n7 4.5005
R15686 VSS.n234 VSS.n7 4.5005
R15687 VSS.n153 VSS.n7 4.5005
R15688 VSS.n235 VSS.n7 4.5005
R15689 VSS.n4506 VSS.n7 4.5005
R15690 VSS.n236 VSS.n7 4.5005
R15691 VSS.n152 VSS.n7 4.5005
R15692 VSS.n237 VSS.n7 4.5005
R15693 VSS.n151 VSS.n7 4.5005
R15694 VSS.n238 VSS.n7 4.5005
R15695 VSS.n150 VSS.n7 4.5005
R15696 VSS.n239 VSS.n7 4.5005
R15697 VSS.n149 VSS.n7 4.5005
R15698 VSS.n240 VSS.n7 4.5005
R15699 VSS.n148 VSS.n7 4.5005
R15700 VSS.n241 VSS.n7 4.5005
R15701 VSS.n147 VSS.n7 4.5005
R15702 VSS.n242 VSS.n7 4.5005
R15703 VSS.n146 VSS.n7 4.5005
R15704 VSS.n243 VSS.n7 4.5005
R15705 VSS.n145 VSS.n7 4.5005
R15706 VSS.n244 VSS.n7 4.5005
R15707 VSS.n144 VSS.n7 4.5005
R15708 VSS.n245 VSS.n7 4.5005
R15709 VSS.n143 VSS.n7 4.5005
R15710 VSS.n246 VSS.n7 4.5005
R15711 VSS.n142 VSS.n7 4.5005
R15712 VSS.n247 VSS.n7 4.5005
R15713 VSS.n141 VSS.n7 4.5005
R15714 VSS.n248 VSS.n7 4.5005
R15715 VSS.n140 VSS.n7 4.5005
R15716 VSS.n249 VSS.n7 4.5005
R15717 VSS.n139 VSS.n7 4.5005
R15718 VSS.n250 VSS.n7 4.5005
R15719 VSS.n138 VSS.n7 4.5005
R15720 VSS.n251 VSS.n7 4.5005
R15721 VSS.n137 VSS.n7 4.5005
R15722 VSS.n252 VSS.n7 4.5005
R15723 VSS.n136 VSS.n7 4.5005
R15724 VSS.n253 VSS.n7 4.5005
R15725 VSS.n135 VSS.n7 4.5005
R15726 VSS.n254 VSS.n7 4.5005
R15727 VSS.n134 VSS.n7 4.5005
R15728 VSS.n255 VSS.n7 4.5005
R15729 VSS.n133 VSS.n7 4.5005
R15730 VSS.n256 VSS.n7 4.5005
R15731 VSS.n132 VSS.n7 4.5005
R15732 VSS.n4502 VSS.n7 4.5005
R15733 VSS.n4504 VSS.n7 4.5005
R15734 VSS.n193 VSS.n130 4.5005
R15735 VSS.n195 VSS.n130 4.5005
R15736 VSS.n192 VSS.n130 4.5005
R15737 VSS.n196 VSS.n130 4.5005
R15738 VSS.n191 VSS.n130 4.5005
R15739 VSS.n197 VSS.n130 4.5005
R15740 VSS.n190 VSS.n130 4.5005
R15741 VSS.n198 VSS.n130 4.5005
R15742 VSS.n189 VSS.n130 4.5005
R15743 VSS.n199 VSS.n130 4.5005
R15744 VSS.n188 VSS.n130 4.5005
R15745 VSS.n200 VSS.n130 4.5005
R15746 VSS.n187 VSS.n130 4.5005
R15747 VSS.n201 VSS.n130 4.5005
R15748 VSS.n186 VSS.n130 4.5005
R15749 VSS.n202 VSS.n130 4.5005
R15750 VSS.n185 VSS.n130 4.5005
R15751 VSS.n203 VSS.n130 4.5005
R15752 VSS.n184 VSS.n130 4.5005
R15753 VSS.n204 VSS.n130 4.5005
R15754 VSS.n183 VSS.n130 4.5005
R15755 VSS.n205 VSS.n130 4.5005
R15756 VSS.n182 VSS.n130 4.5005
R15757 VSS.n206 VSS.n130 4.5005
R15758 VSS.n181 VSS.n130 4.5005
R15759 VSS.n207 VSS.n130 4.5005
R15760 VSS.n180 VSS.n130 4.5005
R15761 VSS.n208 VSS.n130 4.5005
R15762 VSS.n179 VSS.n130 4.5005
R15763 VSS.n209 VSS.n130 4.5005
R15764 VSS.n178 VSS.n130 4.5005
R15765 VSS.n210 VSS.n130 4.5005
R15766 VSS.n177 VSS.n130 4.5005
R15767 VSS.n211 VSS.n130 4.5005
R15768 VSS.n176 VSS.n130 4.5005
R15769 VSS.n212 VSS.n130 4.5005
R15770 VSS.n175 VSS.n130 4.5005
R15771 VSS.n213 VSS.n130 4.5005
R15772 VSS.n174 VSS.n130 4.5005
R15773 VSS.n214 VSS.n130 4.5005
R15774 VSS.n173 VSS.n130 4.5005
R15775 VSS.n215 VSS.n130 4.5005
R15776 VSS.n172 VSS.n130 4.5005
R15777 VSS.n216 VSS.n130 4.5005
R15778 VSS.n171 VSS.n130 4.5005
R15779 VSS.n217 VSS.n130 4.5005
R15780 VSS.n170 VSS.n130 4.5005
R15781 VSS.n218 VSS.n130 4.5005
R15782 VSS.n169 VSS.n130 4.5005
R15783 VSS.n219 VSS.n130 4.5005
R15784 VSS.n168 VSS.n130 4.5005
R15785 VSS.n220 VSS.n130 4.5005
R15786 VSS.n167 VSS.n130 4.5005
R15787 VSS.n221 VSS.n130 4.5005
R15788 VSS.n166 VSS.n130 4.5005
R15789 VSS.n222 VSS.n130 4.5005
R15790 VSS.n165 VSS.n130 4.5005
R15791 VSS.n223 VSS.n130 4.5005
R15792 VSS.n164 VSS.n130 4.5005
R15793 VSS.n224 VSS.n130 4.5005
R15794 VSS.n163 VSS.n130 4.5005
R15795 VSS.n225 VSS.n130 4.5005
R15796 VSS.n162 VSS.n130 4.5005
R15797 VSS.n226 VSS.n130 4.5005
R15798 VSS.n161 VSS.n130 4.5005
R15799 VSS.n227 VSS.n130 4.5005
R15800 VSS.n160 VSS.n130 4.5005
R15801 VSS.n228 VSS.n130 4.5005
R15802 VSS.n159 VSS.n130 4.5005
R15803 VSS.n229 VSS.n130 4.5005
R15804 VSS.n158 VSS.n130 4.5005
R15805 VSS.n230 VSS.n130 4.5005
R15806 VSS.n157 VSS.n130 4.5005
R15807 VSS.n231 VSS.n130 4.5005
R15808 VSS.n156 VSS.n130 4.5005
R15809 VSS.n232 VSS.n130 4.5005
R15810 VSS.n155 VSS.n130 4.5005
R15811 VSS.n233 VSS.n130 4.5005
R15812 VSS.n154 VSS.n130 4.5005
R15813 VSS.n234 VSS.n130 4.5005
R15814 VSS.n153 VSS.n130 4.5005
R15815 VSS.n235 VSS.n130 4.5005
R15816 VSS.n4506 VSS.n130 4.5005
R15817 VSS.n236 VSS.n130 4.5005
R15818 VSS.n152 VSS.n130 4.5005
R15819 VSS.n237 VSS.n130 4.5005
R15820 VSS.n151 VSS.n130 4.5005
R15821 VSS.n238 VSS.n130 4.5005
R15822 VSS.n150 VSS.n130 4.5005
R15823 VSS.n239 VSS.n130 4.5005
R15824 VSS.n149 VSS.n130 4.5005
R15825 VSS.n240 VSS.n130 4.5005
R15826 VSS.n148 VSS.n130 4.5005
R15827 VSS.n241 VSS.n130 4.5005
R15828 VSS.n147 VSS.n130 4.5005
R15829 VSS.n242 VSS.n130 4.5005
R15830 VSS.n146 VSS.n130 4.5005
R15831 VSS.n243 VSS.n130 4.5005
R15832 VSS.n145 VSS.n130 4.5005
R15833 VSS.n244 VSS.n130 4.5005
R15834 VSS.n144 VSS.n130 4.5005
R15835 VSS.n245 VSS.n130 4.5005
R15836 VSS.n143 VSS.n130 4.5005
R15837 VSS.n246 VSS.n130 4.5005
R15838 VSS.n142 VSS.n130 4.5005
R15839 VSS.n247 VSS.n130 4.5005
R15840 VSS.n141 VSS.n130 4.5005
R15841 VSS.n248 VSS.n130 4.5005
R15842 VSS.n140 VSS.n130 4.5005
R15843 VSS.n249 VSS.n130 4.5005
R15844 VSS.n139 VSS.n130 4.5005
R15845 VSS.n250 VSS.n130 4.5005
R15846 VSS.n138 VSS.n130 4.5005
R15847 VSS.n251 VSS.n130 4.5005
R15848 VSS.n137 VSS.n130 4.5005
R15849 VSS.n252 VSS.n130 4.5005
R15850 VSS.n136 VSS.n130 4.5005
R15851 VSS.n253 VSS.n130 4.5005
R15852 VSS.n135 VSS.n130 4.5005
R15853 VSS.n254 VSS.n130 4.5005
R15854 VSS.n134 VSS.n130 4.5005
R15855 VSS.n255 VSS.n130 4.5005
R15856 VSS.n133 VSS.n130 4.5005
R15857 VSS.n256 VSS.n130 4.5005
R15858 VSS.n132 VSS.n130 4.5005
R15859 VSS.n4502 VSS.n130 4.5005
R15860 VSS.n4504 VSS.n130 4.5005
R15861 VSS.n193 VSS.n6 4.5005
R15862 VSS.n195 VSS.n6 4.5005
R15863 VSS.n192 VSS.n6 4.5005
R15864 VSS.n196 VSS.n6 4.5005
R15865 VSS.n191 VSS.n6 4.5005
R15866 VSS.n197 VSS.n6 4.5005
R15867 VSS.n190 VSS.n6 4.5005
R15868 VSS.n198 VSS.n6 4.5005
R15869 VSS.n189 VSS.n6 4.5005
R15870 VSS.n199 VSS.n6 4.5005
R15871 VSS.n188 VSS.n6 4.5005
R15872 VSS.n200 VSS.n6 4.5005
R15873 VSS.n187 VSS.n6 4.5005
R15874 VSS.n201 VSS.n6 4.5005
R15875 VSS.n186 VSS.n6 4.5005
R15876 VSS.n202 VSS.n6 4.5005
R15877 VSS.n185 VSS.n6 4.5005
R15878 VSS.n203 VSS.n6 4.5005
R15879 VSS.n184 VSS.n6 4.5005
R15880 VSS.n204 VSS.n6 4.5005
R15881 VSS.n183 VSS.n6 4.5005
R15882 VSS.n205 VSS.n6 4.5005
R15883 VSS.n182 VSS.n6 4.5005
R15884 VSS.n206 VSS.n6 4.5005
R15885 VSS.n181 VSS.n6 4.5005
R15886 VSS.n207 VSS.n6 4.5005
R15887 VSS.n180 VSS.n6 4.5005
R15888 VSS.n208 VSS.n6 4.5005
R15889 VSS.n179 VSS.n6 4.5005
R15890 VSS.n209 VSS.n6 4.5005
R15891 VSS.n178 VSS.n6 4.5005
R15892 VSS.n210 VSS.n6 4.5005
R15893 VSS.n177 VSS.n6 4.5005
R15894 VSS.n211 VSS.n6 4.5005
R15895 VSS.n176 VSS.n6 4.5005
R15896 VSS.n212 VSS.n6 4.5005
R15897 VSS.n175 VSS.n6 4.5005
R15898 VSS.n213 VSS.n6 4.5005
R15899 VSS.n174 VSS.n6 4.5005
R15900 VSS.n214 VSS.n6 4.5005
R15901 VSS.n173 VSS.n6 4.5005
R15902 VSS.n215 VSS.n6 4.5005
R15903 VSS.n172 VSS.n6 4.5005
R15904 VSS.n216 VSS.n6 4.5005
R15905 VSS.n171 VSS.n6 4.5005
R15906 VSS.n217 VSS.n6 4.5005
R15907 VSS.n170 VSS.n6 4.5005
R15908 VSS.n218 VSS.n6 4.5005
R15909 VSS.n169 VSS.n6 4.5005
R15910 VSS.n219 VSS.n6 4.5005
R15911 VSS.n168 VSS.n6 4.5005
R15912 VSS.n220 VSS.n6 4.5005
R15913 VSS.n167 VSS.n6 4.5005
R15914 VSS.n221 VSS.n6 4.5005
R15915 VSS.n166 VSS.n6 4.5005
R15916 VSS.n222 VSS.n6 4.5005
R15917 VSS.n165 VSS.n6 4.5005
R15918 VSS.n223 VSS.n6 4.5005
R15919 VSS.n164 VSS.n6 4.5005
R15920 VSS.n224 VSS.n6 4.5005
R15921 VSS.n163 VSS.n6 4.5005
R15922 VSS.n225 VSS.n6 4.5005
R15923 VSS.n162 VSS.n6 4.5005
R15924 VSS.n226 VSS.n6 4.5005
R15925 VSS.n161 VSS.n6 4.5005
R15926 VSS.n227 VSS.n6 4.5005
R15927 VSS.n160 VSS.n6 4.5005
R15928 VSS.n228 VSS.n6 4.5005
R15929 VSS.n159 VSS.n6 4.5005
R15930 VSS.n229 VSS.n6 4.5005
R15931 VSS.n158 VSS.n6 4.5005
R15932 VSS.n230 VSS.n6 4.5005
R15933 VSS.n157 VSS.n6 4.5005
R15934 VSS.n231 VSS.n6 4.5005
R15935 VSS.n156 VSS.n6 4.5005
R15936 VSS.n232 VSS.n6 4.5005
R15937 VSS.n155 VSS.n6 4.5005
R15938 VSS.n233 VSS.n6 4.5005
R15939 VSS.n154 VSS.n6 4.5005
R15940 VSS.n234 VSS.n6 4.5005
R15941 VSS.n153 VSS.n6 4.5005
R15942 VSS.n235 VSS.n6 4.5005
R15943 VSS.n4506 VSS.n6 4.5005
R15944 VSS.n236 VSS.n6 4.5005
R15945 VSS.n152 VSS.n6 4.5005
R15946 VSS.n237 VSS.n6 4.5005
R15947 VSS.n151 VSS.n6 4.5005
R15948 VSS.n238 VSS.n6 4.5005
R15949 VSS.n150 VSS.n6 4.5005
R15950 VSS.n239 VSS.n6 4.5005
R15951 VSS.n149 VSS.n6 4.5005
R15952 VSS.n240 VSS.n6 4.5005
R15953 VSS.n148 VSS.n6 4.5005
R15954 VSS.n241 VSS.n6 4.5005
R15955 VSS.n147 VSS.n6 4.5005
R15956 VSS.n242 VSS.n6 4.5005
R15957 VSS.n146 VSS.n6 4.5005
R15958 VSS.n243 VSS.n6 4.5005
R15959 VSS.n145 VSS.n6 4.5005
R15960 VSS.n244 VSS.n6 4.5005
R15961 VSS.n144 VSS.n6 4.5005
R15962 VSS.n245 VSS.n6 4.5005
R15963 VSS.n143 VSS.n6 4.5005
R15964 VSS.n246 VSS.n6 4.5005
R15965 VSS.n142 VSS.n6 4.5005
R15966 VSS.n247 VSS.n6 4.5005
R15967 VSS.n141 VSS.n6 4.5005
R15968 VSS.n248 VSS.n6 4.5005
R15969 VSS.n140 VSS.n6 4.5005
R15970 VSS.n249 VSS.n6 4.5005
R15971 VSS.n139 VSS.n6 4.5005
R15972 VSS.n250 VSS.n6 4.5005
R15973 VSS.n138 VSS.n6 4.5005
R15974 VSS.n251 VSS.n6 4.5005
R15975 VSS.n137 VSS.n6 4.5005
R15976 VSS.n252 VSS.n6 4.5005
R15977 VSS.n136 VSS.n6 4.5005
R15978 VSS.n253 VSS.n6 4.5005
R15979 VSS.n135 VSS.n6 4.5005
R15980 VSS.n254 VSS.n6 4.5005
R15981 VSS.n134 VSS.n6 4.5005
R15982 VSS.n255 VSS.n6 4.5005
R15983 VSS.n133 VSS.n6 4.5005
R15984 VSS.n256 VSS.n6 4.5005
R15985 VSS.n132 VSS.n6 4.5005
R15986 VSS.n4502 VSS.n6 4.5005
R15987 VSS.n4504 VSS.n6 4.5005
R15988 VSS.n193 VSS.n131 4.5005
R15989 VSS.n195 VSS.n131 4.5005
R15990 VSS.n192 VSS.n131 4.5005
R15991 VSS.n196 VSS.n131 4.5005
R15992 VSS.n191 VSS.n131 4.5005
R15993 VSS.n197 VSS.n131 4.5005
R15994 VSS.n190 VSS.n131 4.5005
R15995 VSS.n198 VSS.n131 4.5005
R15996 VSS.n189 VSS.n131 4.5005
R15997 VSS.n199 VSS.n131 4.5005
R15998 VSS.n188 VSS.n131 4.5005
R15999 VSS.n200 VSS.n131 4.5005
R16000 VSS.n187 VSS.n131 4.5005
R16001 VSS.n201 VSS.n131 4.5005
R16002 VSS.n186 VSS.n131 4.5005
R16003 VSS.n202 VSS.n131 4.5005
R16004 VSS.n185 VSS.n131 4.5005
R16005 VSS.n203 VSS.n131 4.5005
R16006 VSS.n184 VSS.n131 4.5005
R16007 VSS.n204 VSS.n131 4.5005
R16008 VSS.n183 VSS.n131 4.5005
R16009 VSS.n205 VSS.n131 4.5005
R16010 VSS.n182 VSS.n131 4.5005
R16011 VSS.n206 VSS.n131 4.5005
R16012 VSS.n181 VSS.n131 4.5005
R16013 VSS.n207 VSS.n131 4.5005
R16014 VSS.n180 VSS.n131 4.5005
R16015 VSS.n208 VSS.n131 4.5005
R16016 VSS.n179 VSS.n131 4.5005
R16017 VSS.n209 VSS.n131 4.5005
R16018 VSS.n178 VSS.n131 4.5005
R16019 VSS.n210 VSS.n131 4.5005
R16020 VSS.n177 VSS.n131 4.5005
R16021 VSS.n211 VSS.n131 4.5005
R16022 VSS.n176 VSS.n131 4.5005
R16023 VSS.n212 VSS.n131 4.5005
R16024 VSS.n175 VSS.n131 4.5005
R16025 VSS.n213 VSS.n131 4.5005
R16026 VSS.n174 VSS.n131 4.5005
R16027 VSS.n214 VSS.n131 4.5005
R16028 VSS.n173 VSS.n131 4.5005
R16029 VSS.n215 VSS.n131 4.5005
R16030 VSS.n172 VSS.n131 4.5005
R16031 VSS.n216 VSS.n131 4.5005
R16032 VSS.n171 VSS.n131 4.5005
R16033 VSS.n217 VSS.n131 4.5005
R16034 VSS.n170 VSS.n131 4.5005
R16035 VSS.n218 VSS.n131 4.5005
R16036 VSS.n169 VSS.n131 4.5005
R16037 VSS.n219 VSS.n131 4.5005
R16038 VSS.n168 VSS.n131 4.5005
R16039 VSS.n220 VSS.n131 4.5005
R16040 VSS.n167 VSS.n131 4.5005
R16041 VSS.n221 VSS.n131 4.5005
R16042 VSS.n166 VSS.n131 4.5005
R16043 VSS.n222 VSS.n131 4.5005
R16044 VSS.n165 VSS.n131 4.5005
R16045 VSS.n223 VSS.n131 4.5005
R16046 VSS.n164 VSS.n131 4.5005
R16047 VSS.n224 VSS.n131 4.5005
R16048 VSS.n163 VSS.n131 4.5005
R16049 VSS.n225 VSS.n131 4.5005
R16050 VSS.n162 VSS.n131 4.5005
R16051 VSS.n226 VSS.n131 4.5005
R16052 VSS.n161 VSS.n131 4.5005
R16053 VSS.n227 VSS.n131 4.5005
R16054 VSS.n160 VSS.n131 4.5005
R16055 VSS.n228 VSS.n131 4.5005
R16056 VSS.n159 VSS.n131 4.5005
R16057 VSS.n229 VSS.n131 4.5005
R16058 VSS.n158 VSS.n131 4.5005
R16059 VSS.n230 VSS.n131 4.5005
R16060 VSS.n157 VSS.n131 4.5005
R16061 VSS.n231 VSS.n131 4.5005
R16062 VSS.n156 VSS.n131 4.5005
R16063 VSS.n232 VSS.n131 4.5005
R16064 VSS.n155 VSS.n131 4.5005
R16065 VSS.n233 VSS.n131 4.5005
R16066 VSS.n154 VSS.n131 4.5005
R16067 VSS.n234 VSS.n131 4.5005
R16068 VSS.n153 VSS.n131 4.5005
R16069 VSS.n235 VSS.n131 4.5005
R16070 VSS.n4506 VSS.n131 4.5005
R16071 VSS.n236 VSS.n131 4.5005
R16072 VSS.n152 VSS.n131 4.5005
R16073 VSS.n237 VSS.n131 4.5005
R16074 VSS.n151 VSS.n131 4.5005
R16075 VSS.n238 VSS.n131 4.5005
R16076 VSS.n150 VSS.n131 4.5005
R16077 VSS.n239 VSS.n131 4.5005
R16078 VSS.n149 VSS.n131 4.5005
R16079 VSS.n240 VSS.n131 4.5005
R16080 VSS.n148 VSS.n131 4.5005
R16081 VSS.n241 VSS.n131 4.5005
R16082 VSS.n147 VSS.n131 4.5005
R16083 VSS.n242 VSS.n131 4.5005
R16084 VSS.n146 VSS.n131 4.5005
R16085 VSS.n243 VSS.n131 4.5005
R16086 VSS.n145 VSS.n131 4.5005
R16087 VSS.n244 VSS.n131 4.5005
R16088 VSS.n144 VSS.n131 4.5005
R16089 VSS.n245 VSS.n131 4.5005
R16090 VSS.n143 VSS.n131 4.5005
R16091 VSS.n246 VSS.n131 4.5005
R16092 VSS.n142 VSS.n131 4.5005
R16093 VSS.n247 VSS.n131 4.5005
R16094 VSS.n141 VSS.n131 4.5005
R16095 VSS.n248 VSS.n131 4.5005
R16096 VSS.n140 VSS.n131 4.5005
R16097 VSS.n249 VSS.n131 4.5005
R16098 VSS.n139 VSS.n131 4.5005
R16099 VSS.n250 VSS.n131 4.5005
R16100 VSS.n138 VSS.n131 4.5005
R16101 VSS.n251 VSS.n131 4.5005
R16102 VSS.n137 VSS.n131 4.5005
R16103 VSS.n252 VSS.n131 4.5005
R16104 VSS.n136 VSS.n131 4.5005
R16105 VSS.n253 VSS.n131 4.5005
R16106 VSS.n135 VSS.n131 4.5005
R16107 VSS.n254 VSS.n131 4.5005
R16108 VSS.n134 VSS.n131 4.5005
R16109 VSS.n255 VSS.n131 4.5005
R16110 VSS.n133 VSS.n131 4.5005
R16111 VSS.n256 VSS.n131 4.5005
R16112 VSS.n132 VSS.n131 4.5005
R16113 VSS.n4502 VSS.n131 4.5005
R16114 VSS.n4504 VSS.n131 4.5005
R16115 VSS.n193 VSS.n5 4.5005
R16116 VSS.n195 VSS.n5 4.5005
R16117 VSS.n192 VSS.n5 4.5005
R16118 VSS.n196 VSS.n5 4.5005
R16119 VSS.n191 VSS.n5 4.5005
R16120 VSS.n197 VSS.n5 4.5005
R16121 VSS.n190 VSS.n5 4.5005
R16122 VSS.n198 VSS.n5 4.5005
R16123 VSS.n189 VSS.n5 4.5005
R16124 VSS.n199 VSS.n5 4.5005
R16125 VSS.n188 VSS.n5 4.5005
R16126 VSS.n200 VSS.n5 4.5005
R16127 VSS.n187 VSS.n5 4.5005
R16128 VSS.n201 VSS.n5 4.5005
R16129 VSS.n186 VSS.n5 4.5005
R16130 VSS.n202 VSS.n5 4.5005
R16131 VSS.n185 VSS.n5 4.5005
R16132 VSS.n203 VSS.n5 4.5005
R16133 VSS.n184 VSS.n5 4.5005
R16134 VSS.n204 VSS.n5 4.5005
R16135 VSS.n183 VSS.n5 4.5005
R16136 VSS.n205 VSS.n5 4.5005
R16137 VSS.n182 VSS.n5 4.5005
R16138 VSS.n206 VSS.n5 4.5005
R16139 VSS.n181 VSS.n5 4.5005
R16140 VSS.n207 VSS.n5 4.5005
R16141 VSS.n180 VSS.n5 4.5005
R16142 VSS.n208 VSS.n5 4.5005
R16143 VSS.n179 VSS.n5 4.5005
R16144 VSS.n209 VSS.n5 4.5005
R16145 VSS.n178 VSS.n5 4.5005
R16146 VSS.n210 VSS.n5 4.5005
R16147 VSS.n177 VSS.n5 4.5005
R16148 VSS.n211 VSS.n5 4.5005
R16149 VSS.n176 VSS.n5 4.5005
R16150 VSS.n212 VSS.n5 4.5005
R16151 VSS.n175 VSS.n5 4.5005
R16152 VSS.n213 VSS.n5 4.5005
R16153 VSS.n174 VSS.n5 4.5005
R16154 VSS.n214 VSS.n5 4.5005
R16155 VSS.n173 VSS.n5 4.5005
R16156 VSS.n215 VSS.n5 4.5005
R16157 VSS.n172 VSS.n5 4.5005
R16158 VSS.n216 VSS.n5 4.5005
R16159 VSS.n171 VSS.n5 4.5005
R16160 VSS.n217 VSS.n5 4.5005
R16161 VSS.n170 VSS.n5 4.5005
R16162 VSS.n218 VSS.n5 4.5005
R16163 VSS.n169 VSS.n5 4.5005
R16164 VSS.n219 VSS.n5 4.5005
R16165 VSS.n168 VSS.n5 4.5005
R16166 VSS.n220 VSS.n5 4.5005
R16167 VSS.n167 VSS.n5 4.5005
R16168 VSS.n221 VSS.n5 4.5005
R16169 VSS.n166 VSS.n5 4.5005
R16170 VSS.n222 VSS.n5 4.5005
R16171 VSS.n165 VSS.n5 4.5005
R16172 VSS.n223 VSS.n5 4.5005
R16173 VSS.n164 VSS.n5 4.5005
R16174 VSS.n224 VSS.n5 4.5005
R16175 VSS.n163 VSS.n5 4.5005
R16176 VSS.n225 VSS.n5 4.5005
R16177 VSS.n162 VSS.n5 4.5005
R16178 VSS.n226 VSS.n5 4.5005
R16179 VSS.n161 VSS.n5 4.5005
R16180 VSS.n227 VSS.n5 4.5005
R16181 VSS.n160 VSS.n5 4.5005
R16182 VSS.n228 VSS.n5 4.5005
R16183 VSS.n159 VSS.n5 4.5005
R16184 VSS.n229 VSS.n5 4.5005
R16185 VSS.n158 VSS.n5 4.5005
R16186 VSS.n230 VSS.n5 4.5005
R16187 VSS.n157 VSS.n5 4.5005
R16188 VSS.n231 VSS.n5 4.5005
R16189 VSS.n156 VSS.n5 4.5005
R16190 VSS.n232 VSS.n5 4.5005
R16191 VSS.n155 VSS.n5 4.5005
R16192 VSS.n233 VSS.n5 4.5005
R16193 VSS.n154 VSS.n5 4.5005
R16194 VSS.n234 VSS.n5 4.5005
R16195 VSS.n153 VSS.n5 4.5005
R16196 VSS.n235 VSS.n5 4.5005
R16197 VSS.n4506 VSS.n5 4.5005
R16198 VSS.n236 VSS.n5 4.5005
R16199 VSS.n152 VSS.n5 4.5005
R16200 VSS.n237 VSS.n5 4.5005
R16201 VSS.n151 VSS.n5 4.5005
R16202 VSS.n238 VSS.n5 4.5005
R16203 VSS.n150 VSS.n5 4.5005
R16204 VSS.n239 VSS.n5 4.5005
R16205 VSS.n149 VSS.n5 4.5005
R16206 VSS.n240 VSS.n5 4.5005
R16207 VSS.n148 VSS.n5 4.5005
R16208 VSS.n241 VSS.n5 4.5005
R16209 VSS.n147 VSS.n5 4.5005
R16210 VSS.n242 VSS.n5 4.5005
R16211 VSS.n146 VSS.n5 4.5005
R16212 VSS.n243 VSS.n5 4.5005
R16213 VSS.n145 VSS.n5 4.5005
R16214 VSS.n244 VSS.n5 4.5005
R16215 VSS.n144 VSS.n5 4.5005
R16216 VSS.n245 VSS.n5 4.5005
R16217 VSS.n143 VSS.n5 4.5005
R16218 VSS.n246 VSS.n5 4.5005
R16219 VSS.n142 VSS.n5 4.5005
R16220 VSS.n247 VSS.n5 4.5005
R16221 VSS.n141 VSS.n5 4.5005
R16222 VSS.n248 VSS.n5 4.5005
R16223 VSS.n140 VSS.n5 4.5005
R16224 VSS.n249 VSS.n5 4.5005
R16225 VSS.n139 VSS.n5 4.5005
R16226 VSS.n250 VSS.n5 4.5005
R16227 VSS.n138 VSS.n5 4.5005
R16228 VSS.n251 VSS.n5 4.5005
R16229 VSS.n137 VSS.n5 4.5005
R16230 VSS.n252 VSS.n5 4.5005
R16231 VSS.n136 VSS.n5 4.5005
R16232 VSS.n253 VSS.n5 4.5005
R16233 VSS.n135 VSS.n5 4.5005
R16234 VSS.n254 VSS.n5 4.5005
R16235 VSS.n134 VSS.n5 4.5005
R16236 VSS.n255 VSS.n5 4.5005
R16237 VSS.n133 VSS.n5 4.5005
R16238 VSS.n256 VSS.n5 4.5005
R16239 VSS.n132 VSS.n5 4.5005
R16240 VSS.n4502 VSS.n5 4.5005
R16241 VSS.n4504 VSS.n5 4.5005
R16242 VSS.n4505 VSS.n193 4.5005
R16243 VSS.n4505 VSS.n195 4.5005
R16244 VSS.n4505 VSS.n192 4.5005
R16245 VSS.n4505 VSS.n196 4.5005
R16246 VSS.n4505 VSS.n191 4.5005
R16247 VSS.n4505 VSS.n197 4.5005
R16248 VSS.n4505 VSS.n190 4.5005
R16249 VSS.n4505 VSS.n198 4.5005
R16250 VSS.n4505 VSS.n189 4.5005
R16251 VSS.n4505 VSS.n199 4.5005
R16252 VSS.n4505 VSS.n188 4.5005
R16253 VSS.n4505 VSS.n200 4.5005
R16254 VSS.n4505 VSS.n187 4.5005
R16255 VSS.n4505 VSS.n201 4.5005
R16256 VSS.n4505 VSS.n186 4.5005
R16257 VSS.n4505 VSS.n202 4.5005
R16258 VSS.n4505 VSS.n185 4.5005
R16259 VSS.n4505 VSS.n203 4.5005
R16260 VSS.n4505 VSS.n184 4.5005
R16261 VSS.n4505 VSS.n204 4.5005
R16262 VSS.n4505 VSS.n183 4.5005
R16263 VSS.n4505 VSS.n205 4.5005
R16264 VSS.n4505 VSS.n182 4.5005
R16265 VSS.n4505 VSS.n206 4.5005
R16266 VSS.n4505 VSS.n181 4.5005
R16267 VSS.n4505 VSS.n207 4.5005
R16268 VSS.n4505 VSS.n180 4.5005
R16269 VSS.n4505 VSS.n208 4.5005
R16270 VSS.n4505 VSS.n179 4.5005
R16271 VSS.n4505 VSS.n209 4.5005
R16272 VSS.n4505 VSS.n178 4.5005
R16273 VSS.n4505 VSS.n210 4.5005
R16274 VSS.n4505 VSS.n177 4.5005
R16275 VSS.n4505 VSS.n211 4.5005
R16276 VSS.n4505 VSS.n176 4.5005
R16277 VSS.n4505 VSS.n212 4.5005
R16278 VSS.n4505 VSS.n175 4.5005
R16279 VSS.n4505 VSS.n213 4.5005
R16280 VSS.n4505 VSS.n174 4.5005
R16281 VSS.n4505 VSS.n214 4.5005
R16282 VSS.n4505 VSS.n173 4.5005
R16283 VSS.n4505 VSS.n215 4.5005
R16284 VSS.n4505 VSS.n172 4.5005
R16285 VSS.n4505 VSS.n216 4.5005
R16286 VSS.n4505 VSS.n171 4.5005
R16287 VSS.n4505 VSS.n217 4.5005
R16288 VSS.n4505 VSS.n170 4.5005
R16289 VSS.n4505 VSS.n218 4.5005
R16290 VSS.n4505 VSS.n169 4.5005
R16291 VSS.n4505 VSS.n219 4.5005
R16292 VSS.n4505 VSS.n168 4.5005
R16293 VSS.n4505 VSS.n220 4.5005
R16294 VSS.n4505 VSS.n167 4.5005
R16295 VSS.n4505 VSS.n221 4.5005
R16296 VSS.n4505 VSS.n166 4.5005
R16297 VSS.n4505 VSS.n222 4.5005
R16298 VSS.n4505 VSS.n165 4.5005
R16299 VSS.n4505 VSS.n223 4.5005
R16300 VSS.n4505 VSS.n164 4.5005
R16301 VSS.n4505 VSS.n224 4.5005
R16302 VSS.n4505 VSS.n163 4.5005
R16303 VSS.n4505 VSS.n225 4.5005
R16304 VSS.n4505 VSS.n162 4.5005
R16305 VSS.n4505 VSS.n226 4.5005
R16306 VSS.n4505 VSS.n161 4.5005
R16307 VSS.n4505 VSS.n227 4.5005
R16308 VSS.n4505 VSS.n160 4.5005
R16309 VSS.n4505 VSS.n228 4.5005
R16310 VSS.n4505 VSS.n159 4.5005
R16311 VSS.n4505 VSS.n229 4.5005
R16312 VSS.n4505 VSS.n158 4.5005
R16313 VSS.n4505 VSS.n230 4.5005
R16314 VSS.n4505 VSS.n157 4.5005
R16315 VSS.n4505 VSS.n231 4.5005
R16316 VSS.n4505 VSS.n156 4.5005
R16317 VSS.n4505 VSS.n232 4.5005
R16318 VSS.n4505 VSS.n155 4.5005
R16319 VSS.n4505 VSS.n233 4.5005
R16320 VSS.n4505 VSS.n154 4.5005
R16321 VSS.n4505 VSS.n234 4.5005
R16322 VSS.n4505 VSS.n153 4.5005
R16323 VSS.n4505 VSS.n235 4.5005
R16324 VSS.n4506 VSS.n4505 4.5005
R16325 VSS.n4505 VSS.n236 4.5005
R16326 VSS.n4505 VSS.n152 4.5005
R16327 VSS.n4505 VSS.n237 4.5005
R16328 VSS.n4505 VSS.n151 4.5005
R16329 VSS.n4505 VSS.n238 4.5005
R16330 VSS.n4505 VSS.n150 4.5005
R16331 VSS.n4505 VSS.n239 4.5005
R16332 VSS.n4505 VSS.n149 4.5005
R16333 VSS.n4505 VSS.n240 4.5005
R16334 VSS.n4505 VSS.n148 4.5005
R16335 VSS.n4505 VSS.n241 4.5005
R16336 VSS.n4505 VSS.n147 4.5005
R16337 VSS.n4505 VSS.n242 4.5005
R16338 VSS.n4505 VSS.n146 4.5005
R16339 VSS.n4505 VSS.n243 4.5005
R16340 VSS.n4505 VSS.n145 4.5005
R16341 VSS.n4505 VSS.n244 4.5005
R16342 VSS.n4505 VSS.n144 4.5005
R16343 VSS.n4505 VSS.n245 4.5005
R16344 VSS.n4505 VSS.n143 4.5005
R16345 VSS.n4505 VSS.n246 4.5005
R16346 VSS.n4505 VSS.n142 4.5005
R16347 VSS.n4505 VSS.n247 4.5005
R16348 VSS.n4505 VSS.n141 4.5005
R16349 VSS.n4505 VSS.n248 4.5005
R16350 VSS.n4505 VSS.n140 4.5005
R16351 VSS.n4505 VSS.n249 4.5005
R16352 VSS.n4505 VSS.n139 4.5005
R16353 VSS.n4505 VSS.n250 4.5005
R16354 VSS.n4505 VSS.n138 4.5005
R16355 VSS.n4505 VSS.n251 4.5005
R16356 VSS.n4505 VSS.n137 4.5005
R16357 VSS.n4505 VSS.n252 4.5005
R16358 VSS.n4505 VSS.n136 4.5005
R16359 VSS.n4505 VSS.n253 4.5005
R16360 VSS.n4505 VSS.n135 4.5005
R16361 VSS.n4505 VSS.n254 4.5005
R16362 VSS.n4505 VSS.n134 4.5005
R16363 VSS.n4505 VSS.n255 4.5005
R16364 VSS.n4505 VSS.n133 4.5005
R16365 VSS.n4505 VSS.n256 4.5005
R16366 VSS.n4505 VSS.n132 4.5005
R16367 VSS.n4505 VSS.n4504 4.5005
R16368 VSS.n3051 VSS.n2416 4.5005
R16369 VSS.n3051 VSS.n2415 4.5005
R16370 VSS.n2415 VSS.n2351 4.5005
R16371 VSS.n2483 VSS.n2415 4.5005
R16372 VSS.n2484 VSS.n2415 4.5005
R16373 VSS.n2486 VSS.n2415 4.5005
R16374 VSS.n2489 VSS.n2415 4.5005
R16375 VSS.n2491 VSS.n2415 4.5005
R16376 VSS.n2492 VSS.n2415 4.5005
R16377 VSS.n2494 VSS.n2415 4.5005
R16378 VSS.n2497 VSS.n2415 4.5005
R16379 VSS.n2499 VSS.n2415 4.5005
R16380 VSS.n2500 VSS.n2415 4.5005
R16381 VSS.n2502 VSS.n2415 4.5005
R16382 VSS.n2505 VSS.n2415 4.5005
R16383 VSS.n2507 VSS.n2415 4.5005
R16384 VSS.n2508 VSS.n2415 4.5005
R16385 VSS.n2510 VSS.n2415 4.5005
R16386 VSS.n2513 VSS.n2415 4.5005
R16387 VSS.n2515 VSS.n2415 4.5005
R16388 VSS.n2516 VSS.n2415 4.5005
R16389 VSS.n2518 VSS.n2415 4.5005
R16390 VSS.n2521 VSS.n2415 4.5005
R16391 VSS.n2523 VSS.n2415 4.5005
R16392 VSS.n2524 VSS.n2415 4.5005
R16393 VSS.n2526 VSS.n2415 4.5005
R16394 VSS.n2529 VSS.n2415 4.5005
R16395 VSS.n2531 VSS.n2415 4.5005
R16396 VSS.n2532 VSS.n2415 4.5005
R16397 VSS.n2534 VSS.n2415 4.5005
R16398 VSS.n2537 VSS.n2415 4.5005
R16399 VSS.n2539 VSS.n2415 4.5005
R16400 VSS.n2540 VSS.n2415 4.5005
R16401 VSS.n2542 VSS.n2415 4.5005
R16402 VSS.n2545 VSS.n2415 4.5005
R16403 VSS.n2547 VSS.n2415 4.5005
R16404 VSS.n2548 VSS.n2415 4.5005
R16405 VSS.n2550 VSS.n2415 4.5005
R16406 VSS.n2553 VSS.n2415 4.5005
R16407 VSS.n2555 VSS.n2415 4.5005
R16408 VSS.n2556 VSS.n2415 4.5005
R16409 VSS.n2558 VSS.n2415 4.5005
R16410 VSS.n2561 VSS.n2415 4.5005
R16411 VSS.n2563 VSS.n2415 4.5005
R16412 VSS.n2564 VSS.n2415 4.5005
R16413 VSS.n2566 VSS.n2415 4.5005
R16414 VSS.n2569 VSS.n2415 4.5005
R16415 VSS.n2571 VSS.n2415 4.5005
R16416 VSS.n2572 VSS.n2415 4.5005
R16417 VSS.n2574 VSS.n2415 4.5005
R16418 VSS.n2577 VSS.n2415 4.5005
R16419 VSS.n2579 VSS.n2415 4.5005
R16420 VSS.n2580 VSS.n2415 4.5005
R16421 VSS.n2582 VSS.n2415 4.5005
R16422 VSS.n2585 VSS.n2415 4.5005
R16423 VSS.n2587 VSS.n2415 4.5005
R16424 VSS.n2588 VSS.n2415 4.5005
R16425 VSS.n2590 VSS.n2415 4.5005
R16426 VSS.n2593 VSS.n2415 4.5005
R16427 VSS.n2595 VSS.n2415 4.5005
R16428 VSS.n2596 VSS.n2415 4.5005
R16429 VSS.n2598 VSS.n2415 4.5005
R16430 VSS.n2601 VSS.n2415 4.5005
R16431 VSS.n2603 VSS.n2415 4.5005
R16432 VSS.n2604 VSS.n2415 4.5005
R16433 VSS.n2606 VSS.n2415 4.5005
R16434 VSS.n2609 VSS.n2415 4.5005
R16435 VSS.n2611 VSS.n2415 4.5005
R16436 VSS.n2612 VSS.n2415 4.5005
R16437 VSS.n2614 VSS.n2415 4.5005
R16438 VSS.n2617 VSS.n2415 4.5005
R16439 VSS.n2619 VSS.n2415 4.5005
R16440 VSS.n2620 VSS.n2415 4.5005
R16441 VSS.n2622 VSS.n2415 4.5005
R16442 VSS.n2625 VSS.n2415 4.5005
R16443 VSS.n2627 VSS.n2415 4.5005
R16444 VSS.n2628 VSS.n2415 4.5005
R16445 VSS.n2630 VSS.n2415 4.5005
R16446 VSS.n2633 VSS.n2415 4.5005
R16447 VSS.n2635 VSS.n2415 4.5005
R16448 VSS.n2636 VSS.n2415 4.5005
R16449 VSS.n2638 VSS.n2415 4.5005
R16450 VSS.n2640 VSS.n2415 4.5005
R16451 VSS.n2642 VSS.n2415 4.5005
R16452 VSS.n2643 VSS.n2415 4.5005
R16453 VSS.n2645 VSS.n2415 4.5005
R16454 VSS.n2648 VSS.n2415 4.5005
R16455 VSS.n2650 VSS.n2415 4.5005
R16456 VSS.n2651 VSS.n2415 4.5005
R16457 VSS.n2653 VSS.n2415 4.5005
R16458 VSS.n2656 VSS.n2415 4.5005
R16459 VSS.n2658 VSS.n2415 4.5005
R16460 VSS.n2659 VSS.n2415 4.5005
R16461 VSS.n2661 VSS.n2415 4.5005
R16462 VSS.n2664 VSS.n2415 4.5005
R16463 VSS.n2666 VSS.n2415 4.5005
R16464 VSS.n2667 VSS.n2415 4.5005
R16465 VSS.n2669 VSS.n2415 4.5005
R16466 VSS.n2672 VSS.n2415 4.5005
R16467 VSS.n2674 VSS.n2415 4.5005
R16468 VSS.n2675 VSS.n2415 4.5005
R16469 VSS.n2677 VSS.n2415 4.5005
R16470 VSS.n2680 VSS.n2415 4.5005
R16471 VSS.n2682 VSS.n2415 4.5005
R16472 VSS.n2683 VSS.n2415 4.5005
R16473 VSS.n2685 VSS.n2415 4.5005
R16474 VSS.n2688 VSS.n2415 4.5005
R16475 VSS.n2690 VSS.n2415 4.5005
R16476 VSS.n2691 VSS.n2415 4.5005
R16477 VSS.n2693 VSS.n2415 4.5005
R16478 VSS.n2696 VSS.n2415 4.5005
R16479 VSS.n2698 VSS.n2415 4.5005
R16480 VSS.n2699 VSS.n2415 4.5005
R16481 VSS.n2701 VSS.n2415 4.5005
R16482 VSS.n2704 VSS.n2415 4.5005
R16483 VSS.n2706 VSS.n2415 4.5005
R16484 VSS.n2707 VSS.n2415 4.5005
R16485 VSS.n2709 VSS.n2415 4.5005
R16486 VSS.n2712 VSS.n2415 4.5005
R16487 VSS.n2714 VSS.n2415 4.5005
R16488 VSS.n2715 VSS.n2415 4.5005
R16489 VSS.n2717 VSS.n2415 4.5005
R16490 VSS.n2720 VSS.n2415 4.5005
R16491 VSS.n2722 VSS.n2415 4.5005
R16492 VSS.n2723 VSS.n2415 4.5005
R16493 VSS.n2725 VSS.n2415 4.5005
R16494 VSS.n2793 VSS.n2415 4.5005
R16495 VSS.n2859 VSS.n2415 4.5005
R16496 VSS.n3051 VSS.n2417 4.5005
R16497 VSS.n2417 VSS.n2351 4.5005
R16498 VSS.n2483 VSS.n2417 4.5005
R16499 VSS.n2484 VSS.n2417 4.5005
R16500 VSS.n2486 VSS.n2417 4.5005
R16501 VSS.n2489 VSS.n2417 4.5005
R16502 VSS.n2491 VSS.n2417 4.5005
R16503 VSS.n2492 VSS.n2417 4.5005
R16504 VSS.n2494 VSS.n2417 4.5005
R16505 VSS.n2497 VSS.n2417 4.5005
R16506 VSS.n2499 VSS.n2417 4.5005
R16507 VSS.n2500 VSS.n2417 4.5005
R16508 VSS.n2502 VSS.n2417 4.5005
R16509 VSS.n2505 VSS.n2417 4.5005
R16510 VSS.n2507 VSS.n2417 4.5005
R16511 VSS.n2508 VSS.n2417 4.5005
R16512 VSS.n2510 VSS.n2417 4.5005
R16513 VSS.n2513 VSS.n2417 4.5005
R16514 VSS.n2515 VSS.n2417 4.5005
R16515 VSS.n2516 VSS.n2417 4.5005
R16516 VSS.n2518 VSS.n2417 4.5005
R16517 VSS.n2521 VSS.n2417 4.5005
R16518 VSS.n2523 VSS.n2417 4.5005
R16519 VSS.n2524 VSS.n2417 4.5005
R16520 VSS.n2526 VSS.n2417 4.5005
R16521 VSS.n2529 VSS.n2417 4.5005
R16522 VSS.n2531 VSS.n2417 4.5005
R16523 VSS.n2532 VSS.n2417 4.5005
R16524 VSS.n2534 VSS.n2417 4.5005
R16525 VSS.n2537 VSS.n2417 4.5005
R16526 VSS.n2539 VSS.n2417 4.5005
R16527 VSS.n2540 VSS.n2417 4.5005
R16528 VSS.n2542 VSS.n2417 4.5005
R16529 VSS.n2545 VSS.n2417 4.5005
R16530 VSS.n2547 VSS.n2417 4.5005
R16531 VSS.n2548 VSS.n2417 4.5005
R16532 VSS.n2550 VSS.n2417 4.5005
R16533 VSS.n2553 VSS.n2417 4.5005
R16534 VSS.n2555 VSS.n2417 4.5005
R16535 VSS.n2556 VSS.n2417 4.5005
R16536 VSS.n2558 VSS.n2417 4.5005
R16537 VSS.n2561 VSS.n2417 4.5005
R16538 VSS.n2563 VSS.n2417 4.5005
R16539 VSS.n2564 VSS.n2417 4.5005
R16540 VSS.n2566 VSS.n2417 4.5005
R16541 VSS.n2569 VSS.n2417 4.5005
R16542 VSS.n2571 VSS.n2417 4.5005
R16543 VSS.n2572 VSS.n2417 4.5005
R16544 VSS.n2574 VSS.n2417 4.5005
R16545 VSS.n2577 VSS.n2417 4.5005
R16546 VSS.n2579 VSS.n2417 4.5005
R16547 VSS.n2580 VSS.n2417 4.5005
R16548 VSS.n2582 VSS.n2417 4.5005
R16549 VSS.n2585 VSS.n2417 4.5005
R16550 VSS.n2587 VSS.n2417 4.5005
R16551 VSS.n2588 VSS.n2417 4.5005
R16552 VSS.n2590 VSS.n2417 4.5005
R16553 VSS.n2593 VSS.n2417 4.5005
R16554 VSS.n2595 VSS.n2417 4.5005
R16555 VSS.n2596 VSS.n2417 4.5005
R16556 VSS.n2598 VSS.n2417 4.5005
R16557 VSS.n2601 VSS.n2417 4.5005
R16558 VSS.n2603 VSS.n2417 4.5005
R16559 VSS.n2604 VSS.n2417 4.5005
R16560 VSS.n2606 VSS.n2417 4.5005
R16561 VSS.n2609 VSS.n2417 4.5005
R16562 VSS.n2611 VSS.n2417 4.5005
R16563 VSS.n2612 VSS.n2417 4.5005
R16564 VSS.n2614 VSS.n2417 4.5005
R16565 VSS.n2617 VSS.n2417 4.5005
R16566 VSS.n2619 VSS.n2417 4.5005
R16567 VSS.n2620 VSS.n2417 4.5005
R16568 VSS.n2622 VSS.n2417 4.5005
R16569 VSS.n2625 VSS.n2417 4.5005
R16570 VSS.n2627 VSS.n2417 4.5005
R16571 VSS.n2628 VSS.n2417 4.5005
R16572 VSS.n2630 VSS.n2417 4.5005
R16573 VSS.n2633 VSS.n2417 4.5005
R16574 VSS.n2635 VSS.n2417 4.5005
R16575 VSS.n2636 VSS.n2417 4.5005
R16576 VSS.n2638 VSS.n2417 4.5005
R16577 VSS.n2640 VSS.n2417 4.5005
R16578 VSS.n2642 VSS.n2417 4.5005
R16579 VSS.n2643 VSS.n2417 4.5005
R16580 VSS.n2645 VSS.n2417 4.5005
R16581 VSS.n2648 VSS.n2417 4.5005
R16582 VSS.n2650 VSS.n2417 4.5005
R16583 VSS.n2651 VSS.n2417 4.5005
R16584 VSS.n2653 VSS.n2417 4.5005
R16585 VSS.n2656 VSS.n2417 4.5005
R16586 VSS.n2658 VSS.n2417 4.5005
R16587 VSS.n2659 VSS.n2417 4.5005
R16588 VSS.n2661 VSS.n2417 4.5005
R16589 VSS.n2664 VSS.n2417 4.5005
R16590 VSS.n2666 VSS.n2417 4.5005
R16591 VSS.n2667 VSS.n2417 4.5005
R16592 VSS.n2669 VSS.n2417 4.5005
R16593 VSS.n2672 VSS.n2417 4.5005
R16594 VSS.n2674 VSS.n2417 4.5005
R16595 VSS.n2675 VSS.n2417 4.5005
R16596 VSS.n2677 VSS.n2417 4.5005
R16597 VSS.n2680 VSS.n2417 4.5005
R16598 VSS.n2682 VSS.n2417 4.5005
R16599 VSS.n2683 VSS.n2417 4.5005
R16600 VSS.n2685 VSS.n2417 4.5005
R16601 VSS.n2688 VSS.n2417 4.5005
R16602 VSS.n2690 VSS.n2417 4.5005
R16603 VSS.n2691 VSS.n2417 4.5005
R16604 VSS.n2693 VSS.n2417 4.5005
R16605 VSS.n2696 VSS.n2417 4.5005
R16606 VSS.n2698 VSS.n2417 4.5005
R16607 VSS.n2699 VSS.n2417 4.5005
R16608 VSS.n2701 VSS.n2417 4.5005
R16609 VSS.n2704 VSS.n2417 4.5005
R16610 VSS.n2706 VSS.n2417 4.5005
R16611 VSS.n2707 VSS.n2417 4.5005
R16612 VSS.n2709 VSS.n2417 4.5005
R16613 VSS.n2712 VSS.n2417 4.5005
R16614 VSS.n2714 VSS.n2417 4.5005
R16615 VSS.n2715 VSS.n2417 4.5005
R16616 VSS.n2717 VSS.n2417 4.5005
R16617 VSS.n2720 VSS.n2417 4.5005
R16618 VSS.n2722 VSS.n2417 4.5005
R16619 VSS.n2723 VSS.n2417 4.5005
R16620 VSS.n2725 VSS.n2417 4.5005
R16621 VSS.n2793 VSS.n2417 4.5005
R16622 VSS.n2859 VSS.n2417 4.5005
R16623 VSS.n3051 VSS.n2414 4.5005
R16624 VSS.n2414 VSS.n2351 4.5005
R16625 VSS.n2483 VSS.n2414 4.5005
R16626 VSS.n2484 VSS.n2414 4.5005
R16627 VSS.n2486 VSS.n2414 4.5005
R16628 VSS.n2489 VSS.n2414 4.5005
R16629 VSS.n2491 VSS.n2414 4.5005
R16630 VSS.n2492 VSS.n2414 4.5005
R16631 VSS.n2494 VSS.n2414 4.5005
R16632 VSS.n2497 VSS.n2414 4.5005
R16633 VSS.n2499 VSS.n2414 4.5005
R16634 VSS.n2500 VSS.n2414 4.5005
R16635 VSS.n2502 VSS.n2414 4.5005
R16636 VSS.n2505 VSS.n2414 4.5005
R16637 VSS.n2507 VSS.n2414 4.5005
R16638 VSS.n2508 VSS.n2414 4.5005
R16639 VSS.n2510 VSS.n2414 4.5005
R16640 VSS.n2513 VSS.n2414 4.5005
R16641 VSS.n2515 VSS.n2414 4.5005
R16642 VSS.n2516 VSS.n2414 4.5005
R16643 VSS.n2518 VSS.n2414 4.5005
R16644 VSS.n2521 VSS.n2414 4.5005
R16645 VSS.n2523 VSS.n2414 4.5005
R16646 VSS.n2524 VSS.n2414 4.5005
R16647 VSS.n2526 VSS.n2414 4.5005
R16648 VSS.n2529 VSS.n2414 4.5005
R16649 VSS.n2531 VSS.n2414 4.5005
R16650 VSS.n2532 VSS.n2414 4.5005
R16651 VSS.n2534 VSS.n2414 4.5005
R16652 VSS.n2537 VSS.n2414 4.5005
R16653 VSS.n2539 VSS.n2414 4.5005
R16654 VSS.n2540 VSS.n2414 4.5005
R16655 VSS.n2542 VSS.n2414 4.5005
R16656 VSS.n2545 VSS.n2414 4.5005
R16657 VSS.n2547 VSS.n2414 4.5005
R16658 VSS.n2548 VSS.n2414 4.5005
R16659 VSS.n2550 VSS.n2414 4.5005
R16660 VSS.n2553 VSS.n2414 4.5005
R16661 VSS.n2555 VSS.n2414 4.5005
R16662 VSS.n2556 VSS.n2414 4.5005
R16663 VSS.n2558 VSS.n2414 4.5005
R16664 VSS.n2561 VSS.n2414 4.5005
R16665 VSS.n2563 VSS.n2414 4.5005
R16666 VSS.n2564 VSS.n2414 4.5005
R16667 VSS.n2566 VSS.n2414 4.5005
R16668 VSS.n2569 VSS.n2414 4.5005
R16669 VSS.n2571 VSS.n2414 4.5005
R16670 VSS.n2572 VSS.n2414 4.5005
R16671 VSS.n2574 VSS.n2414 4.5005
R16672 VSS.n2577 VSS.n2414 4.5005
R16673 VSS.n2579 VSS.n2414 4.5005
R16674 VSS.n2580 VSS.n2414 4.5005
R16675 VSS.n2582 VSS.n2414 4.5005
R16676 VSS.n2585 VSS.n2414 4.5005
R16677 VSS.n2587 VSS.n2414 4.5005
R16678 VSS.n2588 VSS.n2414 4.5005
R16679 VSS.n2590 VSS.n2414 4.5005
R16680 VSS.n2593 VSS.n2414 4.5005
R16681 VSS.n2595 VSS.n2414 4.5005
R16682 VSS.n2596 VSS.n2414 4.5005
R16683 VSS.n2598 VSS.n2414 4.5005
R16684 VSS.n2601 VSS.n2414 4.5005
R16685 VSS.n2603 VSS.n2414 4.5005
R16686 VSS.n2604 VSS.n2414 4.5005
R16687 VSS.n2606 VSS.n2414 4.5005
R16688 VSS.n2609 VSS.n2414 4.5005
R16689 VSS.n2611 VSS.n2414 4.5005
R16690 VSS.n2612 VSS.n2414 4.5005
R16691 VSS.n2614 VSS.n2414 4.5005
R16692 VSS.n2617 VSS.n2414 4.5005
R16693 VSS.n2619 VSS.n2414 4.5005
R16694 VSS.n2620 VSS.n2414 4.5005
R16695 VSS.n2622 VSS.n2414 4.5005
R16696 VSS.n2625 VSS.n2414 4.5005
R16697 VSS.n2627 VSS.n2414 4.5005
R16698 VSS.n2628 VSS.n2414 4.5005
R16699 VSS.n2630 VSS.n2414 4.5005
R16700 VSS.n2633 VSS.n2414 4.5005
R16701 VSS.n2635 VSS.n2414 4.5005
R16702 VSS.n2636 VSS.n2414 4.5005
R16703 VSS.n2638 VSS.n2414 4.5005
R16704 VSS.n2640 VSS.n2414 4.5005
R16705 VSS.n2642 VSS.n2414 4.5005
R16706 VSS.n2643 VSS.n2414 4.5005
R16707 VSS.n2645 VSS.n2414 4.5005
R16708 VSS.n2648 VSS.n2414 4.5005
R16709 VSS.n2650 VSS.n2414 4.5005
R16710 VSS.n2651 VSS.n2414 4.5005
R16711 VSS.n2653 VSS.n2414 4.5005
R16712 VSS.n2656 VSS.n2414 4.5005
R16713 VSS.n2658 VSS.n2414 4.5005
R16714 VSS.n2659 VSS.n2414 4.5005
R16715 VSS.n2661 VSS.n2414 4.5005
R16716 VSS.n2664 VSS.n2414 4.5005
R16717 VSS.n2666 VSS.n2414 4.5005
R16718 VSS.n2667 VSS.n2414 4.5005
R16719 VSS.n2669 VSS.n2414 4.5005
R16720 VSS.n2672 VSS.n2414 4.5005
R16721 VSS.n2674 VSS.n2414 4.5005
R16722 VSS.n2675 VSS.n2414 4.5005
R16723 VSS.n2677 VSS.n2414 4.5005
R16724 VSS.n2680 VSS.n2414 4.5005
R16725 VSS.n2682 VSS.n2414 4.5005
R16726 VSS.n2683 VSS.n2414 4.5005
R16727 VSS.n2685 VSS.n2414 4.5005
R16728 VSS.n2688 VSS.n2414 4.5005
R16729 VSS.n2690 VSS.n2414 4.5005
R16730 VSS.n2691 VSS.n2414 4.5005
R16731 VSS.n2693 VSS.n2414 4.5005
R16732 VSS.n2696 VSS.n2414 4.5005
R16733 VSS.n2698 VSS.n2414 4.5005
R16734 VSS.n2699 VSS.n2414 4.5005
R16735 VSS.n2701 VSS.n2414 4.5005
R16736 VSS.n2704 VSS.n2414 4.5005
R16737 VSS.n2706 VSS.n2414 4.5005
R16738 VSS.n2707 VSS.n2414 4.5005
R16739 VSS.n2709 VSS.n2414 4.5005
R16740 VSS.n2712 VSS.n2414 4.5005
R16741 VSS.n2714 VSS.n2414 4.5005
R16742 VSS.n2715 VSS.n2414 4.5005
R16743 VSS.n2717 VSS.n2414 4.5005
R16744 VSS.n2720 VSS.n2414 4.5005
R16745 VSS.n2722 VSS.n2414 4.5005
R16746 VSS.n2723 VSS.n2414 4.5005
R16747 VSS.n2725 VSS.n2414 4.5005
R16748 VSS.n2793 VSS.n2414 4.5005
R16749 VSS.n2859 VSS.n2414 4.5005
R16750 VSS.n3051 VSS.n2418 4.5005
R16751 VSS.n2418 VSS.n2351 4.5005
R16752 VSS.n2483 VSS.n2418 4.5005
R16753 VSS.n2484 VSS.n2418 4.5005
R16754 VSS.n2486 VSS.n2418 4.5005
R16755 VSS.n2489 VSS.n2418 4.5005
R16756 VSS.n2491 VSS.n2418 4.5005
R16757 VSS.n2492 VSS.n2418 4.5005
R16758 VSS.n2494 VSS.n2418 4.5005
R16759 VSS.n2497 VSS.n2418 4.5005
R16760 VSS.n2499 VSS.n2418 4.5005
R16761 VSS.n2500 VSS.n2418 4.5005
R16762 VSS.n2502 VSS.n2418 4.5005
R16763 VSS.n2505 VSS.n2418 4.5005
R16764 VSS.n2507 VSS.n2418 4.5005
R16765 VSS.n2508 VSS.n2418 4.5005
R16766 VSS.n2510 VSS.n2418 4.5005
R16767 VSS.n2513 VSS.n2418 4.5005
R16768 VSS.n2515 VSS.n2418 4.5005
R16769 VSS.n2516 VSS.n2418 4.5005
R16770 VSS.n2518 VSS.n2418 4.5005
R16771 VSS.n2521 VSS.n2418 4.5005
R16772 VSS.n2523 VSS.n2418 4.5005
R16773 VSS.n2524 VSS.n2418 4.5005
R16774 VSS.n2526 VSS.n2418 4.5005
R16775 VSS.n2529 VSS.n2418 4.5005
R16776 VSS.n2531 VSS.n2418 4.5005
R16777 VSS.n2532 VSS.n2418 4.5005
R16778 VSS.n2534 VSS.n2418 4.5005
R16779 VSS.n2537 VSS.n2418 4.5005
R16780 VSS.n2539 VSS.n2418 4.5005
R16781 VSS.n2540 VSS.n2418 4.5005
R16782 VSS.n2542 VSS.n2418 4.5005
R16783 VSS.n2545 VSS.n2418 4.5005
R16784 VSS.n2547 VSS.n2418 4.5005
R16785 VSS.n2548 VSS.n2418 4.5005
R16786 VSS.n2550 VSS.n2418 4.5005
R16787 VSS.n2553 VSS.n2418 4.5005
R16788 VSS.n2555 VSS.n2418 4.5005
R16789 VSS.n2556 VSS.n2418 4.5005
R16790 VSS.n2558 VSS.n2418 4.5005
R16791 VSS.n2561 VSS.n2418 4.5005
R16792 VSS.n2563 VSS.n2418 4.5005
R16793 VSS.n2564 VSS.n2418 4.5005
R16794 VSS.n2566 VSS.n2418 4.5005
R16795 VSS.n2569 VSS.n2418 4.5005
R16796 VSS.n2571 VSS.n2418 4.5005
R16797 VSS.n2572 VSS.n2418 4.5005
R16798 VSS.n2574 VSS.n2418 4.5005
R16799 VSS.n2577 VSS.n2418 4.5005
R16800 VSS.n2579 VSS.n2418 4.5005
R16801 VSS.n2580 VSS.n2418 4.5005
R16802 VSS.n2582 VSS.n2418 4.5005
R16803 VSS.n2585 VSS.n2418 4.5005
R16804 VSS.n2587 VSS.n2418 4.5005
R16805 VSS.n2588 VSS.n2418 4.5005
R16806 VSS.n2590 VSS.n2418 4.5005
R16807 VSS.n2593 VSS.n2418 4.5005
R16808 VSS.n2595 VSS.n2418 4.5005
R16809 VSS.n2596 VSS.n2418 4.5005
R16810 VSS.n2598 VSS.n2418 4.5005
R16811 VSS.n2601 VSS.n2418 4.5005
R16812 VSS.n2603 VSS.n2418 4.5005
R16813 VSS.n2604 VSS.n2418 4.5005
R16814 VSS.n2606 VSS.n2418 4.5005
R16815 VSS.n2609 VSS.n2418 4.5005
R16816 VSS.n2611 VSS.n2418 4.5005
R16817 VSS.n2612 VSS.n2418 4.5005
R16818 VSS.n2614 VSS.n2418 4.5005
R16819 VSS.n2617 VSS.n2418 4.5005
R16820 VSS.n2619 VSS.n2418 4.5005
R16821 VSS.n2620 VSS.n2418 4.5005
R16822 VSS.n2622 VSS.n2418 4.5005
R16823 VSS.n2625 VSS.n2418 4.5005
R16824 VSS.n2627 VSS.n2418 4.5005
R16825 VSS.n2628 VSS.n2418 4.5005
R16826 VSS.n2630 VSS.n2418 4.5005
R16827 VSS.n2633 VSS.n2418 4.5005
R16828 VSS.n2635 VSS.n2418 4.5005
R16829 VSS.n2636 VSS.n2418 4.5005
R16830 VSS.n2638 VSS.n2418 4.5005
R16831 VSS.n2640 VSS.n2418 4.5005
R16832 VSS.n2642 VSS.n2418 4.5005
R16833 VSS.n2643 VSS.n2418 4.5005
R16834 VSS.n2645 VSS.n2418 4.5005
R16835 VSS.n2648 VSS.n2418 4.5005
R16836 VSS.n2650 VSS.n2418 4.5005
R16837 VSS.n2651 VSS.n2418 4.5005
R16838 VSS.n2653 VSS.n2418 4.5005
R16839 VSS.n2656 VSS.n2418 4.5005
R16840 VSS.n2658 VSS.n2418 4.5005
R16841 VSS.n2659 VSS.n2418 4.5005
R16842 VSS.n2661 VSS.n2418 4.5005
R16843 VSS.n2664 VSS.n2418 4.5005
R16844 VSS.n2666 VSS.n2418 4.5005
R16845 VSS.n2667 VSS.n2418 4.5005
R16846 VSS.n2669 VSS.n2418 4.5005
R16847 VSS.n2672 VSS.n2418 4.5005
R16848 VSS.n2674 VSS.n2418 4.5005
R16849 VSS.n2675 VSS.n2418 4.5005
R16850 VSS.n2677 VSS.n2418 4.5005
R16851 VSS.n2680 VSS.n2418 4.5005
R16852 VSS.n2682 VSS.n2418 4.5005
R16853 VSS.n2683 VSS.n2418 4.5005
R16854 VSS.n2685 VSS.n2418 4.5005
R16855 VSS.n2688 VSS.n2418 4.5005
R16856 VSS.n2690 VSS.n2418 4.5005
R16857 VSS.n2691 VSS.n2418 4.5005
R16858 VSS.n2693 VSS.n2418 4.5005
R16859 VSS.n2696 VSS.n2418 4.5005
R16860 VSS.n2698 VSS.n2418 4.5005
R16861 VSS.n2699 VSS.n2418 4.5005
R16862 VSS.n2701 VSS.n2418 4.5005
R16863 VSS.n2704 VSS.n2418 4.5005
R16864 VSS.n2706 VSS.n2418 4.5005
R16865 VSS.n2707 VSS.n2418 4.5005
R16866 VSS.n2709 VSS.n2418 4.5005
R16867 VSS.n2712 VSS.n2418 4.5005
R16868 VSS.n2714 VSS.n2418 4.5005
R16869 VSS.n2715 VSS.n2418 4.5005
R16870 VSS.n2717 VSS.n2418 4.5005
R16871 VSS.n2720 VSS.n2418 4.5005
R16872 VSS.n2722 VSS.n2418 4.5005
R16873 VSS.n2723 VSS.n2418 4.5005
R16874 VSS.n2725 VSS.n2418 4.5005
R16875 VSS.n2793 VSS.n2418 4.5005
R16876 VSS.n2859 VSS.n2418 4.5005
R16877 VSS.n3051 VSS.n2413 4.5005
R16878 VSS.n2413 VSS.n2351 4.5005
R16879 VSS.n2483 VSS.n2413 4.5005
R16880 VSS.n2484 VSS.n2413 4.5005
R16881 VSS.n2486 VSS.n2413 4.5005
R16882 VSS.n2489 VSS.n2413 4.5005
R16883 VSS.n2491 VSS.n2413 4.5005
R16884 VSS.n2492 VSS.n2413 4.5005
R16885 VSS.n2494 VSS.n2413 4.5005
R16886 VSS.n2497 VSS.n2413 4.5005
R16887 VSS.n2499 VSS.n2413 4.5005
R16888 VSS.n2500 VSS.n2413 4.5005
R16889 VSS.n2502 VSS.n2413 4.5005
R16890 VSS.n2505 VSS.n2413 4.5005
R16891 VSS.n2507 VSS.n2413 4.5005
R16892 VSS.n2508 VSS.n2413 4.5005
R16893 VSS.n2510 VSS.n2413 4.5005
R16894 VSS.n2513 VSS.n2413 4.5005
R16895 VSS.n2515 VSS.n2413 4.5005
R16896 VSS.n2516 VSS.n2413 4.5005
R16897 VSS.n2518 VSS.n2413 4.5005
R16898 VSS.n2521 VSS.n2413 4.5005
R16899 VSS.n2523 VSS.n2413 4.5005
R16900 VSS.n2524 VSS.n2413 4.5005
R16901 VSS.n2526 VSS.n2413 4.5005
R16902 VSS.n2529 VSS.n2413 4.5005
R16903 VSS.n2531 VSS.n2413 4.5005
R16904 VSS.n2532 VSS.n2413 4.5005
R16905 VSS.n2534 VSS.n2413 4.5005
R16906 VSS.n2537 VSS.n2413 4.5005
R16907 VSS.n2539 VSS.n2413 4.5005
R16908 VSS.n2540 VSS.n2413 4.5005
R16909 VSS.n2542 VSS.n2413 4.5005
R16910 VSS.n2545 VSS.n2413 4.5005
R16911 VSS.n2547 VSS.n2413 4.5005
R16912 VSS.n2548 VSS.n2413 4.5005
R16913 VSS.n2550 VSS.n2413 4.5005
R16914 VSS.n2553 VSS.n2413 4.5005
R16915 VSS.n2555 VSS.n2413 4.5005
R16916 VSS.n2556 VSS.n2413 4.5005
R16917 VSS.n2558 VSS.n2413 4.5005
R16918 VSS.n2561 VSS.n2413 4.5005
R16919 VSS.n2563 VSS.n2413 4.5005
R16920 VSS.n2564 VSS.n2413 4.5005
R16921 VSS.n2566 VSS.n2413 4.5005
R16922 VSS.n2569 VSS.n2413 4.5005
R16923 VSS.n2571 VSS.n2413 4.5005
R16924 VSS.n2572 VSS.n2413 4.5005
R16925 VSS.n2574 VSS.n2413 4.5005
R16926 VSS.n2577 VSS.n2413 4.5005
R16927 VSS.n2579 VSS.n2413 4.5005
R16928 VSS.n2580 VSS.n2413 4.5005
R16929 VSS.n2582 VSS.n2413 4.5005
R16930 VSS.n2585 VSS.n2413 4.5005
R16931 VSS.n2587 VSS.n2413 4.5005
R16932 VSS.n2588 VSS.n2413 4.5005
R16933 VSS.n2590 VSS.n2413 4.5005
R16934 VSS.n2593 VSS.n2413 4.5005
R16935 VSS.n2595 VSS.n2413 4.5005
R16936 VSS.n2596 VSS.n2413 4.5005
R16937 VSS.n2598 VSS.n2413 4.5005
R16938 VSS.n2601 VSS.n2413 4.5005
R16939 VSS.n2603 VSS.n2413 4.5005
R16940 VSS.n2604 VSS.n2413 4.5005
R16941 VSS.n2606 VSS.n2413 4.5005
R16942 VSS.n2609 VSS.n2413 4.5005
R16943 VSS.n2611 VSS.n2413 4.5005
R16944 VSS.n2612 VSS.n2413 4.5005
R16945 VSS.n2614 VSS.n2413 4.5005
R16946 VSS.n2617 VSS.n2413 4.5005
R16947 VSS.n2619 VSS.n2413 4.5005
R16948 VSS.n2620 VSS.n2413 4.5005
R16949 VSS.n2622 VSS.n2413 4.5005
R16950 VSS.n2625 VSS.n2413 4.5005
R16951 VSS.n2627 VSS.n2413 4.5005
R16952 VSS.n2628 VSS.n2413 4.5005
R16953 VSS.n2630 VSS.n2413 4.5005
R16954 VSS.n2633 VSS.n2413 4.5005
R16955 VSS.n2635 VSS.n2413 4.5005
R16956 VSS.n2636 VSS.n2413 4.5005
R16957 VSS.n2638 VSS.n2413 4.5005
R16958 VSS.n2640 VSS.n2413 4.5005
R16959 VSS.n2642 VSS.n2413 4.5005
R16960 VSS.n2643 VSS.n2413 4.5005
R16961 VSS.n2645 VSS.n2413 4.5005
R16962 VSS.n2648 VSS.n2413 4.5005
R16963 VSS.n2650 VSS.n2413 4.5005
R16964 VSS.n2651 VSS.n2413 4.5005
R16965 VSS.n2653 VSS.n2413 4.5005
R16966 VSS.n2656 VSS.n2413 4.5005
R16967 VSS.n2658 VSS.n2413 4.5005
R16968 VSS.n2659 VSS.n2413 4.5005
R16969 VSS.n2661 VSS.n2413 4.5005
R16970 VSS.n2664 VSS.n2413 4.5005
R16971 VSS.n2666 VSS.n2413 4.5005
R16972 VSS.n2667 VSS.n2413 4.5005
R16973 VSS.n2669 VSS.n2413 4.5005
R16974 VSS.n2672 VSS.n2413 4.5005
R16975 VSS.n2674 VSS.n2413 4.5005
R16976 VSS.n2675 VSS.n2413 4.5005
R16977 VSS.n2677 VSS.n2413 4.5005
R16978 VSS.n2680 VSS.n2413 4.5005
R16979 VSS.n2682 VSS.n2413 4.5005
R16980 VSS.n2683 VSS.n2413 4.5005
R16981 VSS.n2685 VSS.n2413 4.5005
R16982 VSS.n2688 VSS.n2413 4.5005
R16983 VSS.n2690 VSS.n2413 4.5005
R16984 VSS.n2691 VSS.n2413 4.5005
R16985 VSS.n2693 VSS.n2413 4.5005
R16986 VSS.n2696 VSS.n2413 4.5005
R16987 VSS.n2698 VSS.n2413 4.5005
R16988 VSS.n2699 VSS.n2413 4.5005
R16989 VSS.n2701 VSS.n2413 4.5005
R16990 VSS.n2704 VSS.n2413 4.5005
R16991 VSS.n2706 VSS.n2413 4.5005
R16992 VSS.n2707 VSS.n2413 4.5005
R16993 VSS.n2709 VSS.n2413 4.5005
R16994 VSS.n2712 VSS.n2413 4.5005
R16995 VSS.n2714 VSS.n2413 4.5005
R16996 VSS.n2715 VSS.n2413 4.5005
R16997 VSS.n2717 VSS.n2413 4.5005
R16998 VSS.n2720 VSS.n2413 4.5005
R16999 VSS.n2722 VSS.n2413 4.5005
R17000 VSS.n2723 VSS.n2413 4.5005
R17001 VSS.n2725 VSS.n2413 4.5005
R17002 VSS.n2793 VSS.n2413 4.5005
R17003 VSS.n2859 VSS.n2413 4.5005
R17004 VSS.n3051 VSS.n2419 4.5005
R17005 VSS.n2419 VSS.n2351 4.5005
R17006 VSS.n2483 VSS.n2419 4.5005
R17007 VSS.n2484 VSS.n2419 4.5005
R17008 VSS.n2486 VSS.n2419 4.5005
R17009 VSS.n2489 VSS.n2419 4.5005
R17010 VSS.n2491 VSS.n2419 4.5005
R17011 VSS.n2492 VSS.n2419 4.5005
R17012 VSS.n2494 VSS.n2419 4.5005
R17013 VSS.n2497 VSS.n2419 4.5005
R17014 VSS.n2499 VSS.n2419 4.5005
R17015 VSS.n2500 VSS.n2419 4.5005
R17016 VSS.n2502 VSS.n2419 4.5005
R17017 VSS.n2505 VSS.n2419 4.5005
R17018 VSS.n2507 VSS.n2419 4.5005
R17019 VSS.n2508 VSS.n2419 4.5005
R17020 VSS.n2510 VSS.n2419 4.5005
R17021 VSS.n2513 VSS.n2419 4.5005
R17022 VSS.n2515 VSS.n2419 4.5005
R17023 VSS.n2516 VSS.n2419 4.5005
R17024 VSS.n2518 VSS.n2419 4.5005
R17025 VSS.n2521 VSS.n2419 4.5005
R17026 VSS.n2523 VSS.n2419 4.5005
R17027 VSS.n2524 VSS.n2419 4.5005
R17028 VSS.n2526 VSS.n2419 4.5005
R17029 VSS.n2529 VSS.n2419 4.5005
R17030 VSS.n2531 VSS.n2419 4.5005
R17031 VSS.n2532 VSS.n2419 4.5005
R17032 VSS.n2534 VSS.n2419 4.5005
R17033 VSS.n2537 VSS.n2419 4.5005
R17034 VSS.n2539 VSS.n2419 4.5005
R17035 VSS.n2540 VSS.n2419 4.5005
R17036 VSS.n2542 VSS.n2419 4.5005
R17037 VSS.n2545 VSS.n2419 4.5005
R17038 VSS.n2547 VSS.n2419 4.5005
R17039 VSS.n2548 VSS.n2419 4.5005
R17040 VSS.n2550 VSS.n2419 4.5005
R17041 VSS.n2553 VSS.n2419 4.5005
R17042 VSS.n2555 VSS.n2419 4.5005
R17043 VSS.n2556 VSS.n2419 4.5005
R17044 VSS.n2558 VSS.n2419 4.5005
R17045 VSS.n2561 VSS.n2419 4.5005
R17046 VSS.n2563 VSS.n2419 4.5005
R17047 VSS.n2564 VSS.n2419 4.5005
R17048 VSS.n2566 VSS.n2419 4.5005
R17049 VSS.n2569 VSS.n2419 4.5005
R17050 VSS.n2571 VSS.n2419 4.5005
R17051 VSS.n2572 VSS.n2419 4.5005
R17052 VSS.n2574 VSS.n2419 4.5005
R17053 VSS.n2577 VSS.n2419 4.5005
R17054 VSS.n2579 VSS.n2419 4.5005
R17055 VSS.n2580 VSS.n2419 4.5005
R17056 VSS.n2582 VSS.n2419 4.5005
R17057 VSS.n2585 VSS.n2419 4.5005
R17058 VSS.n2587 VSS.n2419 4.5005
R17059 VSS.n2588 VSS.n2419 4.5005
R17060 VSS.n2590 VSS.n2419 4.5005
R17061 VSS.n2593 VSS.n2419 4.5005
R17062 VSS.n2595 VSS.n2419 4.5005
R17063 VSS.n2596 VSS.n2419 4.5005
R17064 VSS.n2598 VSS.n2419 4.5005
R17065 VSS.n2601 VSS.n2419 4.5005
R17066 VSS.n2603 VSS.n2419 4.5005
R17067 VSS.n2604 VSS.n2419 4.5005
R17068 VSS.n2606 VSS.n2419 4.5005
R17069 VSS.n2609 VSS.n2419 4.5005
R17070 VSS.n2611 VSS.n2419 4.5005
R17071 VSS.n2612 VSS.n2419 4.5005
R17072 VSS.n2614 VSS.n2419 4.5005
R17073 VSS.n2617 VSS.n2419 4.5005
R17074 VSS.n2619 VSS.n2419 4.5005
R17075 VSS.n2620 VSS.n2419 4.5005
R17076 VSS.n2622 VSS.n2419 4.5005
R17077 VSS.n2625 VSS.n2419 4.5005
R17078 VSS.n2627 VSS.n2419 4.5005
R17079 VSS.n2628 VSS.n2419 4.5005
R17080 VSS.n2630 VSS.n2419 4.5005
R17081 VSS.n2633 VSS.n2419 4.5005
R17082 VSS.n2635 VSS.n2419 4.5005
R17083 VSS.n2636 VSS.n2419 4.5005
R17084 VSS.n2638 VSS.n2419 4.5005
R17085 VSS.n2640 VSS.n2419 4.5005
R17086 VSS.n2642 VSS.n2419 4.5005
R17087 VSS.n2643 VSS.n2419 4.5005
R17088 VSS.n2645 VSS.n2419 4.5005
R17089 VSS.n2648 VSS.n2419 4.5005
R17090 VSS.n2650 VSS.n2419 4.5005
R17091 VSS.n2651 VSS.n2419 4.5005
R17092 VSS.n2653 VSS.n2419 4.5005
R17093 VSS.n2656 VSS.n2419 4.5005
R17094 VSS.n2658 VSS.n2419 4.5005
R17095 VSS.n2659 VSS.n2419 4.5005
R17096 VSS.n2661 VSS.n2419 4.5005
R17097 VSS.n2664 VSS.n2419 4.5005
R17098 VSS.n2666 VSS.n2419 4.5005
R17099 VSS.n2667 VSS.n2419 4.5005
R17100 VSS.n2669 VSS.n2419 4.5005
R17101 VSS.n2672 VSS.n2419 4.5005
R17102 VSS.n2674 VSS.n2419 4.5005
R17103 VSS.n2675 VSS.n2419 4.5005
R17104 VSS.n2677 VSS.n2419 4.5005
R17105 VSS.n2680 VSS.n2419 4.5005
R17106 VSS.n2682 VSS.n2419 4.5005
R17107 VSS.n2683 VSS.n2419 4.5005
R17108 VSS.n2685 VSS.n2419 4.5005
R17109 VSS.n2688 VSS.n2419 4.5005
R17110 VSS.n2690 VSS.n2419 4.5005
R17111 VSS.n2691 VSS.n2419 4.5005
R17112 VSS.n2693 VSS.n2419 4.5005
R17113 VSS.n2696 VSS.n2419 4.5005
R17114 VSS.n2698 VSS.n2419 4.5005
R17115 VSS.n2699 VSS.n2419 4.5005
R17116 VSS.n2701 VSS.n2419 4.5005
R17117 VSS.n2704 VSS.n2419 4.5005
R17118 VSS.n2706 VSS.n2419 4.5005
R17119 VSS.n2707 VSS.n2419 4.5005
R17120 VSS.n2709 VSS.n2419 4.5005
R17121 VSS.n2712 VSS.n2419 4.5005
R17122 VSS.n2714 VSS.n2419 4.5005
R17123 VSS.n2715 VSS.n2419 4.5005
R17124 VSS.n2717 VSS.n2419 4.5005
R17125 VSS.n2720 VSS.n2419 4.5005
R17126 VSS.n2722 VSS.n2419 4.5005
R17127 VSS.n2723 VSS.n2419 4.5005
R17128 VSS.n2725 VSS.n2419 4.5005
R17129 VSS.n2793 VSS.n2419 4.5005
R17130 VSS.n2859 VSS.n2419 4.5005
R17131 VSS.n3051 VSS.n2412 4.5005
R17132 VSS.n2412 VSS.n2351 4.5005
R17133 VSS.n2483 VSS.n2412 4.5005
R17134 VSS.n2484 VSS.n2412 4.5005
R17135 VSS.n2486 VSS.n2412 4.5005
R17136 VSS.n2489 VSS.n2412 4.5005
R17137 VSS.n2491 VSS.n2412 4.5005
R17138 VSS.n2492 VSS.n2412 4.5005
R17139 VSS.n2494 VSS.n2412 4.5005
R17140 VSS.n2497 VSS.n2412 4.5005
R17141 VSS.n2499 VSS.n2412 4.5005
R17142 VSS.n2500 VSS.n2412 4.5005
R17143 VSS.n2502 VSS.n2412 4.5005
R17144 VSS.n2505 VSS.n2412 4.5005
R17145 VSS.n2507 VSS.n2412 4.5005
R17146 VSS.n2508 VSS.n2412 4.5005
R17147 VSS.n2510 VSS.n2412 4.5005
R17148 VSS.n2513 VSS.n2412 4.5005
R17149 VSS.n2515 VSS.n2412 4.5005
R17150 VSS.n2516 VSS.n2412 4.5005
R17151 VSS.n2518 VSS.n2412 4.5005
R17152 VSS.n2521 VSS.n2412 4.5005
R17153 VSS.n2523 VSS.n2412 4.5005
R17154 VSS.n2524 VSS.n2412 4.5005
R17155 VSS.n2526 VSS.n2412 4.5005
R17156 VSS.n2529 VSS.n2412 4.5005
R17157 VSS.n2531 VSS.n2412 4.5005
R17158 VSS.n2532 VSS.n2412 4.5005
R17159 VSS.n2534 VSS.n2412 4.5005
R17160 VSS.n2537 VSS.n2412 4.5005
R17161 VSS.n2539 VSS.n2412 4.5005
R17162 VSS.n2540 VSS.n2412 4.5005
R17163 VSS.n2542 VSS.n2412 4.5005
R17164 VSS.n2545 VSS.n2412 4.5005
R17165 VSS.n2547 VSS.n2412 4.5005
R17166 VSS.n2548 VSS.n2412 4.5005
R17167 VSS.n2550 VSS.n2412 4.5005
R17168 VSS.n2553 VSS.n2412 4.5005
R17169 VSS.n2555 VSS.n2412 4.5005
R17170 VSS.n2556 VSS.n2412 4.5005
R17171 VSS.n2558 VSS.n2412 4.5005
R17172 VSS.n2561 VSS.n2412 4.5005
R17173 VSS.n2563 VSS.n2412 4.5005
R17174 VSS.n2564 VSS.n2412 4.5005
R17175 VSS.n2566 VSS.n2412 4.5005
R17176 VSS.n2569 VSS.n2412 4.5005
R17177 VSS.n2571 VSS.n2412 4.5005
R17178 VSS.n2572 VSS.n2412 4.5005
R17179 VSS.n2574 VSS.n2412 4.5005
R17180 VSS.n2577 VSS.n2412 4.5005
R17181 VSS.n2579 VSS.n2412 4.5005
R17182 VSS.n2580 VSS.n2412 4.5005
R17183 VSS.n2582 VSS.n2412 4.5005
R17184 VSS.n2585 VSS.n2412 4.5005
R17185 VSS.n2587 VSS.n2412 4.5005
R17186 VSS.n2588 VSS.n2412 4.5005
R17187 VSS.n2590 VSS.n2412 4.5005
R17188 VSS.n2593 VSS.n2412 4.5005
R17189 VSS.n2595 VSS.n2412 4.5005
R17190 VSS.n2596 VSS.n2412 4.5005
R17191 VSS.n2598 VSS.n2412 4.5005
R17192 VSS.n2601 VSS.n2412 4.5005
R17193 VSS.n2603 VSS.n2412 4.5005
R17194 VSS.n2604 VSS.n2412 4.5005
R17195 VSS.n2606 VSS.n2412 4.5005
R17196 VSS.n2609 VSS.n2412 4.5005
R17197 VSS.n2611 VSS.n2412 4.5005
R17198 VSS.n2612 VSS.n2412 4.5005
R17199 VSS.n2614 VSS.n2412 4.5005
R17200 VSS.n2617 VSS.n2412 4.5005
R17201 VSS.n2619 VSS.n2412 4.5005
R17202 VSS.n2620 VSS.n2412 4.5005
R17203 VSS.n2622 VSS.n2412 4.5005
R17204 VSS.n2625 VSS.n2412 4.5005
R17205 VSS.n2627 VSS.n2412 4.5005
R17206 VSS.n2628 VSS.n2412 4.5005
R17207 VSS.n2630 VSS.n2412 4.5005
R17208 VSS.n2633 VSS.n2412 4.5005
R17209 VSS.n2635 VSS.n2412 4.5005
R17210 VSS.n2636 VSS.n2412 4.5005
R17211 VSS.n2638 VSS.n2412 4.5005
R17212 VSS.n2640 VSS.n2412 4.5005
R17213 VSS.n2642 VSS.n2412 4.5005
R17214 VSS.n2643 VSS.n2412 4.5005
R17215 VSS.n2645 VSS.n2412 4.5005
R17216 VSS.n2648 VSS.n2412 4.5005
R17217 VSS.n2650 VSS.n2412 4.5005
R17218 VSS.n2651 VSS.n2412 4.5005
R17219 VSS.n2653 VSS.n2412 4.5005
R17220 VSS.n2656 VSS.n2412 4.5005
R17221 VSS.n2658 VSS.n2412 4.5005
R17222 VSS.n2659 VSS.n2412 4.5005
R17223 VSS.n2661 VSS.n2412 4.5005
R17224 VSS.n2664 VSS.n2412 4.5005
R17225 VSS.n2666 VSS.n2412 4.5005
R17226 VSS.n2667 VSS.n2412 4.5005
R17227 VSS.n2669 VSS.n2412 4.5005
R17228 VSS.n2672 VSS.n2412 4.5005
R17229 VSS.n2674 VSS.n2412 4.5005
R17230 VSS.n2675 VSS.n2412 4.5005
R17231 VSS.n2677 VSS.n2412 4.5005
R17232 VSS.n2680 VSS.n2412 4.5005
R17233 VSS.n2682 VSS.n2412 4.5005
R17234 VSS.n2683 VSS.n2412 4.5005
R17235 VSS.n2685 VSS.n2412 4.5005
R17236 VSS.n2688 VSS.n2412 4.5005
R17237 VSS.n2690 VSS.n2412 4.5005
R17238 VSS.n2691 VSS.n2412 4.5005
R17239 VSS.n2693 VSS.n2412 4.5005
R17240 VSS.n2696 VSS.n2412 4.5005
R17241 VSS.n2698 VSS.n2412 4.5005
R17242 VSS.n2699 VSS.n2412 4.5005
R17243 VSS.n2701 VSS.n2412 4.5005
R17244 VSS.n2704 VSS.n2412 4.5005
R17245 VSS.n2706 VSS.n2412 4.5005
R17246 VSS.n2707 VSS.n2412 4.5005
R17247 VSS.n2709 VSS.n2412 4.5005
R17248 VSS.n2712 VSS.n2412 4.5005
R17249 VSS.n2714 VSS.n2412 4.5005
R17250 VSS.n2715 VSS.n2412 4.5005
R17251 VSS.n2717 VSS.n2412 4.5005
R17252 VSS.n2720 VSS.n2412 4.5005
R17253 VSS.n2722 VSS.n2412 4.5005
R17254 VSS.n2723 VSS.n2412 4.5005
R17255 VSS.n2725 VSS.n2412 4.5005
R17256 VSS.n2793 VSS.n2412 4.5005
R17257 VSS.n2859 VSS.n2412 4.5005
R17258 VSS.n3051 VSS.n2420 4.5005
R17259 VSS.n2420 VSS.n2351 4.5005
R17260 VSS.n2483 VSS.n2420 4.5005
R17261 VSS.n2484 VSS.n2420 4.5005
R17262 VSS.n2486 VSS.n2420 4.5005
R17263 VSS.n2489 VSS.n2420 4.5005
R17264 VSS.n2491 VSS.n2420 4.5005
R17265 VSS.n2492 VSS.n2420 4.5005
R17266 VSS.n2494 VSS.n2420 4.5005
R17267 VSS.n2497 VSS.n2420 4.5005
R17268 VSS.n2499 VSS.n2420 4.5005
R17269 VSS.n2500 VSS.n2420 4.5005
R17270 VSS.n2502 VSS.n2420 4.5005
R17271 VSS.n2505 VSS.n2420 4.5005
R17272 VSS.n2507 VSS.n2420 4.5005
R17273 VSS.n2508 VSS.n2420 4.5005
R17274 VSS.n2510 VSS.n2420 4.5005
R17275 VSS.n2513 VSS.n2420 4.5005
R17276 VSS.n2515 VSS.n2420 4.5005
R17277 VSS.n2516 VSS.n2420 4.5005
R17278 VSS.n2518 VSS.n2420 4.5005
R17279 VSS.n2521 VSS.n2420 4.5005
R17280 VSS.n2523 VSS.n2420 4.5005
R17281 VSS.n2524 VSS.n2420 4.5005
R17282 VSS.n2526 VSS.n2420 4.5005
R17283 VSS.n2529 VSS.n2420 4.5005
R17284 VSS.n2531 VSS.n2420 4.5005
R17285 VSS.n2532 VSS.n2420 4.5005
R17286 VSS.n2534 VSS.n2420 4.5005
R17287 VSS.n2537 VSS.n2420 4.5005
R17288 VSS.n2539 VSS.n2420 4.5005
R17289 VSS.n2540 VSS.n2420 4.5005
R17290 VSS.n2542 VSS.n2420 4.5005
R17291 VSS.n2545 VSS.n2420 4.5005
R17292 VSS.n2547 VSS.n2420 4.5005
R17293 VSS.n2548 VSS.n2420 4.5005
R17294 VSS.n2550 VSS.n2420 4.5005
R17295 VSS.n2553 VSS.n2420 4.5005
R17296 VSS.n2555 VSS.n2420 4.5005
R17297 VSS.n2556 VSS.n2420 4.5005
R17298 VSS.n2558 VSS.n2420 4.5005
R17299 VSS.n2561 VSS.n2420 4.5005
R17300 VSS.n2563 VSS.n2420 4.5005
R17301 VSS.n2564 VSS.n2420 4.5005
R17302 VSS.n2566 VSS.n2420 4.5005
R17303 VSS.n2569 VSS.n2420 4.5005
R17304 VSS.n2571 VSS.n2420 4.5005
R17305 VSS.n2572 VSS.n2420 4.5005
R17306 VSS.n2574 VSS.n2420 4.5005
R17307 VSS.n2577 VSS.n2420 4.5005
R17308 VSS.n2579 VSS.n2420 4.5005
R17309 VSS.n2580 VSS.n2420 4.5005
R17310 VSS.n2582 VSS.n2420 4.5005
R17311 VSS.n2585 VSS.n2420 4.5005
R17312 VSS.n2587 VSS.n2420 4.5005
R17313 VSS.n2588 VSS.n2420 4.5005
R17314 VSS.n2590 VSS.n2420 4.5005
R17315 VSS.n2593 VSS.n2420 4.5005
R17316 VSS.n2595 VSS.n2420 4.5005
R17317 VSS.n2596 VSS.n2420 4.5005
R17318 VSS.n2598 VSS.n2420 4.5005
R17319 VSS.n2601 VSS.n2420 4.5005
R17320 VSS.n2603 VSS.n2420 4.5005
R17321 VSS.n2604 VSS.n2420 4.5005
R17322 VSS.n2606 VSS.n2420 4.5005
R17323 VSS.n2609 VSS.n2420 4.5005
R17324 VSS.n2611 VSS.n2420 4.5005
R17325 VSS.n2612 VSS.n2420 4.5005
R17326 VSS.n2614 VSS.n2420 4.5005
R17327 VSS.n2617 VSS.n2420 4.5005
R17328 VSS.n2619 VSS.n2420 4.5005
R17329 VSS.n2620 VSS.n2420 4.5005
R17330 VSS.n2622 VSS.n2420 4.5005
R17331 VSS.n2625 VSS.n2420 4.5005
R17332 VSS.n2627 VSS.n2420 4.5005
R17333 VSS.n2628 VSS.n2420 4.5005
R17334 VSS.n2630 VSS.n2420 4.5005
R17335 VSS.n2633 VSS.n2420 4.5005
R17336 VSS.n2635 VSS.n2420 4.5005
R17337 VSS.n2636 VSS.n2420 4.5005
R17338 VSS.n2638 VSS.n2420 4.5005
R17339 VSS.n2640 VSS.n2420 4.5005
R17340 VSS.n2642 VSS.n2420 4.5005
R17341 VSS.n2643 VSS.n2420 4.5005
R17342 VSS.n2645 VSS.n2420 4.5005
R17343 VSS.n2648 VSS.n2420 4.5005
R17344 VSS.n2650 VSS.n2420 4.5005
R17345 VSS.n2651 VSS.n2420 4.5005
R17346 VSS.n2653 VSS.n2420 4.5005
R17347 VSS.n2656 VSS.n2420 4.5005
R17348 VSS.n2658 VSS.n2420 4.5005
R17349 VSS.n2659 VSS.n2420 4.5005
R17350 VSS.n2661 VSS.n2420 4.5005
R17351 VSS.n2664 VSS.n2420 4.5005
R17352 VSS.n2666 VSS.n2420 4.5005
R17353 VSS.n2667 VSS.n2420 4.5005
R17354 VSS.n2669 VSS.n2420 4.5005
R17355 VSS.n2672 VSS.n2420 4.5005
R17356 VSS.n2674 VSS.n2420 4.5005
R17357 VSS.n2675 VSS.n2420 4.5005
R17358 VSS.n2677 VSS.n2420 4.5005
R17359 VSS.n2680 VSS.n2420 4.5005
R17360 VSS.n2682 VSS.n2420 4.5005
R17361 VSS.n2683 VSS.n2420 4.5005
R17362 VSS.n2685 VSS.n2420 4.5005
R17363 VSS.n2688 VSS.n2420 4.5005
R17364 VSS.n2690 VSS.n2420 4.5005
R17365 VSS.n2691 VSS.n2420 4.5005
R17366 VSS.n2693 VSS.n2420 4.5005
R17367 VSS.n2696 VSS.n2420 4.5005
R17368 VSS.n2698 VSS.n2420 4.5005
R17369 VSS.n2699 VSS.n2420 4.5005
R17370 VSS.n2701 VSS.n2420 4.5005
R17371 VSS.n2704 VSS.n2420 4.5005
R17372 VSS.n2706 VSS.n2420 4.5005
R17373 VSS.n2707 VSS.n2420 4.5005
R17374 VSS.n2709 VSS.n2420 4.5005
R17375 VSS.n2712 VSS.n2420 4.5005
R17376 VSS.n2714 VSS.n2420 4.5005
R17377 VSS.n2715 VSS.n2420 4.5005
R17378 VSS.n2717 VSS.n2420 4.5005
R17379 VSS.n2720 VSS.n2420 4.5005
R17380 VSS.n2722 VSS.n2420 4.5005
R17381 VSS.n2723 VSS.n2420 4.5005
R17382 VSS.n2725 VSS.n2420 4.5005
R17383 VSS.n2793 VSS.n2420 4.5005
R17384 VSS.n2859 VSS.n2420 4.5005
R17385 VSS.n3051 VSS.n2411 4.5005
R17386 VSS.n2411 VSS.n2351 4.5005
R17387 VSS.n2483 VSS.n2411 4.5005
R17388 VSS.n2484 VSS.n2411 4.5005
R17389 VSS.n2486 VSS.n2411 4.5005
R17390 VSS.n2489 VSS.n2411 4.5005
R17391 VSS.n2491 VSS.n2411 4.5005
R17392 VSS.n2492 VSS.n2411 4.5005
R17393 VSS.n2494 VSS.n2411 4.5005
R17394 VSS.n2497 VSS.n2411 4.5005
R17395 VSS.n2499 VSS.n2411 4.5005
R17396 VSS.n2500 VSS.n2411 4.5005
R17397 VSS.n2502 VSS.n2411 4.5005
R17398 VSS.n2505 VSS.n2411 4.5005
R17399 VSS.n2507 VSS.n2411 4.5005
R17400 VSS.n2508 VSS.n2411 4.5005
R17401 VSS.n2510 VSS.n2411 4.5005
R17402 VSS.n2513 VSS.n2411 4.5005
R17403 VSS.n2515 VSS.n2411 4.5005
R17404 VSS.n2516 VSS.n2411 4.5005
R17405 VSS.n2518 VSS.n2411 4.5005
R17406 VSS.n2521 VSS.n2411 4.5005
R17407 VSS.n2523 VSS.n2411 4.5005
R17408 VSS.n2524 VSS.n2411 4.5005
R17409 VSS.n2526 VSS.n2411 4.5005
R17410 VSS.n2529 VSS.n2411 4.5005
R17411 VSS.n2531 VSS.n2411 4.5005
R17412 VSS.n2532 VSS.n2411 4.5005
R17413 VSS.n2534 VSS.n2411 4.5005
R17414 VSS.n2537 VSS.n2411 4.5005
R17415 VSS.n2539 VSS.n2411 4.5005
R17416 VSS.n2540 VSS.n2411 4.5005
R17417 VSS.n2542 VSS.n2411 4.5005
R17418 VSS.n2545 VSS.n2411 4.5005
R17419 VSS.n2547 VSS.n2411 4.5005
R17420 VSS.n2548 VSS.n2411 4.5005
R17421 VSS.n2550 VSS.n2411 4.5005
R17422 VSS.n2553 VSS.n2411 4.5005
R17423 VSS.n2555 VSS.n2411 4.5005
R17424 VSS.n2556 VSS.n2411 4.5005
R17425 VSS.n2558 VSS.n2411 4.5005
R17426 VSS.n2561 VSS.n2411 4.5005
R17427 VSS.n2563 VSS.n2411 4.5005
R17428 VSS.n2564 VSS.n2411 4.5005
R17429 VSS.n2566 VSS.n2411 4.5005
R17430 VSS.n2569 VSS.n2411 4.5005
R17431 VSS.n2571 VSS.n2411 4.5005
R17432 VSS.n2572 VSS.n2411 4.5005
R17433 VSS.n2574 VSS.n2411 4.5005
R17434 VSS.n2577 VSS.n2411 4.5005
R17435 VSS.n2579 VSS.n2411 4.5005
R17436 VSS.n2580 VSS.n2411 4.5005
R17437 VSS.n2582 VSS.n2411 4.5005
R17438 VSS.n2585 VSS.n2411 4.5005
R17439 VSS.n2587 VSS.n2411 4.5005
R17440 VSS.n2588 VSS.n2411 4.5005
R17441 VSS.n2590 VSS.n2411 4.5005
R17442 VSS.n2593 VSS.n2411 4.5005
R17443 VSS.n2595 VSS.n2411 4.5005
R17444 VSS.n2596 VSS.n2411 4.5005
R17445 VSS.n2598 VSS.n2411 4.5005
R17446 VSS.n2601 VSS.n2411 4.5005
R17447 VSS.n2603 VSS.n2411 4.5005
R17448 VSS.n2604 VSS.n2411 4.5005
R17449 VSS.n2606 VSS.n2411 4.5005
R17450 VSS.n2609 VSS.n2411 4.5005
R17451 VSS.n2611 VSS.n2411 4.5005
R17452 VSS.n2612 VSS.n2411 4.5005
R17453 VSS.n2614 VSS.n2411 4.5005
R17454 VSS.n2617 VSS.n2411 4.5005
R17455 VSS.n2619 VSS.n2411 4.5005
R17456 VSS.n2620 VSS.n2411 4.5005
R17457 VSS.n2622 VSS.n2411 4.5005
R17458 VSS.n2625 VSS.n2411 4.5005
R17459 VSS.n2627 VSS.n2411 4.5005
R17460 VSS.n2628 VSS.n2411 4.5005
R17461 VSS.n2630 VSS.n2411 4.5005
R17462 VSS.n2633 VSS.n2411 4.5005
R17463 VSS.n2635 VSS.n2411 4.5005
R17464 VSS.n2636 VSS.n2411 4.5005
R17465 VSS.n2638 VSS.n2411 4.5005
R17466 VSS.n2640 VSS.n2411 4.5005
R17467 VSS.n2642 VSS.n2411 4.5005
R17468 VSS.n2643 VSS.n2411 4.5005
R17469 VSS.n2645 VSS.n2411 4.5005
R17470 VSS.n2648 VSS.n2411 4.5005
R17471 VSS.n2650 VSS.n2411 4.5005
R17472 VSS.n2651 VSS.n2411 4.5005
R17473 VSS.n2653 VSS.n2411 4.5005
R17474 VSS.n2656 VSS.n2411 4.5005
R17475 VSS.n2658 VSS.n2411 4.5005
R17476 VSS.n2659 VSS.n2411 4.5005
R17477 VSS.n2661 VSS.n2411 4.5005
R17478 VSS.n2664 VSS.n2411 4.5005
R17479 VSS.n2666 VSS.n2411 4.5005
R17480 VSS.n2667 VSS.n2411 4.5005
R17481 VSS.n2669 VSS.n2411 4.5005
R17482 VSS.n2672 VSS.n2411 4.5005
R17483 VSS.n2674 VSS.n2411 4.5005
R17484 VSS.n2675 VSS.n2411 4.5005
R17485 VSS.n2677 VSS.n2411 4.5005
R17486 VSS.n2680 VSS.n2411 4.5005
R17487 VSS.n2682 VSS.n2411 4.5005
R17488 VSS.n2683 VSS.n2411 4.5005
R17489 VSS.n2685 VSS.n2411 4.5005
R17490 VSS.n2688 VSS.n2411 4.5005
R17491 VSS.n2690 VSS.n2411 4.5005
R17492 VSS.n2691 VSS.n2411 4.5005
R17493 VSS.n2693 VSS.n2411 4.5005
R17494 VSS.n2696 VSS.n2411 4.5005
R17495 VSS.n2698 VSS.n2411 4.5005
R17496 VSS.n2699 VSS.n2411 4.5005
R17497 VSS.n2701 VSS.n2411 4.5005
R17498 VSS.n2704 VSS.n2411 4.5005
R17499 VSS.n2706 VSS.n2411 4.5005
R17500 VSS.n2707 VSS.n2411 4.5005
R17501 VSS.n2709 VSS.n2411 4.5005
R17502 VSS.n2712 VSS.n2411 4.5005
R17503 VSS.n2714 VSS.n2411 4.5005
R17504 VSS.n2715 VSS.n2411 4.5005
R17505 VSS.n2717 VSS.n2411 4.5005
R17506 VSS.n2720 VSS.n2411 4.5005
R17507 VSS.n2722 VSS.n2411 4.5005
R17508 VSS.n2723 VSS.n2411 4.5005
R17509 VSS.n2725 VSS.n2411 4.5005
R17510 VSS.n2793 VSS.n2411 4.5005
R17511 VSS.n2859 VSS.n2411 4.5005
R17512 VSS.n3051 VSS.n2421 4.5005
R17513 VSS.n2421 VSS.n2351 4.5005
R17514 VSS.n2483 VSS.n2421 4.5005
R17515 VSS.n2484 VSS.n2421 4.5005
R17516 VSS.n2486 VSS.n2421 4.5005
R17517 VSS.n2489 VSS.n2421 4.5005
R17518 VSS.n2491 VSS.n2421 4.5005
R17519 VSS.n2492 VSS.n2421 4.5005
R17520 VSS.n2494 VSS.n2421 4.5005
R17521 VSS.n2497 VSS.n2421 4.5005
R17522 VSS.n2499 VSS.n2421 4.5005
R17523 VSS.n2500 VSS.n2421 4.5005
R17524 VSS.n2502 VSS.n2421 4.5005
R17525 VSS.n2505 VSS.n2421 4.5005
R17526 VSS.n2507 VSS.n2421 4.5005
R17527 VSS.n2508 VSS.n2421 4.5005
R17528 VSS.n2510 VSS.n2421 4.5005
R17529 VSS.n2513 VSS.n2421 4.5005
R17530 VSS.n2515 VSS.n2421 4.5005
R17531 VSS.n2516 VSS.n2421 4.5005
R17532 VSS.n2518 VSS.n2421 4.5005
R17533 VSS.n2521 VSS.n2421 4.5005
R17534 VSS.n2523 VSS.n2421 4.5005
R17535 VSS.n2524 VSS.n2421 4.5005
R17536 VSS.n2526 VSS.n2421 4.5005
R17537 VSS.n2529 VSS.n2421 4.5005
R17538 VSS.n2531 VSS.n2421 4.5005
R17539 VSS.n2532 VSS.n2421 4.5005
R17540 VSS.n2534 VSS.n2421 4.5005
R17541 VSS.n2537 VSS.n2421 4.5005
R17542 VSS.n2539 VSS.n2421 4.5005
R17543 VSS.n2540 VSS.n2421 4.5005
R17544 VSS.n2542 VSS.n2421 4.5005
R17545 VSS.n2545 VSS.n2421 4.5005
R17546 VSS.n2547 VSS.n2421 4.5005
R17547 VSS.n2548 VSS.n2421 4.5005
R17548 VSS.n2550 VSS.n2421 4.5005
R17549 VSS.n2553 VSS.n2421 4.5005
R17550 VSS.n2555 VSS.n2421 4.5005
R17551 VSS.n2556 VSS.n2421 4.5005
R17552 VSS.n2558 VSS.n2421 4.5005
R17553 VSS.n2561 VSS.n2421 4.5005
R17554 VSS.n2563 VSS.n2421 4.5005
R17555 VSS.n2564 VSS.n2421 4.5005
R17556 VSS.n2566 VSS.n2421 4.5005
R17557 VSS.n2569 VSS.n2421 4.5005
R17558 VSS.n2571 VSS.n2421 4.5005
R17559 VSS.n2572 VSS.n2421 4.5005
R17560 VSS.n2574 VSS.n2421 4.5005
R17561 VSS.n2577 VSS.n2421 4.5005
R17562 VSS.n2579 VSS.n2421 4.5005
R17563 VSS.n2580 VSS.n2421 4.5005
R17564 VSS.n2582 VSS.n2421 4.5005
R17565 VSS.n2585 VSS.n2421 4.5005
R17566 VSS.n2587 VSS.n2421 4.5005
R17567 VSS.n2588 VSS.n2421 4.5005
R17568 VSS.n2590 VSS.n2421 4.5005
R17569 VSS.n2593 VSS.n2421 4.5005
R17570 VSS.n2595 VSS.n2421 4.5005
R17571 VSS.n2596 VSS.n2421 4.5005
R17572 VSS.n2598 VSS.n2421 4.5005
R17573 VSS.n2601 VSS.n2421 4.5005
R17574 VSS.n2603 VSS.n2421 4.5005
R17575 VSS.n2604 VSS.n2421 4.5005
R17576 VSS.n2606 VSS.n2421 4.5005
R17577 VSS.n2609 VSS.n2421 4.5005
R17578 VSS.n2611 VSS.n2421 4.5005
R17579 VSS.n2612 VSS.n2421 4.5005
R17580 VSS.n2614 VSS.n2421 4.5005
R17581 VSS.n2617 VSS.n2421 4.5005
R17582 VSS.n2619 VSS.n2421 4.5005
R17583 VSS.n2620 VSS.n2421 4.5005
R17584 VSS.n2622 VSS.n2421 4.5005
R17585 VSS.n2625 VSS.n2421 4.5005
R17586 VSS.n2627 VSS.n2421 4.5005
R17587 VSS.n2628 VSS.n2421 4.5005
R17588 VSS.n2630 VSS.n2421 4.5005
R17589 VSS.n2633 VSS.n2421 4.5005
R17590 VSS.n2635 VSS.n2421 4.5005
R17591 VSS.n2636 VSS.n2421 4.5005
R17592 VSS.n2638 VSS.n2421 4.5005
R17593 VSS.n2640 VSS.n2421 4.5005
R17594 VSS.n2642 VSS.n2421 4.5005
R17595 VSS.n2643 VSS.n2421 4.5005
R17596 VSS.n2645 VSS.n2421 4.5005
R17597 VSS.n2648 VSS.n2421 4.5005
R17598 VSS.n2650 VSS.n2421 4.5005
R17599 VSS.n2651 VSS.n2421 4.5005
R17600 VSS.n2653 VSS.n2421 4.5005
R17601 VSS.n2656 VSS.n2421 4.5005
R17602 VSS.n2658 VSS.n2421 4.5005
R17603 VSS.n2659 VSS.n2421 4.5005
R17604 VSS.n2661 VSS.n2421 4.5005
R17605 VSS.n2664 VSS.n2421 4.5005
R17606 VSS.n2666 VSS.n2421 4.5005
R17607 VSS.n2667 VSS.n2421 4.5005
R17608 VSS.n2669 VSS.n2421 4.5005
R17609 VSS.n2672 VSS.n2421 4.5005
R17610 VSS.n2674 VSS.n2421 4.5005
R17611 VSS.n2675 VSS.n2421 4.5005
R17612 VSS.n2677 VSS.n2421 4.5005
R17613 VSS.n2680 VSS.n2421 4.5005
R17614 VSS.n2682 VSS.n2421 4.5005
R17615 VSS.n2683 VSS.n2421 4.5005
R17616 VSS.n2685 VSS.n2421 4.5005
R17617 VSS.n2688 VSS.n2421 4.5005
R17618 VSS.n2690 VSS.n2421 4.5005
R17619 VSS.n2691 VSS.n2421 4.5005
R17620 VSS.n2693 VSS.n2421 4.5005
R17621 VSS.n2696 VSS.n2421 4.5005
R17622 VSS.n2698 VSS.n2421 4.5005
R17623 VSS.n2699 VSS.n2421 4.5005
R17624 VSS.n2701 VSS.n2421 4.5005
R17625 VSS.n2704 VSS.n2421 4.5005
R17626 VSS.n2706 VSS.n2421 4.5005
R17627 VSS.n2707 VSS.n2421 4.5005
R17628 VSS.n2709 VSS.n2421 4.5005
R17629 VSS.n2712 VSS.n2421 4.5005
R17630 VSS.n2714 VSS.n2421 4.5005
R17631 VSS.n2715 VSS.n2421 4.5005
R17632 VSS.n2717 VSS.n2421 4.5005
R17633 VSS.n2720 VSS.n2421 4.5005
R17634 VSS.n2722 VSS.n2421 4.5005
R17635 VSS.n2723 VSS.n2421 4.5005
R17636 VSS.n2725 VSS.n2421 4.5005
R17637 VSS.n2793 VSS.n2421 4.5005
R17638 VSS.n2859 VSS.n2421 4.5005
R17639 VSS.n3051 VSS.n2410 4.5005
R17640 VSS.n2410 VSS.n2351 4.5005
R17641 VSS.n2483 VSS.n2410 4.5005
R17642 VSS.n2484 VSS.n2410 4.5005
R17643 VSS.n2486 VSS.n2410 4.5005
R17644 VSS.n2489 VSS.n2410 4.5005
R17645 VSS.n2491 VSS.n2410 4.5005
R17646 VSS.n2492 VSS.n2410 4.5005
R17647 VSS.n2494 VSS.n2410 4.5005
R17648 VSS.n2497 VSS.n2410 4.5005
R17649 VSS.n2499 VSS.n2410 4.5005
R17650 VSS.n2500 VSS.n2410 4.5005
R17651 VSS.n2502 VSS.n2410 4.5005
R17652 VSS.n2505 VSS.n2410 4.5005
R17653 VSS.n2507 VSS.n2410 4.5005
R17654 VSS.n2508 VSS.n2410 4.5005
R17655 VSS.n2510 VSS.n2410 4.5005
R17656 VSS.n2513 VSS.n2410 4.5005
R17657 VSS.n2515 VSS.n2410 4.5005
R17658 VSS.n2516 VSS.n2410 4.5005
R17659 VSS.n2518 VSS.n2410 4.5005
R17660 VSS.n2521 VSS.n2410 4.5005
R17661 VSS.n2523 VSS.n2410 4.5005
R17662 VSS.n2524 VSS.n2410 4.5005
R17663 VSS.n2526 VSS.n2410 4.5005
R17664 VSS.n2529 VSS.n2410 4.5005
R17665 VSS.n2531 VSS.n2410 4.5005
R17666 VSS.n2532 VSS.n2410 4.5005
R17667 VSS.n2534 VSS.n2410 4.5005
R17668 VSS.n2537 VSS.n2410 4.5005
R17669 VSS.n2539 VSS.n2410 4.5005
R17670 VSS.n2540 VSS.n2410 4.5005
R17671 VSS.n2542 VSS.n2410 4.5005
R17672 VSS.n2545 VSS.n2410 4.5005
R17673 VSS.n2547 VSS.n2410 4.5005
R17674 VSS.n2548 VSS.n2410 4.5005
R17675 VSS.n2550 VSS.n2410 4.5005
R17676 VSS.n2553 VSS.n2410 4.5005
R17677 VSS.n2555 VSS.n2410 4.5005
R17678 VSS.n2556 VSS.n2410 4.5005
R17679 VSS.n2558 VSS.n2410 4.5005
R17680 VSS.n2561 VSS.n2410 4.5005
R17681 VSS.n2563 VSS.n2410 4.5005
R17682 VSS.n2564 VSS.n2410 4.5005
R17683 VSS.n2566 VSS.n2410 4.5005
R17684 VSS.n2569 VSS.n2410 4.5005
R17685 VSS.n2571 VSS.n2410 4.5005
R17686 VSS.n2572 VSS.n2410 4.5005
R17687 VSS.n2574 VSS.n2410 4.5005
R17688 VSS.n2577 VSS.n2410 4.5005
R17689 VSS.n2579 VSS.n2410 4.5005
R17690 VSS.n2580 VSS.n2410 4.5005
R17691 VSS.n2582 VSS.n2410 4.5005
R17692 VSS.n2585 VSS.n2410 4.5005
R17693 VSS.n2587 VSS.n2410 4.5005
R17694 VSS.n2588 VSS.n2410 4.5005
R17695 VSS.n2590 VSS.n2410 4.5005
R17696 VSS.n2593 VSS.n2410 4.5005
R17697 VSS.n2595 VSS.n2410 4.5005
R17698 VSS.n2596 VSS.n2410 4.5005
R17699 VSS.n2598 VSS.n2410 4.5005
R17700 VSS.n2601 VSS.n2410 4.5005
R17701 VSS.n2603 VSS.n2410 4.5005
R17702 VSS.n2604 VSS.n2410 4.5005
R17703 VSS.n2606 VSS.n2410 4.5005
R17704 VSS.n2609 VSS.n2410 4.5005
R17705 VSS.n2611 VSS.n2410 4.5005
R17706 VSS.n2612 VSS.n2410 4.5005
R17707 VSS.n2614 VSS.n2410 4.5005
R17708 VSS.n2617 VSS.n2410 4.5005
R17709 VSS.n2619 VSS.n2410 4.5005
R17710 VSS.n2620 VSS.n2410 4.5005
R17711 VSS.n2622 VSS.n2410 4.5005
R17712 VSS.n2625 VSS.n2410 4.5005
R17713 VSS.n2627 VSS.n2410 4.5005
R17714 VSS.n2628 VSS.n2410 4.5005
R17715 VSS.n2630 VSS.n2410 4.5005
R17716 VSS.n2633 VSS.n2410 4.5005
R17717 VSS.n2635 VSS.n2410 4.5005
R17718 VSS.n2636 VSS.n2410 4.5005
R17719 VSS.n2638 VSS.n2410 4.5005
R17720 VSS.n2640 VSS.n2410 4.5005
R17721 VSS.n2642 VSS.n2410 4.5005
R17722 VSS.n2643 VSS.n2410 4.5005
R17723 VSS.n2645 VSS.n2410 4.5005
R17724 VSS.n2648 VSS.n2410 4.5005
R17725 VSS.n2650 VSS.n2410 4.5005
R17726 VSS.n2651 VSS.n2410 4.5005
R17727 VSS.n2653 VSS.n2410 4.5005
R17728 VSS.n2656 VSS.n2410 4.5005
R17729 VSS.n2658 VSS.n2410 4.5005
R17730 VSS.n2659 VSS.n2410 4.5005
R17731 VSS.n2661 VSS.n2410 4.5005
R17732 VSS.n2664 VSS.n2410 4.5005
R17733 VSS.n2666 VSS.n2410 4.5005
R17734 VSS.n2667 VSS.n2410 4.5005
R17735 VSS.n2669 VSS.n2410 4.5005
R17736 VSS.n2672 VSS.n2410 4.5005
R17737 VSS.n2674 VSS.n2410 4.5005
R17738 VSS.n2675 VSS.n2410 4.5005
R17739 VSS.n2677 VSS.n2410 4.5005
R17740 VSS.n2680 VSS.n2410 4.5005
R17741 VSS.n2682 VSS.n2410 4.5005
R17742 VSS.n2683 VSS.n2410 4.5005
R17743 VSS.n2685 VSS.n2410 4.5005
R17744 VSS.n2688 VSS.n2410 4.5005
R17745 VSS.n2690 VSS.n2410 4.5005
R17746 VSS.n2691 VSS.n2410 4.5005
R17747 VSS.n2693 VSS.n2410 4.5005
R17748 VSS.n2696 VSS.n2410 4.5005
R17749 VSS.n2698 VSS.n2410 4.5005
R17750 VSS.n2699 VSS.n2410 4.5005
R17751 VSS.n2701 VSS.n2410 4.5005
R17752 VSS.n2704 VSS.n2410 4.5005
R17753 VSS.n2706 VSS.n2410 4.5005
R17754 VSS.n2707 VSS.n2410 4.5005
R17755 VSS.n2709 VSS.n2410 4.5005
R17756 VSS.n2712 VSS.n2410 4.5005
R17757 VSS.n2714 VSS.n2410 4.5005
R17758 VSS.n2715 VSS.n2410 4.5005
R17759 VSS.n2717 VSS.n2410 4.5005
R17760 VSS.n2720 VSS.n2410 4.5005
R17761 VSS.n2722 VSS.n2410 4.5005
R17762 VSS.n2723 VSS.n2410 4.5005
R17763 VSS.n2725 VSS.n2410 4.5005
R17764 VSS.n2793 VSS.n2410 4.5005
R17765 VSS.n2859 VSS.n2410 4.5005
R17766 VSS.n3051 VSS.n2422 4.5005
R17767 VSS.n2422 VSS.n2351 4.5005
R17768 VSS.n2483 VSS.n2422 4.5005
R17769 VSS.n2484 VSS.n2422 4.5005
R17770 VSS.n2486 VSS.n2422 4.5005
R17771 VSS.n2489 VSS.n2422 4.5005
R17772 VSS.n2491 VSS.n2422 4.5005
R17773 VSS.n2492 VSS.n2422 4.5005
R17774 VSS.n2494 VSS.n2422 4.5005
R17775 VSS.n2497 VSS.n2422 4.5005
R17776 VSS.n2499 VSS.n2422 4.5005
R17777 VSS.n2500 VSS.n2422 4.5005
R17778 VSS.n2502 VSS.n2422 4.5005
R17779 VSS.n2505 VSS.n2422 4.5005
R17780 VSS.n2507 VSS.n2422 4.5005
R17781 VSS.n2508 VSS.n2422 4.5005
R17782 VSS.n2510 VSS.n2422 4.5005
R17783 VSS.n2513 VSS.n2422 4.5005
R17784 VSS.n2515 VSS.n2422 4.5005
R17785 VSS.n2516 VSS.n2422 4.5005
R17786 VSS.n2518 VSS.n2422 4.5005
R17787 VSS.n2521 VSS.n2422 4.5005
R17788 VSS.n2523 VSS.n2422 4.5005
R17789 VSS.n2524 VSS.n2422 4.5005
R17790 VSS.n2526 VSS.n2422 4.5005
R17791 VSS.n2529 VSS.n2422 4.5005
R17792 VSS.n2531 VSS.n2422 4.5005
R17793 VSS.n2532 VSS.n2422 4.5005
R17794 VSS.n2534 VSS.n2422 4.5005
R17795 VSS.n2537 VSS.n2422 4.5005
R17796 VSS.n2539 VSS.n2422 4.5005
R17797 VSS.n2540 VSS.n2422 4.5005
R17798 VSS.n2542 VSS.n2422 4.5005
R17799 VSS.n2545 VSS.n2422 4.5005
R17800 VSS.n2547 VSS.n2422 4.5005
R17801 VSS.n2548 VSS.n2422 4.5005
R17802 VSS.n2550 VSS.n2422 4.5005
R17803 VSS.n2553 VSS.n2422 4.5005
R17804 VSS.n2555 VSS.n2422 4.5005
R17805 VSS.n2556 VSS.n2422 4.5005
R17806 VSS.n2558 VSS.n2422 4.5005
R17807 VSS.n2561 VSS.n2422 4.5005
R17808 VSS.n2563 VSS.n2422 4.5005
R17809 VSS.n2564 VSS.n2422 4.5005
R17810 VSS.n2566 VSS.n2422 4.5005
R17811 VSS.n2569 VSS.n2422 4.5005
R17812 VSS.n2571 VSS.n2422 4.5005
R17813 VSS.n2572 VSS.n2422 4.5005
R17814 VSS.n2574 VSS.n2422 4.5005
R17815 VSS.n2577 VSS.n2422 4.5005
R17816 VSS.n2579 VSS.n2422 4.5005
R17817 VSS.n2580 VSS.n2422 4.5005
R17818 VSS.n2582 VSS.n2422 4.5005
R17819 VSS.n2585 VSS.n2422 4.5005
R17820 VSS.n2587 VSS.n2422 4.5005
R17821 VSS.n2588 VSS.n2422 4.5005
R17822 VSS.n2590 VSS.n2422 4.5005
R17823 VSS.n2593 VSS.n2422 4.5005
R17824 VSS.n2595 VSS.n2422 4.5005
R17825 VSS.n2596 VSS.n2422 4.5005
R17826 VSS.n2598 VSS.n2422 4.5005
R17827 VSS.n2601 VSS.n2422 4.5005
R17828 VSS.n2603 VSS.n2422 4.5005
R17829 VSS.n2604 VSS.n2422 4.5005
R17830 VSS.n2606 VSS.n2422 4.5005
R17831 VSS.n2609 VSS.n2422 4.5005
R17832 VSS.n2611 VSS.n2422 4.5005
R17833 VSS.n2612 VSS.n2422 4.5005
R17834 VSS.n2614 VSS.n2422 4.5005
R17835 VSS.n2617 VSS.n2422 4.5005
R17836 VSS.n2619 VSS.n2422 4.5005
R17837 VSS.n2620 VSS.n2422 4.5005
R17838 VSS.n2622 VSS.n2422 4.5005
R17839 VSS.n2625 VSS.n2422 4.5005
R17840 VSS.n2627 VSS.n2422 4.5005
R17841 VSS.n2628 VSS.n2422 4.5005
R17842 VSS.n2630 VSS.n2422 4.5005
R17843 VSS.n2633 VSS.n2422 4.5005
R17844 VSS.n2635 VSS.n2422 4.5005
R17845 VSS.n2636 VSS.n2422 4.5005
R17846 VSS.n2638 VSS.n2422 4.5005
R17847 VSS.n2640 VSS.n2422 4.5005
R17848 VSS.n2642 VSS.n2422 4.5005
R17849 VSS.n2643 VSS.n2422 4.5005
R17850 VSS.n2645 VSS.n2422 4.5005
R17851 VSS.n2648 VSS.n2422 4.5005
R17852 VSS.n2650 VSS.n2422 4.5005
R17853 VSS.n2651 VSS.n2422 4.5005
R17854 VSS.n2653 VSS.n2422 4.5005
R17855 VSS.n2656 VSS.n2422 4.5005
R17856 VSS.n2658 VSS.n2422 4.5005
R17857 VSS.n2659 VSS.n2422 4.5005
R17858 VSS.n2661 VSS.n2422 4.5005
R17859 VSS.n2664 VSS.n2422 4.5005
R17860 VSS.n2666 VSS.n2422 4.5005
R17861 VSS.n2667 VSS.n2422 4.5005
R17862 VSS.n2669 VSS.n2422 4.5005
R17863 VSS.n2672 VSS.n2422 4.5005
R17864 VSS.n2674 VSS.n2422 4.5005
R17865 VSS.n2675 VSS.n2422 4.5005
R17866 VSS.n2677 VSS.n2422 4.5005
R17867 VSS.n2680 VSS.n2422 4.5005
R17868 VSS.n2682 VSS.n2422 4.5005
R17869 VSS.n2683 VSS.n2422 4.5005
R17870 VSS.n2685 VSS.n2422 4.5005
R17871 VSS.n2688 VSS.n2422 4.5005
R17872 VSS.n2690 VSS.n2422 4.5005
R17873 VSS.n2691 VSS.n2422 4.5005
R17874 VSS.n2693 VSS.n2422 4.5005
R17875 VSS.n2696 VSS.n2422 4.5005
R17876 VSS.n2698 VSS.n2422 4.5005
R17877 VSS.n2699 VSS.n2422 4.5005
R17878 VSS.n2701 VSS.n2422 4.5005
R17879 VSS.n2704 VSS.n2422 4.5005
R17880 VSS.n2706 VSS.n2422 4.5005
R17881 VSS.n2707 VSS.n2422 4.5005
R17882 VSS.n2709 VSS.n2422 4.5005
R17883 VSS.n2712 VSS.n2422 4.5005
R17884 VSS.n2714 VSS.n2422 4.5005
R17885 VSS.n2715 VSS.n2422 4.5005
R17886 VSS.n2717 VSS.n2422 4.5005
R17887 VSS.n2720 VSS.n2422 4.5005
R17888 VSS.n2722 VSS.n2422 4.5005
R17889 VSS.n2723 VSS.n2422 4.5005
R17890 VSS.n2725 VSS.n2422 4.5005
R17891 VSS.n2793 VSS.n2422 4.5005
R17892 VSS.n2859 VSS.n2422 4.5005
R17893 VSS.n3051 VSS.n2409 4.5005
R17894 VSS.n2409 VSS.n2351 4.5005
R17895 VSS.n2483 VSS.n2409 4.5005
R17896 VSS.n2484 VSS.n2409 4.5005
R17897 VSS.n2486 VSS.n2409 4.5005
R17898 VSS.n2489 VSS.n2409 4.5005
R17899 VSS.n2491 VSS.n2409 4.5005
R17900 VSS.n2492 VSS.n2409 4.5005
R17901 VSS.n2494 VSS.n2409 4.5005
R17902 VSS.n2497 VSS.n2409 4.5005
R17903 VSS.n2499 VSS.n2409 4.5005
R17904 VSS.n2500 VSS.n2409 4.5005
R17905 VSS.n2502 VSS.n2409 4.5005
R17906 VSS.n2505 VSS.n2409 4.5005
R17907 VSS.n2507 VSS.n2409 4.5005
R17908 VSS.n2508 VSS.n2409 4.5005
R17909 VSS.n2510 VSS.n2409 4.5005
R17910 VSS.n2513 VSS.n2409 4.5005
R17911 VSS.n2515 VSS.n2409 4.5005
R17912 VSS.n2516 VSS.n2409 4.5005
R17913 VSS.n2518 VSS.n2409 4.5005
R17914 VSS.n2521 VSS.n2409 4.5005
R17915 VSS.n2523 VSS.n2409 4.5005
R17916 VSS.n2524 VSS.n2409 4.5005
R17917 VSS.n2526 VSS.n2409 4.5005
R17918 VSS.n2529 VSS.n2409 4.5005
R17919 VSS.n2531 VSS.n2409 4.5005
R17920 VSS.n2532 VSS.n2409 4.5005
R17921 VSS.n2534 VSS.n2409 4.5005
R17922 VSS.n2537 VSS.n2409 4.5005
R17923 VSS.n2539 VSS.n2409 4.5005
R17924 VSS.n2540 VSS.n2409 4.5005
R17925 VSS.n2542 VSS.n2409 4.5005
R17926 VSS.n2545 VSS.n2409 4.5005
R17927 VSS.n2547 VSS.n2409 4.5005
R17928 VSS.n2548 VSS.n2409 4.5005
R17929 VSS.n2550 VSS.n2409 4.5005
R17930 VSS.n2553 VSS.n2409 4.5005
R17931 VSS.n2555 VSS.n2409 4.5005
R17932 VSS.n2556 VSS.n2409 4.5005
R17933 VSS.n2558 VSS.n2409 4.5005
R17934 VSS.n2561 VSS.n2409 4.5005
R17935 VSS.n2563 VSS.n2409 4.5005
R17936 VSS.n2564 VSS.n2409 4.5005
R17937 VSS.n2566 VSS.n2409 4.5005
R17938 VSS.n2569 VSS.n2409 4.5005
R17939 VSS.n2571 VSS.n2409 4.5005
R17940 VSS.n2572 VSS.n2409 4.5005
R17941 VSS.n2574 VSS.n2409 4.5005
R17942 VSS.n2577 VSS.n2409 4.5005
R17943 VSS.n2579 VSS.n2409 4.5005
R17944 VSS.n2580 VSS.n2409 4.5005
R17945 VSS.n2582 VSS.n2409 4.5005
R17946 VSS.n2585 VSS.n2409 4.5005
R17947 VSS.n2587 VSS.n2409 4.5005
R17948 VSS.n2588 VSS.n2409 4.5005
R17949 VSS.n2590 VSS.n2409 4.5005
R17950 VSS.n2593 VSS.n2409 4.5005
R17951 VSS.n2595 VSS.n2409 4.5005
R17952 VSS.n2596 VSS.n2409 4.5005
R17953 VSS.n2598 VSS.n2409 4.5005
R17954 VSS.n2601 VSS.n2409 4.5005
R17955 VSS.n2603 VSS.n2409 4.5005
R17956 VSS.n2604 VSS.n2409 4.5005
R17957 VSS.n2606 VSS.n2409 4.5005
R17958 VSS.n2609 VSS.n2409 4.5005
R17959 VSS.n2611 VSS.n2409 4.5005
R17960 VSS.n2612 VSS.n2409 4.5005
R17961 VSS.n2614 VSS.n2409 4.5005
R17962 VSS.n2617 VSS.n2409 4.5005
R17963 VSS.n2619 VSS.n2409 4.5005
R17964 VSS.n2620 VSS.n2409 4.5005
R17965 VSS.n2622 VSS.n2409 4.5005
R17966 VSS.n2625 VSS.n2409 4.5005
R17967 VSS.n2627 VSS.n2409 4.5005
R17968 VSS.n2628 VSS.n2409 4.5005
R17969 VSS.n2630 VSS.n2409 4.5005
R17970 VSS.n2633 VSS.n2409 4.5005
R17971 VSS.n2635 VSS.n2409 4.5005
R17972 VSS.n2636 VSS.n2409 4.5005
R17973 VSS.n2638 VSS.n2409 4.5005
R17974 VSS.n2640 VSS.n2409 4.5005
R17975 VSS.n2642 VSS.n2409 4.5005
R17976 VSS.n2643 VSS.n2409 4.5005
R17977 VSS.n2645 VSS.n2409 4.5005
R17978 VSS.n2648 VSS.n2409 4.5005
R17979 VSS.n2650 VSS.n2409 4.5005
R17980 VSS.n2651 VSS.n2409 4.5005
R17981 VSS.n2653 VSS.n2409 4.5005
R17982 VSS.n2656 VSS.n2409 4.5005
R17983 VSS.n2658 VSS.n2409 4.5005
R17984 VSS.n2659 VSS.n2409 4.5005
R17985 VSS.n2661 VSS.n2409 4.5005
R17986 VSS.n2664 VSS.n2409 4.5005
R17987 VSS.n2666 VSS.n2409 4.5005
R17988 VSS.n2667 VSS.n2409 4.5005
R17989 VSS.n2669 VSS.n2409 4.5005
R17990 VSS.n2672 VSS.n2409 4.5005
R17991 VSS.n2674 VSS.n2409 4.5005
R17992 VSS.n2675 VSS.n2409 4.5005
R17993 VSS.n2677 VSS.n2409 4.5005
R17994 VSS.n2680 VSS.n2409 4.5005
R17995 VSS.n2682 VSS.n2409 4.5005
R17996 VSS.n2683 VSS.n2409 4.5005
R17997 VSS.n2685 VSS.n2409 4.5005
R17998 VSS.n2688 VSS.n2409 4.5005
R17999 VSS.n2690 VSS.n2409 4.5005
R18000 VSS.n2691 VSS.n2409 4.5005
R18001 VSS.n2693 VSS.n2409 4.5005
R18002 VSS.n2696 VSS.n2409 4.5005
R18003 VSS.n2698 VSS.n2409 4.5005
R18004 VSS.n2699 VSS.n2409 4.5005
R18005 VSS.n2701 VSS.n2409 4.5005
R18006 VSS.n2704 VSS.n2409 4.5005
R18007 VSS.n2706 VSS.n2409 4.5005
R18008 VSS.n2707 VSS.n2409 4.5005
R18009 VSS.n2709 VSS.n2409 4.5005
R18010 VSS.n2712 VSS.n2409 4.5005
R18011 VSS.n2714 VSS.n2409 4.5005
R18012 VSS.n2715 VSS.n2409 4.5005
R18013 VSS.n2717 VSS.n2409 4.5005
R18014 VSS.n2720 VSS.n2409 4.5005
R18015 VSS.n2722 VSS.n2409 4.5005
R18016 VSS.n2723 VSS.n2409 4.5005
R18017 VSS.n2725 VSS.n2409 4.5005
R18018 VSS.n2793 VSS.n2409 4.5005
R18019 VSS.n2859 VSS.n2409 4.5005
R18020 VSS.n3051 VSS.n2423 4.5005
R18021 VSS.n2423 VSS.n2351 4.5005
R18022 VSS.n2483 VSS.n2423 4.5005
R18023 VSS.n2484 VSS.n2423 4.5005
R18024 VSS.n2486 VSS.n2423 4.5005
R18025 VSS.n2489 VSS.n2423 4.5005
R18026 VSS.n2491 VSS.n2423 4.5005
R18027 VSS.n2492 VSS.n2423 4.5005
R18028 VSS.n2494 VSS.n2423 4.5005
R18029 VSS.n2497 VSS.n2423 4.5005
R18030 VSS.n2499 VSS.n2423 4.5005
R18031 VSS.n2500 VSS.n2423 4.5005
R18032 VSS.n2502 VSS.n2423 4.5005
R18033 VSS.n2505 VSS.n2423 4.5005
R18034 VSS.n2507 VSS.n2423 4.5005
R18035 VSS.n2508 VSS.n2423 4.5005
R18036 VSS.n2510 VSS.n2423 4.5005
R18037 VSS.n2513 VSS.n2423 4.5005
R18038 VSS.n2515 VSS.n2423 4.5005
R18039 VSS.n2516 VSS.n2423 4.5005
R18040 VSS.n2518 VSS.n2423 4.5005
R18041 VSS.n2521 VSS.n2423 4.5005
R18042 VSS.n2523 VSS.n2423 4.5005
R18043 VSS.n2524 VSS.n2423 4.5005
R18044 VSS.n2526 VSS.n2423 4.5005
R18045 VSS.n2529 VSS.n2423 4.5005
R18046 VSS.n2531 VSS.n2423 4.5005
R18047 VSS.n2532 VSS.n2423 4.5005
R18048 VSS.n2534 VSS.n2423 4.5005
R18049 VSS.n2537 VSS.n2423 4.5005
R18050 VSS.n2539 VSS.n2423 4.5005
R18051 VSS.n2540 VSS.n2423 4.5005
R18052 VSS.n2542 VSS.n2423 4.5005
R18053 VSS.n2545 VSS.n2423 4.5005
R18054 VSS.n2547 VSS.n2423 4.5005
R18055 VSS.n2548 VSS.n2423 4.5005
R18056 VSS.n2550 VSS.n2423 4.5005
R18057 VSS.n2553 VSS.n2423 4.5005
R18058 VSS.n2555 VSS.n2423 4.5005
R18059 VSS.n2556 VSS.n2423 4.5005
R18060 VSS.n2558 VSS.n2423 4.5005
R18061 VSS.n2561 VSS.n2423 4.5005
R18062 VSS.n2563 VSS.n2423 4.5005
R18063 VSS.n2564 VSS.n2423 4.5005
R18064 VSS.n2566 VSS.n2423 4.5005
R18065 VSS.n2569 VSS.n2423 4.5005
R18066 VSS.n2571 VSS.n2423 4.5005
R18067 VSS.n2572 VSS.n2423 4.5005
R18068 VSS.n2574 VSS.n2423 4.5005
R18069 VSS.n2577 VSS.n2423 4.5005
R18070 VSS.n2579 VSS.n2423 4.5005
R18071 VSS.n2580 VSS.n2423 4.5005
R18072 VSS.n2582 VSS.n2423 4.5005
R18073 VSS.n2585 VSS.n2423 4.5005
R18074 VSS.n2587 VSS.n2423 4.5005
R18075 VSS.n2588 VSS.n2423 4.5005
R18076 VSS.n2590 VSS.n2423 4.5005
R18077 VSS.n2593 VSS.n2423 4.5005
R18078 VSS.n2595 VSS.n2423 4.5005
R18079 VSS.n2596 VSS.n2423 4.5005
R18080 VSS.n2598 VSS.n2423 4.5005
R18081 VSS.n2601 VSS.n2423 4.5005
R18082 VSS.n2603 VSS.n2423 4.5005
R18083 VSS.n2604 VSS.n2423 4.5005
R18084 VSS.n2606 VSS.n2423 4.5005
R18085 VSS.n2609 VSS.n2423 4.5005
R18086 VSS.n2611 VSS.n2423 4.5005
R18087 VSS.n2612 VSS.n2423 4.5005
R18088 VSS.n2614 VSS.n2423 4.5005
R18089 VSS.n2617 VSS.n2423 4.5005
R18090 VSS.n2619 VSS.n2423 4.5005
R18091 VSS.n2620 VSS.n2423 4.5005
R18092 VSS.n2622 VSS.n2423 4.5005
R18093 VSS.n2625 VSS.n2423 4.5005
R18094 VSS.n2627 VSS.n2423 4.5005
R18095 VSS.n2628 VSS.n2423 4.5005
R18096 VSS.n2630 VSS.n2423 4.5005
R18097 VSS.n2633 VSS.n2423 4.5005
R18098 VSS.n2635 VSS.n2423 4.5005
R18099 VSS.n2636 VSS.n2423 4.5005
R18100 VSS.n2638 VSS.n2423 4.5005
R18101 VSS.n2640 VSS.n2423 4.5005
R18102 VSS.n2642 VSS.n2423 4.5005
R18103 VSS.n2643 VSS.n2423 4.5005
R18104 VSS.n2645 VSS.n2423 4.5005
R18105 VSS.n2648 VSS.n2423 4.5005
R18106 VSS.n2650 VSS.n2423 4.5005
R18107 VSS.n2651 VSS.n2423 4.5005
R18108 VSS.n2653 VSS.n2423 4.5005
R18109 VSS.n2656 VSS.n2423 4.5005
R18110 VSS.n2658 VSS.n2423 4.5005
R18111 VSS.n2659 VSS.n2423 4.5005
R18112 VSS.n2661 VSS.n2423 4.5005
R18113 VSS.n2664 VSS.n2423 4.5005
R18114 VSS.n2666 VSS.n2423 4.5005
R18115 VSS.n2667 VSS.n2423 4.5005
R18116 VSS.n2669 VSS.n2423 4.5005
R18117 VSS.n2672 VSS.n2423 4.5005
R18118 VSS.n2674 VSS.n2423 4.5005
R18119 VSS.n2675 VSS.n2423 4.5005
R18120 VSS.n2677 VSS.n2423 4.5005
R18121 VSS.n2680 VSS.n2423 4.5005
R18122 VSS.n2682 VSS.n2423 4.5005
R18123 VSS.n2683 VSS.n2423 4.5005
R18124 VSS.n2685 VSS.n2423 4.5005
R18125 VSS.n2688 VSS.n2423 4.5005
R18126 VSS.n2690 VSS.n2423 4.5005
R18127 VSS.n2691 VSS.n2423 4.5005
R18128 VSS.n2693 VSS.n2423 4.5005
R18129 VSS.n2696 VSS.n2423 4.5005
R18130 VSS.n2698 VSS.n2423 4.5005
R18131 VSS.n2699 VSS.n2423 4.5005
R18132 VSS.n2701 VSS.n2423 4.5005
R18133 VSS.n2704 VSS.n2423 4.5005
R18134 VSS.n2706 VSS.n2423 4.5005
R18135 VSS.n2707 VSS.n2423 4.5005
R18136 VSS.n2709 VSS.n2423 4.5005
R18137 VSS.n2712 VSS.n2423 4.5005
R18138 VSS.n2714 VSS.n2423 4.5005
R18139 VSS.n2715 VSS.n2423 4.5005
R18140 VSS.n2717 VSS.n2423 4.5005
R18141 VSS.n2720 VSS.n2423 4.5005
R18142 VSS.n2722 VSS.n2423 4.5005
R18143 VSS.n2723 VSS.n2423 4.5005
R18144 VSS.n2725 VSS.n2423 4.5005
R18145 VSS.n2793 VSS.n2423 4.5005
R18146 VSS.n2859 VSS.n2423 4.5005
R18147 VSS.n3051 VSS.n2408 4.5005
R18148 VSS.n2408 VSS.n2351 4.5005
R18149 VSS.n2483 VSS.n2408 4.5005
R18150 VSS.n2484 VSS.n2408 4.5005
R18151 VSS.n2486 VSS.n2408 4.5005
R18152 VSS.n2489 VSS.n2408 4.5005
R18153 VSS.n2491 VSS.n2408 4.5005
R18154 VSS.n2492 VSS.n2408 4.5005
R18155 VSS.n2494 VSS.n2408 4.5005
R18156 VSS.n2497 VSS.n2408 4.5005
R18157 VSS.n2499 VSS.n2408 4.5005
R18158 VSS.n2500 VSS.n2408 4.5005
R18159 VSS.n2502 VSS.n2408 4.5005
R18160 VSS.n2505 VSS.n2408 4.5005
R18161 VSS.n2507 VSS.n2408 4.5005
R18162 VSS.n2508 VSS.n2408 4.5005
R18163 VSS.n2510 VSS.n2408 4.5005
R18164 VSS.n2513 VSS.n2408 4.5005
R18165 VSS.n2515 VSS.n2408 4.5005
R18166 VSS.n2516 VSS.n2408 4.5005
R18167 VSS.n2518 VSS.n2408 4.5005
R18168 VSS.n2521 VSS.n2408 4.5005
R18169 VSS.n2523 VSS.n2408 4.5005
R18170 VSS.n2524 VSS.n2408 4.5005
R18171 VSS.n2526 VSS.n2408 4.5005
R18172 VSS.n2529 VSS.n2408 4.5005
R18173 VSS.n2531 VSS.n2408 4.5005
R18174 VSS.n2532 VSS.n2408 4.5005
R18175 VSS.n2534 VSS.n2408 4.5005
R18176 VSS.n2537 VSS.n2408 4.5005
R18177 VSS.n2539 VSS.n2408 4.5005
R18178 VSS.n2540 VSS.n2408 4.5005
R18179 VSS.n2542 VSS.n2408 4.5005
R18180 VSS.n2545 VSS.n2408 4.5005
R18181 VSS.n2547 VSS.n2408 4.5005
R18182 VSS.n2548 VSS.n2408 4.5005
R18183 VSS.n2550 VSS.n2408 4.5005
R18184 VSS.n2553 VSS.n2408 4.5005
R18185 VSS.n2555 VSS.n2408 4.5005
R18186 VSS.n2556 VSS.n2408 4.5005
R18187 VSS.n2558 VSS.n2408 4.5005
R18188 VSS.n2561 VSS.n2408 4.5005
R18189 VSS.n2563 VSS.n2408 4.5005
R18190 VSS.n2564 VSS.n2408 4.5005
R18191 VSS.n2566 VSS.n2408 4.5005
R18192 VSS.n2569 VSS.n2408 4.5005
R18193 VSS.n2571 VSS.n2408 4.5005
R18194 VSS.n2572 VSS.n2408 4.5005
R18195 VSS.n2574 VSS.n2408 4.5005
R18196 VSS.n2577 VSS.n2408 4.5005
R18197 VSS.n2579 VSS.n2408 4.5005
R18198 VSS.n2580 VSS.n2408 4.5005
R18199 VSS.n2582 VSS.n2408 4.5005
R18200 VSS.n2585 VSS.n2408 4.5005
R18201 VSS.n2587 VSS.n2408 4.5005
R18202 VSS.n2588 VSS.n2408 4.5005
R18203 VSS.n2590 VSS.n2408 4.5005
R18204 VSS.n2593 VSS.n2408 4.5005
R18205 VSS.n2595 VSS.n2408 4.5005
R18206 VSS.n2596 VSS.n2408 4.5005
R18207 VSS.n2598 VSS.n2408 4.5005
R18208 VSS.n2601 VSS.n2408 4.5005
R18209 VSS.n2603 VSS.n2408 4.5005
R18210 VSS.n2604 VSS.n2408 4.5005
R18211 VSS.n2606 VSS.n2408 4.5005
R18212 VSS.n2609 VSS.n2408 4.5005
R18213 VSS.n2611 VSS.n2408 4.5005
R18214 VSS.n2612 VSS.n2408 4.5005
R18215 VSS.n2614 VSS.n2408 4.5005
R18216 VSS.n2617 VSS.n2408 4.5005
R18217 VSS.n2619 VSS.n2408 4.5005
R18218 VSS.n2620 VSS.n2408 4.5005
R18219 VSS.n2622 VSS.n2408 4.5005
R18220 VSS.n2625 VSS.n2408 4.5005
R18221 VSS.n2627 VSS.n2408 4.5005
R18222 VSS.n2628 VSS.n2408 4.5005
R18223 VSS.n2630 VSS.n2408 4.5005
R18224 VSS.n2633 VSS.n2408 4.5005
R18225 VSS.n2635 VSS.n2408 4.5005
R18226 VSS.n2636 VSS.n2408 4.5005
R18227 VSS.n2638 VSS.n2408 4.5005
R18228 VSS.n2640 VSS.n2408 4.5005
R18229 VSS.n2642 VSS.n2408 4.5005
R18230 VSS.n2643 VSS.n2408 4.5005
R18231 VSS.n2645 VSS.n2408 4.5005
R18232 VSS.n2648 VSS.n2408 4.5005
R18233 VSS.n2650 VSS.n2408 4.5005
R18234 VSS.n2651 VSS.n2408 4.5005
R18235 VSS.n2653 VSS.n2408 4.5005
R18236 VSS.n2656 VSS.n2408 4.5005
R18237 VSS.n2658 VSS.n2408 4.5005
R18238 VSS.n2659 VSS.n2408 4.5005
R18239 VSS.n2661 VSS.n2408 4.5005
R18240 VSS.n2664 VSS.n2408 4.5005
R18241 VSS.n2666 VSS.n2408 4.5005
R18242 VSS.n2667 VSS.n2408 4.5005
R18243 VSS.n2669 VSS.n2408 4.5005
R18244 VSS.n2672 VSS.n2408 4.5005
R18245 VSS.n2674 VSS.n2408 4.5005
R18246 VSS.n2675 VSS.n2408 4.5005
R18247 VSS.n2677 VSS.n2408 4.5005
R18248 VSS.n2680 VSS.n2408 4.5005
R18249 VSS.n2682 VSS.n2408 4.5005
R18250 VSS.n2683 VSS.n2408 4.5005
R18251 VSS.n2685 VSS.n2408 4.5005
R18252 VSS.n2688 VSS.n2408 4.5005
R18253 VSS.n2690 VSS.n2408 4.5005
R18254 VSS.n2691 VSS.n2408 4.5005
R18255 VSS.n2693 VSS.n2408 4.5005
R18256 VSS.n2696 VSS.n2408 4.5005
R18257 VSS.n2698 VSS.n2408 4.5005
R18258 VSS.n2699 VSS.n2408 4.5005
R18259 VSS.n2701 VSS.n2408 4.5005
R18260 VSS.n2704 VSS.n2408 4.5005
R18261 VSS.n2706 VSS.n2408 4.5005
R18262 VSS.n2707 VSS.n2408 4.5005
R18263 VSS.n2709 VSS.n2408 4.5005
R18264 VSS.n2712 VSS.n2408 4.5005
R18265 VSS.n2714 VSS.n2408 4.5005
R18266 VSS.n2715 VSS.n2408 4.5005
R18267 VSS.n2717 VSS.n2408 4.5005
R18268 VSS.n2720 VSS.n2408 4.5005
R18269 VSS.n2722 VSS.n2408 4.5005
R18270 VSS.n2723 VSS.n2408 4.5005
R18271 VSS.n2725 VSS.n2408 4.5005
R18272 VSS.n2793 VSS.n2408 4.5005
R18273 VSS.n2859 VSS.n2408 4.5005
R18274 VSS.n3051 VSS.n2424 4.5005
R18275 VSS.n2424 VSS.n2351 4.5005
R18276 VSS.n2483 VSS.n2424 4.5005
R18277 VSS.n2484 VSS.n2424 4.5005
R18278 VSS.n2486 VSS.n2424 4.5005
R18279 VSS.n2489 VSS.n2424 4.5005
R18280 VSS.n2491 VSS.n2424 4.5005
R18281 VSS.n2492 VSS.n2424 4.5005
R18282 VSS.n2494 VSS.n2424 4.5005
R18283 VSS.n2497 VSS.n2424 4.5005
R18284 VSS.n2499 VSS.n2424 4.5005
R18285 VSS.n2500 VSS.n2424 4.5005
R18286 VSS.n2502 VSS.n2424 4.5005
R18287 VSS.n2505 VSS.n2424 4.5005
R18288 VSS.n2507 VSS.n2424 4.5005
R18289 VSS.n2508 VSS.n2424 4.5005
R18290 VSS.n2510 VSS.n2424 4.5005
R18291 VSS.n2513 VSS.n2424 4.5005
R18292 VSS.n2515 VSS.n2424 4.5005
R18293 VSS.n2516 VSS.n2424 4.5005
R18294 VSS.n2518 VSS.n2424 4.5005
R18295 VSS.n2521 VSS.n2424 4.5005
R18296 VSS.n2523 VSS.n2424 4.5005
R18297 VSS.n2524 VSS.n2424 4.5005
R18298 VSS.n2526 VSS.n2424 4.5005
R18299 VSS.n2529 VSS.n2424 4.5005
R18300 VSS.n2531 VSS.n2424 4.5005
R18301 VSS.n2532 VSS.n2424 4.5005
R18302 VSS.n2534 VSS.n2424 4.5005
R18303 VSS.n2537 VSS.n2424 4.5005
R18304 VSS.n2539 VSS.n2424 4.5005
R18305 VSS.n2540 VSS.n2424 4.5005
R18306 VSS.n2542 VSS.n2424 4.5005
R18307 VSS.n2545 VSS.n2424 4.5005
R18308 VSS.n2547 VSS.n2424 4.5005
R18309 VSS.n2548 VSS.n2424 4.5005
R18310 VSS.n2550 VSS.n2424 4.5005
R18311 VSS.n2553 VSS.n2424 4.5005
R18312 VSS.n2555 VSS.n2424 4.5005
R18313 VSS.n2556 VSS.n2424 4.5005
R18314 VSS.n2558 VSS.n2424 4.5005
R18315 VSS.n2561 VSS.n2424 4.5005
R18316 VSS.n2563 VSS.n2424 4.5005
R18317 VSS.n2564 VSS.n2424 4.5005
R18318 VSS.n2566 VSS.n2424 4.5005
R18319 VSS.n2569 VSS.n2424 4.5005
R18320 VSS.n2571 VSS.n2424 4.5005
R18321 VSS.n2572 VSS.n2424 4.5005
R18322 VSS.n2574 VSS.n2424 4.5005
R18323 VSS.n2577 VSS.n2424 4.5005
R18324 VSS.n2579 VSS.n2424 4.5005
R18325 VSS.n2580 VSS.n2424 4.5005
R18326 VSS.n2582 VSS.n2424 4.5005
R18327 VSS.n2585 VSS.n2424 4.5005
R18328 VSS.n2587 VSS.n2424 4.5005
R18329 VSS.n2588 VSS.n2424 4.5005
R18330 VSS.n2590 VSS.n2424 4.5005
R18331 VSS.n2593 VSS.n2424 4.5005
R18332 VSS.n2595 VSS.n2424 4.5005
R18333 VSS.n2596 VSS.n2424 4.5005
R18334 VSS.n2598 VSS.n2424 4.5005
R18335 VSS.n2601 VSS.n2424 4.5005
R18336 VSS.n2603 VSS.n2424 4.5005
R18337 VSS.n2604 VSS.n2424 4.5005
R18338 VSS.n2606 VSS.n2424 4.5005
R18339 VSS.n2609 VSS.n2424 4.5005
R18340 VSS.n2611 VSS.n2424 4.5005
R18341 VSS.n2612 VSS.n2424 4.5005
R18342 VSS.n2614 VSS.n2424 4.5005
R18343 VSS.n2617 VSS.n2424 4.5005
R18344 VSS.n2619 VSS.n2424 4.5005
R18345 VSS.n2620 VSS.n2424 4.5005
R18346 VSS.n2622 VSS.n2424 4.5005
R18347 VSS.n2625 VSS.n2424 4.5005
R18348 VSS.n2627 VSS.n2424 4.5005
R18349 VSS.n2628 VSS.n2424 4.5005
R18350 VSS.n2630 VSS.n2424 4.5005
R18351 VSS.n2633 VSS.n2424 4.5005
R18352 VSS.n2635 VSS.n2424 4.5005
R18353 VSS.n2636 VSS.n2424 4.5005
R18354 VSS.n2638 VSS.n2424 4.5005
R18355 VSS.n2640 VSS.n2424 4.5005
R18356 VSS.n2642 VSS.n2424 4.5005
R18357 VSS.n2643 VSS.n2424 4.5005
R18358 VSS.n2645 VSS.n2424 4.5005
R18359 VSS.n2648 VSS.n2424 4.5005
R18360 VSS.n2650 VSS.n2424 4.5005
R18361 VSS.n2651 VSS.n2424 4.5005
R18362 VSS.n2653 VSS.n2424 4.5005
R18363 VSS.n2656 VSS.n2424 4.5005
R18364 VSS.n2658 VSS.n2424 4.5005
R18365 VSS.n2659 VSS.n2424 4.5005
R18366 VSS.n2661 VSS.n2424 4.5005
R18367 VSS.n2664 VSS.n2424 4.5005
R18368 VSS.n2666 VSS.n2424 4.5005
R18369 VSS.n2667 VSS.n2424 4.5005
R18370 VSS.n2669 VSS.n2424 4.5005
R18371 VSS.n2672 VSS.n2424 4.5005
R18372 VSS.n2674 VSS.n2424 4.5005
R18373 VSS.n2675 VSS.n2424 4.5005
R18374 VSS.n2677 VSS.n2424 4.5005
R18375 VSS.n2680 VSS.n2424 4.5005
R18376 VSS.n2682 VSS.n2424 4.5005
R18377 VSS.n2683 VSS.n2424 4.5005
R18378 VSS.n2685 VSS.n2424 4.5005
R18379 VSS.n2688 VSS.n2424 4.5005
R18380 VSS.n2690 VSS.n2424 4.5005
R18381 VSS.n2691 VSS.n2424 4.5005
R18382 VSS.n2693 VSS.n2424 4.5005
R18383 VSS.n2696 VSS.n2424 4.5005
R18384 VSS.n2698 VSS.n2424 4.5005
R18385 VSS.n2699 VSS.n2424 4.5005
R18386 VSS.n2701 VSS.n2424 4.5005
R18387 VSS.n2704 VSS.n2424 4.5005
R18388 VSS.n2706 VSS.n2424 4.5005
R18389 VSS.n2707 VSS.n2424 4.5005
R18390 VSS.n2709 VSS.n2424 4.5005
R18391 VSS.n2712 VSS.n2424 4.5005
R18392 VSS.n2714 VSS.n2424 4.5005
R18393 VSS.n2715 VSS.n2424 4.5005
R18394 VSS.n2717 VSS.n2424 4.5005
R18395 VSS.n2720 VSS.n2424 4.5005
R18396 VSS.n2722 VSS.n2424 4.5005
R18397 VSS.n2723 VSS.n2424 4.5005
R18398 VSS.n2725 VSS.n2424 4.5005
R18399 VSS.n2793 VSS.n2424 4.5005
R18400 VSS.n2859 VSS.n2424 4.5005
R18401 VSS.n3051 VSS.n2407 4.5005
R18402 VSS.n2407 VSS.n2351 4.5005
R18403 VSS.n2483 VSS.n2407 4.5005
R18404 VSS.n2484 VSS.n2407 4.5005
R18405 VSS.n2486 VSS.n2407 4.5005
R18406 VSS.n2489 VSS.n2407 4.5005
R18407 VSS.n2491 VSS.n2407 4.5005
R18408 VSS.n2492 VSS.n2407 4.5005
R18409 VSS.n2494 VSS.n2407 4.5005
R18410 VSS.n2497 VSS.n2407 4.5005
R18411 VSS.n2499 VSS.n2407 4.5005
R18412 VSS.n2500 VSS.n2407 4.5005
R18413 VSS.n2502 VSS.n2407 4.5005
R18414 VSS.n2505 VSS.n2407 4.5005
R18415 VSS.n2507 VSS.n2407 4.5005
R18416 VSS.n2508 VSS.n2407 4.5005
R18417 VSS.n2510 VSS.n2407 4.5005
R18418 VSS.n2513 VSS.n2407 4.5005
R18419 VSS.n2515 VSS.n2407 4.5005
R18420 VSS.n2516 VSS.n2407 4.5005
R18421 VSS.n2518 VSS.n2407 4.5005
R18422 VSS.n2521 VSS.n2407 4.5005
R18423 VSS.n2523 VSS.n2407 4.5005
R18424 VSS.n2524 VSS.n2407 4.5005
R18425 VSS.n2526 VSS.n2407 4.5005
R18426 VSS.n2529 VSS.n2407 4.5005
R18427 VSS.n2531 VSS.n2407 4.5005
R18428 VSS.n2532 VSS.n2407 4.5005
R18429 VSS.n2534 VSS.n2407 4.5005
R18430 VSS.n2537 VSS.n2407 4.5005
R18431 VSS.n2539 VSS.n2407 4.5005
R18432 VSS.n2540 VSS.n2407 4.5005
R18433 VSS.n2542 VSS.n2407 4.5005
R18434 VSS.n2545 VSS.n2407 4.5005
R18435 VSS.n2547 VSS.n2407 4.5005
R18436 VSS.n2548 VSS.n2407 4.5005
R18437 VSS.n2550 VSS.n2407 4.5005
R18438 VSS.n2553 VSS.n2407 4.5005
R18439 VSS.n2555 VSS.n2407 4.5005
R18440 VSS.n2556 VSS.n2407 4.5005
R18441 VSS.n2558 VSS.n2407 4.5005
R18442 VSS.n2561 VSS.n2407 4.5005
R18443 VSS.n2563 VSS.n2407 4.5005
R18444 VSS.n2564 VSS.n2407 4.5005
R18445 VSS.n2566 VSS.n2407 4.5005
R18446 VSS.n2569 VSS.n2407 4.5005
R18447 VSS.n2571 VSS.n2407 4.5005
R18448 VSS.n2572 VSS.n2407 4.5005
R18449 VSS.n2574 VSS.n2407 4.5005
R18450 VSS.n2577 VSS.n2407 4.5005
R18451 VSS.n2579 VSS.n2407 4.5005
R18452 VSS.n2580 VSS.n2407 4.5005
R18453 VSS.n2582 VSS.n2407 4.5005
R18454 VSS.n2585 VSS.n2407 4.5005
R18455 VSS.n2587 VSS.n2407 4.5005
R18456 VSS.n2588 VSS.n2407 4.5005
R18457 VSS.n2590 VSS.n2407 4.5005
R18458 VSS.n2593 VSS.n2407 4.5005
R18459 VSS.n2595 VSS.n2407 4.5005
R18460 VSS.n2596 VSS.n2407 4.5005
R18461 VSS.n2598 VSS.n2407 4.5005
R18462 VSS.n2601 VSS.n2407 4.5005
R18463 VSS.n2603 VSS.n2407 4.5005
R18464 VSS.n2604 VSS.n2407 4.5005
R18465 VSS.n2606 VSS.n2407 4.5005
R18466 VSS.n2609 VSS.n2407 4.5005
R18467 VSS.n2611 VSS.n2407 4.5005
R18468 VSS.n2612 VSS.n2407 4.5005
R18469 VSS.n2614 VSS.n2407 4.5005
R18470 VSS.n2617 VSS.n2407 4.5005
R18471 VSS.n2619 VSS.n2407 4.5005
R18472 VSS.n2620 VSS.n2407 4.5005
R18473 VSS.n2622 VSS.n2407 4.5005
R18474 VSS.n2625 VSS.n2407 4.5005
R18475 VSS.n2627 VSS.n2407 4.5005
R18476 VSS.n2628 VSS.n2407 4.5005
R18477 VSS.n2630 VSS.n2407 4.5005
R18478 VSS.n2633 VSS.n2407 4.5005
R18479 VSS.n2635 VSS.n2407 4.5005
R18480 VSS.n2636 VSS.n2407 4.5005
R18481 VSS.n2638 VSS.n2407 4.5005
R18482 VSS.n2640 VSS.n2407 4.5005
R18483 VSS.n2642 VSS.n2407 4.5005
R18484 VSS.n2643 VSS.n2407 4.5005
R18485 VSS.n2645 VSS.n2407 4.5005
R18486 VSS.n2648 VSS.n2407 4.5005
R18487 VSS.n2650 VSS.n2407 4.5005
R18488 VSS.n2651 VSS.n2407 4.5005
R18489 VSS.n2653 VSS.n2407 4.5005
R18490 VSS.n2656 VSS.n2407 4.5005
R18491 VSS.n2658 VSS.n2407 4.5005
R18492 VSS.n2659 VSS.n2407 4.5005
R18493 VSS.n2661 VSS.n2407 4.5005
R18494 VSS.n2664 VSS.n2407 4.5005
R18495 VSS.n2666 VSS.n2407 4.5005
R18496 VSS.n2667 VSS.n2407 4.5005
R18497 VSS.n2669 VSS.n2407 4.5005
R18498 VSS.n2672 VSS.n2407 4.5005
R18499 VSS.n2674 VSS.n2407 4.5005
R18500 VSS.n2675 VSS.n2407 4.5005
R18501 VSS.n2677 VSS.n2407 4.5005
R18502 VSS.n2680 VSS.n2407 4.5005
R18503 VSS.n2682 VSS.n2407 4.5005
R18504 VSS.n2683 VSS.n2407 4.5005
R18505 VSS.n2685 VSS.n2407 4.5005
R18506 VSS.n2688 VSS.n2407 4.5005
R18507 VSS.n2690 VSS.n2407 4.5005
R18508 VSS.n2691 VSS.n2407 4.5005
R18509 VSS.n2693 VSS.n2407 4.5005
R18510 VSS.n2696 VSS.n2407 4.5005
R18511 VSS.n2698 VSS.n2407 4.5005
R18512 VSS.n2699 VSS.n2407 4.5005
R18513 VSS.n2701 VSS.n2407 4.5005
R18514 VSS.n2704 VSS.n2407 4.5005
R18515 VSS.n2706 VSS.n2407 4.5005
R18516 VSS.n2707 VSS.n2407 4.5005
R18517 VSS.n2709 VSS.n2407 4.5005
R18518 VSS.n2712 VSS.n2407 4.5005
R18519 VSS.n2714 VSS.n2407 4.5005
R18520 VSS.n2715 VSS.n2407 4.5005
R18521 VSS.n2717 VSS.n2407 4.5005
R18522 VSS.n2720 VSS.n2407 4.5005
R18523 VSS.n2722 VSS.n2407 4.5005
R18524 VSS.n2723 VSS.n2407 4.5005
R18525 VSS.n2725 VSS.n2407 4.5005
R18526 VSS.n2793 VSS.n2407 4.5005
R18527 VSS.n2859 VSS.n2407 4.5005
R18528 VSS.n3051 VSS.n2425 4.5005
R18529 VSS.n2425 VSS.n2351 4.5005
R18530 VSS.n2483 VSS.n2425 4.5005
R18531 VSS.n2484 VSS.n2425 4.5005
R18532 VSS.n2486 VSS.n2425 4.5005
R18533 VSS.n2489 VSS.n2425 4.5005
R18534 VSS.n2491 VSS.n2425 4.5005
R18535 VSS.n2492 VSS.n2425 4.5005
R18536 VSS.n2494 VSS.n2425 4.5005
R18537 VSS.n2497 VSS.n2425 4.5005
R18538 VSS.n2499 VSS.n2425 4.5005
R18539 VSS.n2500 VSS.n2425 4.5005
R18540 VSS.n2502 VSS.n2425 4.5005
R18541 VSS.n2505 VSS.n2425 4.5005
R18542 VSS.n2507 VSS.n2425 4.5005
R18543 VSS.n2508 VSS.n2425 4.5005
R18544 VSS.n2510 VSS.n2425 4.5005
R18545 VSS.n2513 VSS.n2425 4.5005
R18546 VSS.n2515 VSS.n2425 4.5005
R18547 VSS.n2516 VSS.n2425 4.5005
R18548 VSS.n2518 VSS.n2425 4.5005
R18549 VSS.n2521 VSS.n2425 4.5005
R18550 VSS.n2523 VSS.n2425 4.5005
R18551 VSS.n2524 VSS.n2425 4.5005
R18552 VSS.n2526 VSS.n2425 4.5005
R18553 VSS.n2529 VSS.n2425 4.5005
R18554 VSS.n2531 VSS.n2425 4.5005
R18555 VSS.n2532 VSS.n2425 4.5005
R18556 VSS.n2534 VSS.n2425 4.5005
R18557 VSS.n2537 VSS.n2425 4.5005
R18558 VSS.n2539 VSS.n2425 4.5005
R18559 VSS.n2540 VSS.n2425 4.5005
R18560 VSS.n2542 VSS.n2425 4.5005
R18561 VSS.n2545 VSS.n2425 4.5005
R18562 VSS.n2547 VSS.n2425 4.5005
R18563 VSS.n2548 VSS.n2425 4.5005
R18564 VSS.n2550 VSS.n2425 4.5005
R18565 VSS.n2553 VSS.n2425 4.5005
R18566 VSS.n2555 VSS.n2425 4.5005
R18567 VSS.n2556 VSS.n2425 4.5005
R18568 VSS.n2558 VSS.n2425 4.5005
R18569 VSS.n2561 VSS.n2425 4.5005
R18570 VSS.n2563 VSS.n2425 4.5005
R18571 VSS.n2564 VSS.n2425 4.5005
R18572 VSS.n2566 VSS.n2425 4.5005
R18573 VSS.n2569 VSS.n2425 4.5005
R18574 VSS.n2571 VSS.n2425 4.5005
R18575 VSS.n2572 VSS.n2425 4.5005
R18576 VSS.n2574 VSS.n2425 4.5005
R18577 VSS.n2577 VSS.n2425 4.5005
R18578 VSS.n2579 VSS.n2425 4.5005
R18579 VSS.n2580 VSS.n2425 4.5005
R18580 VSS.n2582 VSS.n2425 4.5005
R18581 VSS.n2585 VSS.n2425 4.5005
R18582 VSS.n2587 VSS.n2425 4.5005
R18583 VSS.n2588 VSS.n2425 4.5005
R18584 VSS.n2590 VSS.n2425 4.5005
R18585 VSS.n2593 VSS.n2425 4.5005
R18586 VSS.n2595 VSS.n2425 4.5005
R18587 VSS.n2596 VSS.n2425 4.5005
R18588 VSS.n2598 VSS.n2425 4.5005
R18589 VSS.n2601 VSS.n2425 4.5005
R18590 VSS.n2603 VSS.n2425 4.5005
R18591 VSS.n2604 VSS.n2425 4.5005
R18592 VSS.n2606 VSS.n2425 4.5005
R18593 VSS.n2609 VSS.n2425 4.5005
R18594 VSS.n2611 VSS.n2425 4.5005
R18595 VSS.n2612 VSS.n2425 4.5005
R18596 VSS.n2614 VSS.n2425 4.5005
R18597 VSS.n2617 VSS.n2425 4.5005
R18598 VSS.n2619 VSS.n2425 4.5005
R18599 VSS.n2620 VSS.n2425 4.5005
R18600 VSS.n2622 VSS.n2425 4.5005
R18601 VSS.n2625 VSS.n2425 4.5005
R18602 VSS.n2627 VSS.n2425 4.5005
R18603 VSS.n2628 VSS.n2425 4.5005
R18604 VSS.n2630 VSS.n2425 4.5005
R18605 VSS.n2633 VSS.n2425 4.5005
R18606 VSS.n2635 VSS.n2425 4.5005
R18607 VSS.n2636 VSS.n2425 4.5005
R18608 VSS.n2638 VSS.n2425 4.5005
R18609 VSS.n2640 VSS.n2425 4.5005
R18610 VSS.n2642 VSS.n2425 4.5005
R18611 VSS.n2643 VSS.n2425 4.5005
R18612 VSS.n2645 VSS.n2425 4.5005
R18613 VSS.n2648 VSS.n2425 4.5005
R18614 VSS.n2650 VSS.n2425 4.5005
R18615 VSS.n2651 VSS.n2425 4.5005
R18616 VSS.n2653 VSS.n2425 4.5005
R18617 VSS.n2656 VSS.n2425 4.5005
R18618 VSS.n2658 VSS.n2425 4.5005
R18619 VSS.n2659 VSS.n2425 4.5005
R18620 VSS.n2661 VSS.n2425 4.5005
R18621 VSS.n2664 VSS.n2425 4.5005
R18622 VSS.n2666 VSS.n2425 4.5005
R18623 VSS.n2667 VSS.n2425 4.5005
R18624 VSS.n2669 VSS.n2425 4.5005
R18625 VSS.n2672 VSS.n2425 4.5005
R18626 VSS.n2674 VSS.n2425 4.5005
R18627 VSS.n2675 VSS.n2425 4.5005
R18628 VSS.n2677 VSS.n2425 4.5005
R18629 VSS.n2680 VSS.n2425 4.5005
R18630 VSS.n2682 VSS.n2425 4.5005
R18631 VSS.n2683 VSS.n2425 4.5005
R18632 VSS.n2685 VSS.n2425 4.5005
R18633 VSS.n2688 VSS.n2425 4.5005
R18634 VSS.n2690 VSS.n2425 4.5005
R18635 VSS.n2691 VSS.n2425 4.5005
R18636 VSS.n2693 VSS.n2425 4.5005
R18637 VSS.n2696 VSS.n2425 4.5005
R18638 VSS.n2698 VSS.n2425 4.5005
R18639 VSS.n2699 VSS.n2425 4.5005
R18640 VSS.n2701 VSS.n2425 4.5005
R18641 VSS.n2704 VSS.n2425 4.5005
R18642 VSS.n2706 VSS.n2425 4.5005
R18643 VSS.n2707 VSS.n2425 4.5005
R18644 VSS.n2709 VSS.n2425 4.5005
R18645 VSS.n2712 VSS.n2425 4.5005
R18646 VSS.n2714 VSS.n2425 4.5005
R18647 VSS.n2715 VSS.n2425 4.5005
R18648 VSS.n2717 VSS.n2425 4.5005
R18649 VSS.n2720 VSS.n2425 4.5005
R18650 VSS.n2722 VSS.n2425 4.5005
R18651 VSS.n2723 VSS.n2425 4.5005
R18652 VSS.n2725 VSS.n2425 4.5005
R18653 VSS.n2793 VSS.n2425 4.5005
R18654 VSS.n2859 VSS.n2425 4.5005
R18655 VSS.n3051 VSS.n2406 4.5005
R18656 VSS.n2406 VSS.n2351 4.5005
R18657 VSS.n2483 VSS.n2406 4.5005
R18658 VSS.n2484 VSS.n2406 4.5005
R18659 VSS.n2486 VSS.n2406 4.5005
R18660 VSS.n2489 VSS.n2406 4.5005
R18661 VSS.n2491 VSS.n2406 4.5005
R18662 VSS.n2492 VSS.n2406 4.5005
R18663 VSS.n2494 VSS.n2406 4.5005
R18664 VSS.n2497 VSS.n2406 4.5005
R18665 VSS.n2499 VSS.n2406 4.5005
R18666 VSS.n2500 VSS.n2406 4.5005
R18667 VSS.n2502 VSS.n2406 4.5005
R18668 VSS.n2505 VSS.n2406 4.5005
R18669 VSS.n2507 VSS.n2406 4.5005
R18670 VSS.n2508 VSS.n2406 4.5005
R18671 VSS.n2510 VSS.n2406 4.5005
R18672 VSS.n2513 VSS.n2406 4.5005
R18673 VSS.n2515 VSS.n2406 4.5005
R18674 VSS.n2516 VSS.n2406 4.5005
R18675 VSS.n2518 VSS.n2406 4.5005
R18676 VSS.n2521 VSS.n2406 4.5005
R18677 VSS.n2523 VSS.n2406 4.5005
R18678 VSS.n2524 VSS.n2406 4.5005
R18679 VSS.n2526 VSS.n2406 4.5005
R18680 VSS.n2529 VSS.n2406 4.5005
R18681 VSS.n2531 VSS.n2406 4.5005
R18682 VSS.n2532 VSS.n2406 4.5005
R18683 VSS.n2534 VSS.n2406 4.5005
R18684 VSS.n2537 VSS.n2406 4.5005
R18685 VSS.n2539 VSS.n2406 4.5005
R18686 VSS.n2540 VSS.n2406 4.5005
R18687 VSS.n2542 VSS.n2406 4.5005
R18688 VSS.n2545 VSS.n2406 4.5005
R18689 VSS.n2547 VSS.n2406 4.5005
R18690 VSS.n2548 VSS.n2406 4.5005
R18691 VSS.n2550 VSS.n2406 4.5005
R18692 VSS.n2553 VSS.n2406 4.5005
R18693 VSS.n2555 VSS.n2406 4.5005
R18694 VSS.n2556 VSS.n2406 4.5005
R18695 VSS.n2558 VSS.n2406 4.5005
R18696 VSS.n2561 VSS.n2406 4.5005
R18697 VSS.n2563 VSS.n2406 4.5005
R18698 VSS.n2564 VSS.n2406 4.5005
R18699 VSS.n2566 VSS.n2406 4.5005
R18700 VSS.n2569 VSS.n2406 4.5005
R18701 VSS.n2571 VSS.n2406 4.5005
R18702 VSS.n2572 VSS.n2406 4.5005
R18703 VSS.n2574 VSS.n2406 4.5005
R18704 VSS.n2577 VSS.n2406 4.5005
R18705 VSS.n2579 VSS.n2406 4.5005
R18706 VSS.n2580 VSS.n2406 4.5005
R18707 VSS.n2582 VSS.n2406 4.5005
R18708 VSS.n2585 VSS.n2406 4.5005
R18709 VSS.n2587 VSS.n2406 4.5005
R18710 VSS.n2588 VSS.n2406 4.5005
R18711 VSS.n2590 VSS.n2406 4.5005
R18712 VSS.n2593 VSS.n2406 4.5005
R18713 VSS.n2595 VSS.n2406 4.5005
R18714 VSS.n2596 VSS.n2406 4.5005
R18715 VSS.n2598 VSS.n2406 4.5005
R18716 VSS.n2601 VSS.n2406 4.5005
R18717 VSS.n2603 VSS.n2406 4.5005
R18718 VSS.n2604 VSS.n2406 4.5005
R18719 VSS.n2606 VSS.n2406 4.5005
R18720 VSS.n2609 VSS.n2406 4.5005
R18721 VSS.n2611 VSS.n2406 4.5005
R18722 VSS.n2612 VSS.n2406 4.5005
R18723 VSS.n2614 VSS.n2406 4.5005
R18724 VSS.n2617 VSS.n2406 4.5005
R18725 VSS.n2619 VSS.n2406 4.5005
R18726 VSS.n2620 VSS.n2406 4.5005
R18727 VSS.n2622 VSS.n2406 4.5005
R18728 VSS.n2625 VSS.n2406 4.5005
R18729 VSS.n2627 VSS.n2406 4.5005
R18730 VSS.n2628 VSS.n2406 4.5005
R18731 VSS.n2630 VSS.n2406 4.5005
R18732 VSS.n2633 VSS.n2406 4.5005
R18733 VSS.n2635 VSS.n2406 4.5005
R18734 VSS.n2636 VSS.n2406 4.5005
R18735 VSS.n2638 VSS.n2406 4.5005
R18736 VSS.n2640 VSS.n2406 4.5005
R18737 VSS.n2642 VSS.n2406 4.5005
R18738 VSS.n2643 VSS.n2406 4.5005
R18739 VSS.n2645 VSS.n2406 4.5005
R18740 VSS.n2648 VSS.n2406 4.5005
R18741 VSS.n2650 VSS.n2406 4.5005
R18742 VSS.n2651 VSS.n2406 4.5005
R18743 VSS.n2653 VSS.n2406 4.5005
R18744 VSS.n2656 VSS.n2406 4.5005
R18745 VSS.n2658 VSS.n2406 4.5005
R18746 VSS.n2659 VSS.n2406 4.5005
R18747 VSS.n2661 VSS.n2406 4.5005
R18748 VSS.n2664 VSS.n2406 4.5005
R18749 VSS.n2666 VSS.n2406 4.5005
R18750 VSS.n2667 VSS.n2406 4.5005
R18751 VSS.n2669 VSS.n2406 4.5005
R18752 VSS.n2672 VSS.n2406 4.5005
R18753 VSS.n2674 VSS.n2406 4.5005
R18754 VSS.n2675 VSS.n2406 4.5005
R18755 VSS.n2677 VSS.n2406 4.5005
R18756 VSS.n2680 VSS.n2406 4.5005
R18757 VSS.n2682 VSS.n2406 4.5005
R18758 VSS.n2683 VSS.n2406 4.5005
R18759 VSS.n2685 VSS.n2406 4.5005
R18760 VSS.n2688 VSS.n2406 4.5005
R18761 VSS.n2690 VSS.n2406 4.5005
R18762 VSS.n2691 VSS.n2406 4.5005
R18763 VSS.n2693 VSS.n2406 4.5005
R18764 VSS.n2696 VSS.n2406 4.5005
R18765 VSS.n2698 VSS.n2406 4.5005
R18766 VSS.n2699 VSS.n2406 4.5005
R18767 VSS.n2701 VSS.n2406 4.5005
R18768 VSS.n2704 VSS.n2406 4.5005
R18769 VSS.n2706 VSS.n2406 4.5005
R18770 VSS.n2707 VSS.n2406 4.5005
R18771 VSS.n2709 VSS.n2406 4.5005
R18772 VSS.n2712 VSS.n2406 4.5005
R18773 VSS.n2714 VSS.n2406 4.5005
R18774 VSS.n2715 VSS.n2406 4.5005
R18775 VSS.n2717 VSS.n2406 4.5005
R18776 VSS.n2720 VSS.n2406 4.5005
R18777 VSS.n2722 VSS.n2406 4.5005
R18778 VSS.n2723 VSS.n2406 4.5005
R18779 VSS.n2725 VSS.n2406 4.5005
R18780 VSS.n2793 VSS.n2406 4.5005
R18781 VSS.n2859 VSS.n2406 4.5005
R18782 VSS.n3051 VSS.n2426 4.5005
R18783 VSS.n2426 VSS.n2351 4.5005
R18784 VSS.n2483 VSS.n2426 4.5005
R18785 VSS.n2484 VSS.n2426 4.5005
R18786 VSS.n2486 VSS.n2426 4.5005
R18787 VSS.n2489 VSS.n2426 4.5005
R18788 VSS.n2491 VSS.n2426 4.5005
R18789 VSS.n2492 VSS.n2426 4.5005
R18790 VSS.n2494 VSS.n2426 4.5005
R18791 VSS.n2497 VSS.n2426 4.5005
R18792 VSS.n2499 VSS.n2426 4.5005
R18793 VSS.n2500 VSS.n2426 4.5005
R18794 VSS.n2502 VSS.n2426 4.5005
R18795 VSS.n2505 VSS.n2426 4.5005
R18796 VSS.n2507 VSS.n2426 4.5005
R18797 VSS.n2508 VSS.n2426 4.5005
R18798 VSS.n2510 VSS.n2426 4.5005
R18799 VSS.n2513 VSS.n2426 4.5005
R18800 VSS.n2515 VSS.n2426 4.5005
R18801 VSS.n2516 VSS.n2426 4.5005
R18802 VSS.n2518 VSS.n2426 4.5005
R18803 VSS.n2521 VSS.n2426 4.5005
R18804 VSS.n2523 VSS.n2426 4.5005
R18805 VSS.n2524 VSS.n2426 4.5005
R18806 VSS.n2526 VSS.n2426 4.5005
R18807 VSS.n2529 VSS.n2426 4.5005
R18808 VSS.n2531 VSS.n2426 4.5005
R18809 VSS.n2532 VSS.n2426 4.5005
R18810 VSS.n2534 VSS.n2426 4.5005
R18811 VSS.n2537 VSS.n2426 4.5005
R18812 VSS.n2539 VSS.n2426 4.5005
R18813 VSS.n2540 VSS.n2426 4.5005
R18814 VSS.n2542 VSS.n2426 4.5005
R18815 VSS.n2545 VSS.n2426 4.5005
R18816 VSS.n2547 VSS.n2426 4.5005
R18817 VSS.n2548 VSS.n2426 4.5005
R18818 VSS.n2550 VSS.n2426 4.5005
R18819 VSS.n2553 VSS.n2426 4.5005
R18820 VSS.n2555 VSS.n2426 4.5005
R18821 VSS.n2556 VSS.n2426 4.5005
R18822 VSS.n2558 VSS.n2426 4.5005
R18823 VSS.n2561 VSS.n2426 4.5005
R18824 VSS.n2563 VSS.n2426 4.5005
R18825 VSS.n2564 VSS.n2426 4.5005
R18826 VSS.n2566 VSS.n2426 4.5005
R18827 VSS.n2569 VSS.n2426 4.5005
R18828 VSS.n2571 VSS.n2426 4.5005
R18829 VSS.n2572 VSS.n2426 4.5005
R18830 VSS.n2574 VSS.n2426 4.5005
R18831 VSS.n2577 VSS.n2426 4.5005
R18832 VSS.n2579 VSS.n2426 4.5005
R18833 VSS.n2580 VSS.n2426 4.5005
R18834 VSS.n2582 VSS.n2426 4.5005
R18835 VSS.n2585 VSS.n2426 4.5005
R18836 VSS.n2587 VSS.n2426 4.5005
R18837 VSS.n2588 VSS.n2426 4.5005
R18838 VSS.n2590 VSS.n2426 4.5005
R18839 VSS.n2593 VSS.n2426 4.5005
R18840 VSS.n2595 VSS.n2426 4.5005
R18841 VSS.n2596 VSS.n2426 4.5005
R18842 VSS.n2598 VSS.n2426 4.5005
R18843 VSS.n2601 VSS.n2426 4.5005
R18844 VSS.n2603 VSS.n2426 4.5005
R18845 VSS.n2604 VSS.n2426 4.5005
R18846 VSS.n2606 VSS.n2426 4.5005
R18847 VSS.n2609 VSS.n2426 4.5005
R18848 VSS.n2611 VSS.n2426 4.5005
R18849 VSS.n2612 VSS.n2426 4.5005
R18850 VSS.n2614 VSS.n2426 4.5005
R18851 VSS.n2617 VSS.n2426 4.5005
R18852 VSS.n2619 VSS.n2426 4.5005
R18853 VSS.n2620 VSS.n2426 4.5005
R18854 VSS.n2622 VSS.n2426 4.5005
R18855 VSS.n2625 VSS.n2426 4.5005
R18856 VSS.n2627 VSS.n2426 4.5005
R18857 VSS.n2628 VSS.n2426 4.5005
R18858 VSS.n2630 VSS.n2426 4.5005
R18859 VSS.n2633 VSS.n2426 4.5005
R18860 VSS.n2635 VSS.n2426 4.5005
R18861 VSS.n2636 VSS.n2426 4.5005
R18862 VSS.n2638 VSS.n2426 4.5005
R18863 VSS.n2640 VSS.n2426 4.5005
R18864 VSS.n2642 VSS.n2426 4.5005
R18865 VSS.n2643 VSS.n2426 4.5005
R18866 VSS.n2645 VSS.n2426 4.5005
R18867 VSS.n2648 VSS.n2426 4.5005
R18868 VSS.n2650 VSS.n2426 4.5005
R18869 VSS.n2651 VSS.n2426 4.5005
R18870 VSS.n2653 VSS.n2426 4.5005
R18871 VSS.n2656 VSS.n2426 4.5005
R18872 VSS.n2658 VSS.n2426 4.5005
R18873 VSS.n2659 VSS.n2426 4.5005
R18874 VSS.n2661 VSS.n2426 4.5005
R18875 VSS.n2664 VSS.n2426 4.5005
R18876 VSS.n2666 VSS.n2426 4.5005
R18877 VSS.n2667 VSS.n2426 4.5005
R18878 VSS.n2669 VSS.n2426 4.5005
R18879 VSS.n2672 VSS.n2426 4.5005
R18880 VSS.n2674 VSS.n2426 4.5005
R18881 VSS.n2675 VSS.n2426 4.5005
R18882 VSS.n2677 VSS.n2426 4.5005
R18883 VSS.n2680 VSS.n2426 4.5005
R18884 VSS.n2682 VSS.n2426 4.5005
R18885 VSS.n2683 VSS.n2426 4.5005
R18886 VSS.n2685 VSS.n2426 4.5005
R18887 VSS.n2688 VSS.n2426 4.5005
R18888 VSS.n2690 VSS.n2426 4.5005
R18889 VSS.n2691 VSS.n2426 4.5005
R18890 VSS.n2693 VSS.n2426 4.5005
R18891 VSS.n2696 VSS.n2426 4.5005
R18892 VSS.n2698 VSS.n2426 4.5005
R18893 VSS.n2699 VSS.n2426 4.5005
R18894 VSS.n2701 VSS.n2426 4.5005
R18895 VSS.n2704 VSS.n2426 4.5005
R18896 VSS.n2706 VSS.n2426 4.5005
R18897 VSS.n2707 VSS.n2426 4.5005
R18898 VSS.n2709 VSS.n2426 4.5005
R18899 VSS.n2712 VSS.n2426 4.5005
R18900 VSS.n2714 VSS.n2426 4.5005
R18901 VSS.n2715 VSS.n2426 4.5005
R18902 VSS.n2717 VSS.n2426 4.5005
R18903 VSS.n2720 VSS.n2426 4.5005
R18904 VSS.n2722 VSS.n2426 4.5005
R18905 VSS.n2723 VSS.n2426 4.5005
R18906 VSS.n2725 VSS.n2426 4.5005
R18907 VSS.n2793 VSS.n2426 4.5005
R18908 VSS.n2859 VSS.n2426 4.5005
R18909 VSS.n3051 VSS.n2405 4.5005
R18910 VSS.n2405 VSS.n2351 4.5005
R18911 VSS.n2483 VSS.n2405 4.5005
R18912 VSS.n2484 VSS.n2405 4.5005
R18913 VSS.n2486 VSS.n2405 4.5005
R18914 VSS.n2489 VSS.n2405 4.5005
R18915 VSS.n2491 VSS.n2405 4.5005
R18916 VSS.n2492 VSS.n2405 4.5005
R18917 VSS.n2494 VSS.n2405 4.5005
R18918 VSS.n2497 VSS.n2405 4.5005
R18919 VSS.n2499 VSS.n2405 4.5005
R18920 VSS.n2500 VSS.n2405 4.5005
R18921 VSS.n2502 VSS.n2405 4.5005
R18922 VSS.n2505 VSS.n2405 4.5005
R18923 VSS.n2507 VSS.n2405 4.5005
R18924 VSS.n2508 VSS.n2405 4.5005
R18925 VSS.n2510 VSS.n2405 4.5005
R18926 VSS.n2513 VSS.n2405 4.5005
R18927 VSS.n2515 VSS.n2405 4.5005
R18928 VSS.n2516 VSS.n2405 4.5005
R18929 VSS.n2518 VSS.n2405 4.5005
R18930 VSS.n2521 VSS.n2405 4.5005
R18931 VSS.n2523 VSS.n2405 4.5005
R18932 VSS.n2524 VSS.n2405 4.5005
R18933 VSS.n2526 VSS.n2405 4.5005
R18934 VSS.n2529 VSS.n2405 4.5005
R18935 VSS.n2531 VSS.n2405 4.5005
R18936 VSS.n2532 VSS.n2405 4.5005
R18937 VSS.n2534 VSS.n2405 4.5005
R18938 VSS.n2537 VSS.n2405 4.5005
R18939 VSS.n2539 VSS.n2405 4.5005
R18940 VSS.n2540 VSS.n2405 4.5005
R18941 VSS.n2542 VSS.n2405 4.5005
R18942 VSS.n2545 VSS.n2405 4.5005
R18943 VSS.n2547 VSS.n2405 4.5005
R18944 VSS.n2548 VSS.n2405 4.5005
R18945 VSS.n2550 VSS.n2405 4.5005
R18946 VSS.n2553 VSS.n2405 4.5005
R18947 VSS.n2555 VSS.n2405 4.5005
R18948 VSS.n2556 VSS.n2405 4.5005
R18949 VSS.n2558 VSS.n2405 4.5005
R18950 VSS.n2561 VSS.n2405 4.5005
R18951 VSS.n2563 VSS.n2405 4.5005
R18952 VSS.n2564 VSS.n2405 4.5005
R18953 VSS.n2566 VSS.n2405 4.5005
R18954 VSS.n2569 VSS.n2405 4.5005
R18955 VSS.n2571 VSS.n2405 4.5005
R18956 VSS.n2572 VSS.n2405 4.5005
R18957 VSS.n2574 VSS.n2405 4.5005
R18958 VSS.n2577 VSS.n2405 4.5005
R18959 VSS.n2579 VSS.n2405 4.5005
R18960 VSS.n2580 VSS.n2405 4.5005
R18961 VSS.n2582 VSS.n2405 4.5005
R18962 VSS.n2585 VSS.n2405 4.5005
R18963 VSS.n2587 VSS.n2405 4.5005
R18964 VSS.n2588 VSS.n2405 4.5005
R18965 VSS.n2590 VSS.n2405 4.5005
R18966 VSS.n2593 VSS.n2405 4.5005
R18967 VSS.n2595 VSS.n2405 4.5005
R18968 VSS.n2596 VSS.n2405 4.5005
R18969 VSS.n2598 VSS.n2405 4.5005
R18970 VSS.n2601 VSS.n2405 4.5005
R18971 VSS.n2603 VSS.n2405 4.5005
R18972 VSS.n2604 VSS.n2405 4.5005
R18973 VSS.n2606 VSS.n2405 4.5005
R18974 VSS.n2609 VSS.n2405 4.5005
R18975 VSS.n2611 VSS.n2405 4.5005
R18976 VSS.n2612 VSS.n2405 4.5005
R18977 VSS.n2614 VSS.n2405 4.5005
R18978 VSS.n2617 VSS.n2405 4.5005
R18979 VSS.n2619 VSS.n2405 4.5005
R18980 VSS.n2620 VSS.n2405 4.5005
R18981 VSS.n2622 VSS.n2405 4.5005
R18982 VSS.n2625 VSS.n2405 4.5005
R18983 VSS.n2627 VSS.n2405 4.5005
R18984 VSS.n2628 VSS.n2405 4.5005
R18985 VSS.n2630 VSS.n2405 4.5005
R18986 VSS.n2633 VSS.n2405 4.5005
R18987 VSS.n2635 VSS.n2405 4.5005
R18988 VSS.n2636 VSS.n2405 4.5005
R18989 VSS.n2638 VSS.n2405 4.5005
R18990 VSS.n2640 VSS.n2405 4.5005
R18991 VSS.n2642 VSS.n2405 4.5005
R18992 VSS.n2643 VSS.n2405 4.5005
R18993 VSS.n2645 VSS.n2405 4.5005
R18994 VSS.n2648 VSS.n2405 4.5005
R18995 VSS.n2650 VSS.n2405 4.5005
R18996 VSS.n2651 VSS.n2405 4.5005
R18997 VSS.n2653 VSS.n2405 4.5005
R18998 VSS.n2656 VSS.n2405 4.5005
R18999 VSS.n2658 VSS.n2405 4.5005
R19000 VSS.n2659 VSS.n2405 4.5005
R19001 VSS.n2661 VSS.n2405 4.5005
R19002 VSS.n2664 VSS.n2405 4.5005
R19003 VSS.n2666 VSS.n2405 4.5005
R19004 VSS.n2667 VSS.n2405 4.5005
R19005 VSS.n2669 VSS.n2405 4.5005
R19006 VSS.n2672 VSS.n2405 4.5005
R19007 VSS.n2674 VSS.n2405 4.5005
R19008 VSS.n2675 VSS.n2405 4.5005
R19009 VSS.n2677 VSS.n2405 4.5005
R19010 VSS.n2680 VSS.n2405 4.5005
R19011 VSS.n2682 VSS.n2405 4.5005
R19012 VSS.n2683 VSS.n2405 4.5005
R19013 VSS.n2685 VSS.n2405 4.5005
R19014 VSS.n2688 VSS.n2405 4.5005
R19015 VSS.n2690 VSS.n2405 4.5005
R19016 VSS.n2691 VSS.n2405 4.5005
R19017 VSS.n2693 VSS.n2405 4.5005
R19018 VSS.n2696 VSS.n2405 4.5005
R19019 VSS.n2698 VSS.n2405 4.5005
R19020 VSS.n2699 VSS.n2405 4.5005
R19021 VSS.n2701 VSS.n2405 4.5005
R19022 VSS.n2704 VSS.n2405 4.5005
R19023 VSS.n2706 VSS.n2405 4.5005
R19024 VSS.n2707 VSS.n2405 4.5005
R19025 VSS.n2709 VSS.n2405 4.5005
R19026 VSS.n2712 VSS.n2405 4.5005
R19027 VSS.n2714 VSS.n2405 4.5005
R19028 VSS.n2715 VSS.n2405 4.5005
R19029 VSS.n2717 VSS.n2405 4.5005
R19030 VSS.n2720 VSS.n2405 4.5005
R19031 VSS.n2722 VSS.n2405 4.5005
R19032 VSS.n2723 VSS.n2405 4.5005
R19033 VSS.n2725 VSS.n2405 4.5005
R19034 VSS.n2793 VSS.n2405 4.5005
R19035 VSS.n2859 VSS.n2405 4.5005
R19036 VSS.n3051 VSS.n2427 4.5005
R19037 VSS.n2427 VSS.n2351 4.5005
R19038 VSS.n2483 VSS.n2427 4.5005
R19039 VSS.n2484 VSS.n2427 4.5005
R19040 VSS.n2486 VSS.n2427 4.5005
R19041 VSS.n2489 VSS.n2427 4.5005
R19042 VSS.n2491 VSS.n2427 4.5005
R19043 VSS.n2492 VSS.n2427 4.5005
R19044 VSS.n2494 VSS.n2427 4.5005
R19045 VSS.n2497 VSS.n2427 4.5005
R19046 VSS.n2499 VSS.n2427 4.5005
R19047 VSS.n2500 VSS.n2427 4.5005
R19048 VSS.n2502 VSS.n2427 4.5005
R19049 VSS.n2505 VSS.n2427 4.5005
R19050 VSS.n2507 VSS.n2427 4.5005
R19051 VSS.n2508 VSS.n2427 4.5005
R19052 VSS.n2510 VSS.n2427 4.5005
R19053 VSS.n2513 VSS.n2427 4.5005
R19054 VSS.n2515 VSS.n2427 4.5005
R19055 VSS.n2516 VSS.n2427 4.5005
R19056 VSS.n2518 VSS.n2427 4.5005
R19057 VSS.n2521 VSS.n2427 4.5005
R19058 VSS.n2523 VSS.n2427 4.5005
R19059 VSS.n2524 VSS.n2427 4.5005
R19060 VSS.n2526 VSS.n2427 4.5005
R19061 VSS.n2529 VSS.n2427 4.5005
R19062 VSS.n2531 VSS.n2427 4.5005
R19063 VSS.n2532 VSS.n2427 4.5005
R19064 VSS.n2534 VSS.n2427 4.5005
R19065 VSS.n2537 VSS.n2427 4.5005
R19066 VSS.n2539 VSS.n2427 4.5005
R19067 VSS.n2540 VSS.n2427 4.5005
R19068 VSS.n2542 VSS.n2427 4.5005
R19069 VSS.n2545 VSS.n2427 4.5005
R19070 VSS.n2547 VSS.n2427 4.5005
R19071 VSS.n2548 VSS.n2427 4.5005
R19072 VSS.n2550 VSS.n2427 4.5005
R19073 VSS.n2553 VSS.n2427 4.5005
R19074 VSS.n2555 VSS.n2427 4.5005
R19075 VSS.n2556 VSS.n2427 4.5005
R19076 VSS.n2558 VSS.n2427 4.5005
R19077 VSS.n2561 VSS.n2427 4.5005
R19078 VSS.n2563 VSS.n2427 4.5005
R19079 VSS.n2564 VSS.n2427 4.5005
R19080 VSS.n2566 VSS.n2427 4.5005
R19081 VSS.n2569 VSS.n2427 4.5005
R19082 VSS.n2571 VSS.n2427 4.5005
R19083 VSS.n2572 VSS.n2427 4.5005
R19084 VSS.n2574 VSS.n2427 4.5005
R19085 VSS.n2577 VSS.n2427 4.5005
R19086 VSS.n2579 VSS.n2427 4.5005
R19087 VSS.n2580 VSS.n2427 4.5005
R19088 VSS.n2582 VSS.n2427 4.5005
R19089 VSS.n2585 VSS.n2427 4.5005
R19090 VSS.n2587 VSS.n2427 4.5005
R19091 VSS.n2588 VSS.n2427 4.5005
R19092 VSS.n2590 VSS.n2427 4.5005
R19093 VSS.n2593 VSS.n2427 4.5005
R19094 VSS.n2595 VSS.n2427 4.5005
R19095 VSS.n2596 VSS.n2427 4.5005
R19096 VSS.n2598 VSS.n2427 4.5005
R19097 VSS.n2601 VSS.n2427 4.5005
R19098 VSS.n2603 VSS.n2427 4.5005
R19099 VSS.n2604 VSS.n2427 4.5005
R19100 VSS.n2606 VSS.n2427 4.5005
R19101 VSS.n2609 VSS.n2427 4.5005
R19102 VSS.n2611 VSS.n2427 4.5005
R19103 VSS.n2612 VSS.n2427 4.5005
R19104 VSS.n2614 VSS.n2427 4.5005
R19105 VSS.n2617 VSS.n2427 4.5005
R19106 VSS.n2619 VSS.n2427 4.5005
R19107 VSS.n2620 VSS.n2427 4.5005
R19108 VSS.n2622 VSS.n2427 4.5005
R19109 VSS.n2625 VSS.n2427 4.5005
R19110 VSS.n2627 VSS.n2427 4.5005
R19111 VSS.n2628 VSS.n2427 4.5005
R19112 VSS.n2630 VSS.n2427 4.5005
R19113 VSS.n2633 VSS.n2427 4.5005
R19114 VSS.n2635 VSS.n2427 4.5005
R19115 VSS.n2636 VSS.n2427 4.5005
R19116 VSS.n2638 VSS.n2427 4.5005
R19117 VSS.n2640 VSS.n2427 4.5005
R19118 VSS.n2642 VSS.n2427 4.5005
R19119 VSS.n2643 VSS.n2427 4.5005
R19120 VSS.n2645 VSS.n2427 4.5005
R19121 VSS.n2648 VSS.n2427 4.5005
R19122 VSS.n2650 VSS.n2427 4.5005
R19123 VSS.n2651 VSS.n2427 4.5005
R19124 VSS.n2653 VSS.n2427 4.5005
R19125 VSS.n2656 VSS.n2427 4.5005
R19126 VSS.n2658 VSS.n2427 4.5005
R19127 VSS.n2659 VSS.n2427 4.5005
R19128 VSS.n2661 VSS.n2427 4.5005
R19129 VSS.n2664 VSS.n2427 4.5005
R19130 VSS.n2666 VSS.n2427 4.5005
R19131 VSS.n2667 VSS.n2427 4.5005
R19132 VSS.n2669 VSS.n2427 4.5005
R19133 VSS.n2672 VSS.n2427 4.5005
R19134 VSS.n2674 VSS.n2427 4.5005
R19135 VSS.n2675 VSS.n2427 4.5005
R19136 VSS.n2677 VSS.n2427 4.5005
R19137 VSS.n2680 VSS.n2427 4.5005
R19138 VSS.n2682 VSS.n2427 4.5005
R19139 VSS.n2683 VSS.n2427 4.5005
R19140 VSS.n2685 VSS.n2427 4.5005
R19141 VSS.n2688 VSS.n2427 4.5005
R19142 VSS.n2690 VSS.n2427 4.5005
R19143 VSS.n2691 VSS.n2427 4.5005
R19144 VSS.n2693 VSS.n2427 4.5005
R19145 VSS.n2696 VSS.n2427 4.5005
R19146 VSS.n2698 VSS.n2427 4.5005
R19147 VSS.n2699 VSS.n2427 4.5005
R19148 VSS.n2701 VSS.n2427 4.5005
R19149 VSS.n2704 VSS.n2427 4.5005
R19150 VSS.n2706 VSS.n2427 4.5005
R19151 VSS.n2707 VSS.n2427 4.5005
R19152 VSS.n2709 VSS.n2427 4.5005
R19153 VSS.n2712 VSS.n2427 4.5005
R19154 VSS.n2714 VSS.n2427 4.5005
R19155 VSS.n2715 VSS.n2427 4.5005
R19156 VSS.n2717 VSS.n2427 4.5005
R19157 VSS.n2720 VSS.n2427 4.5005
R19158 VSS.n2722 VSS.n2427 4.5005
R19159 VSS.n2723 VSS.n2427 4.5005
R19160 VSS.n2725 VSS.n2427 4.5005
R19161 VSS.n2793 VSS.n2427 4.5005
R19162 VSS.n2859 VSS.n2427 4.5005
R19163 VSS.n3051 VSS.n2404 4.5005
R19164 VSS.n2404 VSS.n2351 4.5005
R19165 VSS.n2483 VSS.n2404 4.5005
R19166 VSS.n2484 VSS.n2404 4.5005
R19167 VSS.n2486 VSS.n2404 4.5005
R19168 VSS.n2489 VSS.n2404 4.5005
R19169 VSS.n2491 VSS.n2404 4.5005
R19170 VSS.n2492 VSS.n2404 4.5005
R19171 VSS.n2494 VSS.n2404 4.5005
R19172 VSS.n2497 VSS.n2404 4.5005
R19173 VSS.n2499 VSS.n2404 4.5005
R19174 VSS.n2500 VSS.n2404 4.5005
R19175 VSS.n2502 VSS.n2404 4.5005
R19176 VSS.n2505 VSS.n2404 4.5005
R19177 VSS.n2507 VSS.n2404 4.5005
R19178 VSS.n2508 VSS.n2404 4.5005
R19179 VSS.n2510 VSS.n2404 4.5005
R19180 VSS.n2513 VSS.n2404 4.5005
R19181 VSS.n2515 VSS.n2404 4.5005
R19182 VSS.n2516 VSS.n2404 4.5005
R19183 VSS.n2518 VSS.n2404 4.5005
R19184 VSS.n2521 VSS.n2404 4.5005
R19185 VSS.n2523 VSS.n2404 4.5005
R19186 VSS.n2524 VSS.n2404 4.5005
R19187 VSS.n2526 VSS.n2404 4.5005
R19188 VSS.n2529 VSS.n2404 4.5005
R19189 VSS.n2531 VSS.n2404 4.5005
R19190 VSS.n2532 VSS.n2404 4.5005
R19191 VSS.n2534 VSS.n2404 4.5005
R19192 VSS.n2537 VSS.n2404 4.5005
R19193 VSS.n2539 VSS.n2404 4.5005
R19194 VSS.n2540 VSS.n2404 4.5005
R19195 VSS.n2542 VSS.n2404 4.5005
R19196 VSS.n2545 VSS.n2404 4.5005
R19197 VSS.n2547 VSS.n2404 4.5005
R19198 VSS.n2548 VSS.n2404 4.5005
R19199 VSS.n2550 VSS.n2404 4.5005
R19200 VSS.n2553 VSS.n2404 4.5005
R19201 VSS.n2555 VSS.n2404 4.5005
R19202 VSS.n2556 VSS.n2404 4.5005
R19203 VSS.n2558 VSS.n2404 4.5005
R19204 VSS.n2561 VSS.n2404 4.5005
R19205 VSS.n2563 VSS.n2404 4.5005
R19206 VSS.n2564 VSS.n2404 4.5005
R19207 VSS.n2566 VSS.n2404 4.5005
R19208 VSS.n2569 VSS.n2404 4.5005
R19209 VSS.n2571 VSS.n2404 4.5005
R19210 VSS.n2572 VSS.n2404 4.5005
R19211 VSS.n2574 VSS.n2404 4.5005
R19212 VSS.n2577 VSS.n2404 4.5005
R19213 VSS.n2579 VSS.n2404 4.5005
R19214 VSS.n2580 VSS.n2404 4.5005
R19215 VSS.n2582 VSS.n2404 4.5005
R19216 VSS.n2585 VSS.n2404 4.5005
R19217 VSS.n2587 VSS.n2404 4.5005
R19218 VSS.n2588 VSS.n2404 4.5005
R19219 VSS.n2590 VSS.n2404 4.5005
R19220 VSS.n2593 VSS.n2404 4.5005
R19221 VSS.n2595 VSS.n2404 4.5005
R19222 VSS.n2596 VSS.n2404 4.5005
R19223 VSS.n2598 VSS.n2404 4.5005
R19224 VSS.n2601 VSS.n2404 4.5005
R19225 VSS.n2603 VSS.n2404 4.5005
R19226 VSS.n2604 VSS.n2404 4.5005
R19227 VSS.n2606 VSS.n2404 4.5005
R19228 VSS.n2609 VSS.n2404 4.5005
R19229 VSS.n2611 VSS.n2404 4.5005
R19230 VSS.n2612 VSS.n2404 4.5005
R19231 VSS.n2614 VSS.n2404 4.5005
R19232 VSS.n2617 VSS.n2404 4.5005
R19233 VSS.n2619 VSS.n2404 4.5005
R19234 VSS.n2620 VSS.n2404 4.5005
R19235 VSS.n2622 VSS.n2404 4.5005
R19236 VSS.n2625 VSS.n2404 4.5005
R19237 VSS.n2627 VSS.n2404 4.5005
R19238 VSS.n2628 VSS.n2404 4.5005
R19239 VSS.n2630 VSS.n2404 4.5005
R19240 VSS.n2633 VSS.n2404 4.5005
R19241 VSS.n2635 VSS.n2404 4.5005
R19242 VSS.n2636 VSS.n2404 4.5005
R19243 VSS.n2638 VSS.n2404 4.5005
R19244 VSS.n2640 VSS.n2404 4.5005
R19245 VSS.n2642 VSS.n2404 4.5005
R19246 VSS.n2643 VSS.n2404 4.5005
R19247 VSS.n2645 VSS.n2404 4.5005
R19248 VSS.n2648 VSS.n2404 4.5005
R19249 VSS.n2650 VSS.n2404 4.5005
R19250 VSS.n2651 VSS.n2404 4.5005
R19251 VSS.n2653 VSS.n2404 4.5005
R19252 VSS.n2656 VSS.n2404 4.5005
R19253 VSS.n2658 VSS.n2404 4.5005
R19254 VSS.n2659 VSS.n2404 4.5005
R19255 VSS.n2661 VSS.n2404 4.5005
R19256 VSS.n2664 VSS.n2404 4.5005
R19257 VSS.n2666 VSS.n2404 4.5005
R19258 VSS.n2667 VSS.n2404 4.5005
R19259 VSS.n2669 VSS.n2404 4.5005
R19260 VSS.n2672 VSS.n2404 4.5005
R19261 VSS.n2674 VSS.n2404 4.5005
R19262 VSS.n2675 VSS.n2404 4.5005
R19263 VSS.n2677 VSS.n2404 4.5005
R19264 VSS.n2680 VSS.n2404 4.5005
R19265 VSS.n2682 VSS.n2404 4.5005
R19266 VSS.n2683 VSS.n2404 4.5005
R19267 VSS.n2685 VSS.n2404 4.5005
R19268 VSS.n2688 VSS.n2404 4.5005
R19269 VSS.n2690 VSS.n2404 4.5005
R19270 VSS.n2691 VSS.n2404 4.5005
R19271 VSS.n2693 VSS.n2404 4.5005
R19272 VSS.n2696 VSS.n2404 4.5005
R19273 VSS.n2698 VSS.n2404 4.5005
R19274 VSS.n2699 VSS.n2404 4.5005
R19275 VSS.n2701 VSS.n2404 4.5005
R19276 VSS.n2704 VSS.n2404 4.5005
R19277 VSS.n2706 VSS.n2404 4.5005
R19278 VSS.n2707 VSS.n2404 4.5005
R19279 VSS.n2709 VSS.n2404 4.5005
R19280 VSS.n2712 VSS.n2404 4.5005
R19281 VSS.n2714 VSS.n2404 4.5005
R19282 VSS.n2715 VSS.n2404 4.5005
R19283 VSS.n2717 VSS.n2404 4.5005
R19284 VSS.n2720 VSS.n2404 4.5005
R19285 VSS.n2722 VSS.n2404 4.5005
R19286 VSS.n2723 VSS.n2404 4.5005
R19287 VSS.n2725 VSS.n2404 4.5005
R19288 VSS.n2793 VSS.n2404 4.5005
R19289 VSS.n2859 VSS.n2404 4.5005
R19290 VSS.n3051 VSS.n2428 4.5005
R19291 VSS.n2428 VSS.n2351 4.5005
R19292 VSS.n2483 VSS.n2428 4.5005
R19293 VSS.n2484 VSS.n2428 4.5005
R19294 VSS.n2486 VSS.n2428 4.5005
R19295 VSS.n2489 VSS.n2428 4.5005
R19296 VSS.n2491 VSS.n2428 4.5005
R19297 VSS.n2492 VSS.n2428 4.5005
R19298 VSS.n2494 VSS.n2428 4.5005
R19299 VSS.n2497 VSS.n2428 4.5005
R19300 VSS.n2499 VSS.n2428 4.5005
R19301 VSS.n2500 VSS.n2428 4.5005
R19302 VSS.n2502 VSS.n2428 4.5005
R19303 VSS.n2505 VSS.n2428 4.5005
R19304 VSS.n2507 VSS.n2428 4.5005
R19305 VSS.n2508 VSS.n2428 4.5005
R19306 VSS.n2510 VSS.n2428 4.5005
R19307 VSS.n2513 VSS.n2428 4.5005
R19308 VSS.n2515 VSS.n2428 4.5005
R19309 VSS.n2516 VSS.n2428 4.5005
R19310 VSS.n2518 VSS.n2428 4.5005
R19311 VSS.n2521 VSS.n2428 4.5005
R19312 VSS.n2523 VSS.n2428 4.5005
R19313 VSS.n2524 VSS.n2428 4.5005
R19314 VSS.n2526 VSS.n2428 4.5005
R19315 VSS.n2529 VSS.n2428 4.5005
R19316 VSS.n2531 VSS.n2428 4.5005
R19317 VSS.n2532 VSS.n2428 4.5005
R19318 VSS.n2534 VSS.n2428 4.5005
R19319 VSS.n2537 VSS.n2428 4.5005
R19320 VSS.n2539 VSS.n2428 4.5005
R19321 VSS.n2540 VSS.n2428 4.5005
R19322 VSS.n2542 VSS.n2428 4.5005
R19323 VSS.n2545 VSS.n2428 4.5005
R19324 VSS.n2547 VSS.n2428 4.5005
R19325 VSS.n2548 VSS.n2428 4.5005
R19326 VSS.n2550 VSS.n2428 4.5005
R19327 VSS.n2553 VSS.n2428 4.5005
R19328 VSS.n2555 VSS.n2428 4.5005
R19329 VSS.n2556 VSS.n2428 4.5005
R19330 VSS.n2558 VSS.n2428 4.5005
R19331 VSS.n2561 VSS.n2428 4.5005
R19332 VSS.n2563 VSS.n2428 4.5005
R19333 VSS.n2564 VSS.n2428 4.5005
R19334 VSS.n2566 VSS.n2428 4.5005
R19335 VSS.n2569 VSS.n2428 4.5005
R19336 VSS.n2571 VSS.n2428 4.5005
R19337 VSS.n2572 VSS.n2428 4.5005
R19338 VSS.n2574 VSS.n2428 4.5005
R19339 VSS.n2577 VSS.n2428 4.5005
R19340 VSS.n2579 VSS.n2428 4.5005
R19341 VSS.n2580 VSS.n2428 4.5005
R19342 VSS.n2582 VSS.n2428 4.5005
R19343 VSS.n2585 VSS.n2428 4.5005
R19344 VSS.n2587 VSS.n2428 4.5005
R19345 VSS.n2588 VSS.n2428 4.5005
R19346 VSS.n2590 VSS.n2428 4.5005
R19347 VSS.n2593 VSS.n2428 4.5005
R19348 VSS.n2595 VSS.n2428 4.5005
R19349 VSS.n2596 VSS.n2428 4.5005
R19350 VSS.n2598 VSS.n2428 4.5005
R19351 VSS.n2601 VSS.n2428 4.5005
R19352 VSS.n2603 VSS.n2428 4.5005
R19353 VSS.n2604 VSS.n2428 4.5005
R19354 VSS.n2606 VSS.n2428 4.5005
R19355 VSS.n2609 VSS.n2428 4.5005
R19356 VSS.n2611 VSS.n2428 4.5005
R19357 VSS.n2612 VSS.n2428 4.5005
R19358 VSS.n2614 VSS.n2428 4.5005
R19359 VSS.n2617 VSS.n2428 4.5005
R19360 VSS.n2619 VSS.n2428 4.5005
R19361 VSS.n2620 VSS.n2428 4.5005
R19362 VSS.n2622 VSS.n2428 4.5005
R19363 VSS.n2625 VSS.n2428 4.5005
R19364 VSS.n2627 VSS.n2428 4.5005
R19365 VSS.n2628 VSS.n2428 4.5005
R19366 VSS.n2630 VSS.n2428 4.5005
R19367 VSS.n2633 VSS.n2428 4.5005
R19368 VSS.n2635 VSS.n2428 4.5005
R19369 VSS.n2636 VSS.n2428 4.5005
R19370 VSS.n2638 VSS.n2428 4.5005
R19371 VSS.n2640 VSS.n2428 4.5005
R19372 VSS.n2642 VSS.n2428 4.5005
R19373 VSS.n2643 VSS.n2428 4.5005
R19374 VSS.n2645 VSS.n2428 4.5005
R19375 VSS.n2648 VSS.n2428 4.5005
R19376 VSS.n2650 VSS.n2428 4.5005
R19377 VSS.n2651 VSS.n2428 4.5005
R19378 VSS.n2653 VSS.n2428 4.5005
R19379 VSS.n2656 VSS.n2428 4.5005
R19380 VSS.n2658 VSS.n2428 4.5005
R19381 VSS.n2659 VSS.n2428 4.5005
R19382 VSS.n2661 VSS.n2428 4.5005
R19383 VSS.n2664 VSS.n2428 4.5005
R19384 VSS.n2666 VSS.n2428 4.5005
R19385 VSS.n2667 VSS.n2428 4.5005
R19386 VSS.n2669 VSS.n2428 4.5005
R19387 VSS.n2672 VSS.n2428 4.5005
R19388 VSS.n2674 VSS.n2428 4.5005
R19389 VSS.n2675 VSS.n2428 4.5005
R19390 VSS.n2677 VSS.n2428 4.5005
R19391 VSS.n2680 VSS.n2428 4.5005
R19392 VSS.n2682 VSS.n2428 4.5005
R19393 VSS.n2683 VSS.n2428 4.5005
R19394 VSS.n2685 VSS.n2428 4.5005
R19395 VSS.n2688 VSS.n2428 4.5005
R19396 VSS.n2690 VSS.n2428 4.5005
R19397 VSS.n2691 VSS.n2428 4.5005
R19398 VSS.n2693 VSS.n2428 4.5005
R19399 VSS.n2696 VSS.n2428 4.5005
R19400 VSS.n2698 VSS.n2428 4.5005
R19401 VSS.n2699 VSS.n2428 4.5005
R19402 VSS.n2701 VSS.n2428 4.5005
R19403 VSS.n2704 VSS.n2428 4.5005
R19404 VSS.n2706 VSS.n2428 4.5005
R19405 VSS.n2707 VSS.n2428 4.5005
R19406 VSS.n2709 VSS.n2428 4.5005
R19407 VSS.n2712 VSS.n2428 4.5005
R19408 VSS.n2714 VSS.n2428 4.5005
R19409 VSS.n2715 VSS.n2428 4.5005
R19410 VSS.n2717 VSS.n2428 4.5005
R19411 VSS.n2720 VSS.n2428 4.5005
R19412 VSS.n2722 VSS.n2428 4.5005
R19413 VSS.n2723 VSS.n2428 4.5005
R19414 VSS.n2725 VSS.n2428 4.5005
R19415 VSS.n2793 VSS.n2428 4.5005
R19416 VSS.n2859 VSS.n2428 4.5005
R19417 VSS.n3051 VSS.n2403 4.5005
R19418 VSS.n2403 VSS.n2351 4.5005
R19419 VSS.n2483 VSS.n2403 4.5005
R19420 VSS.n2484 VSS.n2403 4.5005
R19421 VSS.n2486 VSS.n2403 4.5005
R19422 VSS.n2489 VSS.n2403 4.5005
R19423 VSS.n2491 VSS.n2403 4.5005
R19424 VSS.n2492 VSS.n2403 4.5005
R19425 VSS.n2494 VSS.n2403 4.5005
R19426 VSS.n2497 VSS.n2403 4.5005
R19427 VSS.n2499 VSS.n2403 4.5005
R19428 VSS.n2500 VSS.n2403 4.5005
R19429 VSS.n2502 VSS.n2403 4.5005
R19430 VSS.n2505 VSS.n2403 4.5005
R19431 VSS.n2507 VSS.n2403 4.5005
R19432 VSS.n2508 VSS.n2403 4.5005
R19433 VSS.n2510 VSS.n2403 4.5005
R19434 VSS.n2513 VSS.n2403 4.5005
R19435 VSS.n2515 VSS.n2403 4.5005
R19436 VSS.n2516 VSS.n2403 4.5005
R19437 VSS.n2518 VSS.n2403 4.5005
R19438 VSS.n2521 VSS.n2403 4.5005
R19439 VSS.n2523 VSS.n2403 4.5005
R19440 VSS.n2524 VSS.n2403 4.5005
R19441 VSS.n2526 VSS.n2403 4.5005
R19442 VSS.n2529 VSS.n2403 4.5005
R19443 VSS.n2531 VSS.n2403 4.5005
R19444 VSS.n2532 VSS.n2403 4.5005
R19445 VSS.n2534 VSS.n2403 4.5005
R19446 VSS.n2537 VSS.n2403 4.5005
R19447 VSS.n2539 VSS.n2403 4.5005
R19448 VSS.n2540 VSS.n2403 4.5005
R19449 VSS.n2542 VSS.n2403 4.5005
R19450 VSS.n2545 VSS.n2403 4.5005
R19451 VSS.n2547 VSS.n2403 4.5005
R19452 VSS.n2548 VSS.n2403 4.5005
R19453 VSS.n2550 VSS.n2403 4.5005
R19454 VSS.n2553 VSS.n2403 4.5005
R19455 VSS.n2555 VSS.n2403 4.5005
R19456 VSS.n2556 VSS.n2403 4.5005
R19457 VSS.n2558 VSS.n2403 4.5005
R19458 VSS.n2561 VSS.n2403 4.5005
R19459 VSS.n2563 VSS.n2403 4.5005
R19460 VSS.n2564 VSS.n2403 4.5005
R19461 VSS.n2566 VSS.n2403 4.5005
R19462 VSS.n2569 VSS.n2403 4.5005
R19463 VSS.n2571 VSS.n2403 4.5005
R19464 VSS.n2572 VSS.n2403 4.5005
R19465 VSS.n2574 VSS.n2403 4.5005
R19466 VSS.n2577 VSS.n2403 4.5005
R19467 VSS.n2579 VSS.n2403 4.5005
R19468 VSS.n2580 VSS.n2403 4.5005
R19469 VSS.n2582 VSS.n2403 4.5005
R19470 VSS.n2585 VSS.n2403 4.5005
R19471 VSS.n2587 VSS.n2403 4.5005
R19472 VSS.n2588 VSS.n2403 4.5005
R19473 VSS.n2590 VSS.n2403 4.5005
R19474 VSS.n2593 VSS.n2403 4.5005
R19475 VSS.n2595 VSS.n2403 4.5005
R19476 VSS.n2596 VSS.n2403 4.5005
R19477 VSS.n2598 VSS.n2403 4.5005
R19478 VSS.n2601 VSS.n2403 4.5005
R19479 VSS.n2603 VSS.n2403 4.5005
R19480 VSS.n2604 VSS.n2403 4.5005
R19481 VSS.n2606 VSS.n2403 4.5005
R19482 VSS.n2609 VSS.n2403 4.5005
R19483 VSS.n2611 VSS.n2403 4.5005
R19484 VSS.n2612 VSS.n2403 4.5005
R19485 VSS.n2614 VSS.n2403 4.5005
R19486 VSS.n2617 VSS.n2403 4.5005
R19487 VSS.n2619 VSS.n2403 4.5005
R19488 VSS.n2620 VSS.n2403 4.5005
R19489 VSS.n2622 VSS.n2403 4.5005
R19490 VSS.n2625 VSS.n2403 4.5005
R19491 VSS.n2627 VSS.n2403 4.5005
R19492 VSS.n2628 VSS.n2403 4.5005
R19493 VSS.n2630 VSS.n2403 4.5005
R19494 VSS.n2633 VSS.n2403 4.5005
R19495 VSS.n2635 VSS.n2403 4.5005
R19496 VSS.n2636 VSS.n2403 4.5005
R19497 VSS.n2638 VSS.n2403 4.5005
R19498 VSS.n2640 VSS.n2403 4.5005
R19499 VSS.n2642 VSS.n2403 4.5005
R19500 VSS.n2643 VSS.n2403 4.5005
R19501 VSS.n2645 VSS.n2403 4.5005
R19502 VSS.n2648 VSS.n2403 4.5005
R19503 VSS.n2650 VSS.n2403 4.5005
R19504 VSS.n2651 VSS.n2403 4.5005
R19505 VSS.n2653 VSS.n2403 4.5005
R19506 VSS.n2656 VSS.n2403 4.5005
R19507 VSS.n2658 VSS.n2403 4.5005
R19508 VSS.n2659 VSS.n2403 4.5005
R19509 VSS.n2661 VSS.n2403 4.5005
R19510 VSS.n2664 VSS.n2403 4.5005
R19511 VSS.n2666 VSS.n2403 4.5005
R19512 VSS.n2667 VSS.n2403 4.5005
R19513 VSS.n2669 VSS.n2403 4.5005
R19514 VSS.n2672 VSS.n2403 4.5005
R19515 VSS.n2674 VSS.n2403 4.5005
R19516 VSS.n2675 VSS.n2403 4.5005
R19517 VSS.n2677 VSS.n2403 4.5005
R19518 VSS.n2680 VSS.n2403 4.5005
R19519 VSS.n2682 VSS.n2403 4.5005
R19520 VSS.n2683 VSS.n2403 4.5005
R19521 VSS.n2685 VSS.n2403 4.5005
R19522 VSS.n2688 VSS.n2403 4.5005
R19523 VSS.n2690 VSS.n2403 4.5005
R19524 VSS.n2691 VSS.n2403 4.5005
R19525 VSS.n2693 VSS.n2403 4.5005
R19526 VSS.n2696 VSS.n2403 4.5005
R19527 VSS.n2698 VSS.n2403 4.5005
R19528 VSS.n2699 VSS.n2403 4.5005
R19529 VSS.n2701 VSS.n2403 4.5005
R19530 VSS.n2704 VSS.n2403 4.5005
R19531 VSS.n2706 VSS.n2403 4.5005
R19532 VSS.n2707 VSS.n2403 4.5005
R19533 VSS.n2709 VSS.n2403 4.5005
R19534 VSS.n2712 VSS.n2403 4.5005
R19535 VSS.n2714 VSS.n2403 4.5005
R19536 VSS.n2715 VSS.n2403 4.5005
R19537 VSS.n2717 VSS.n2403 4.5005
R19538 VSS.n2720 VSS.n2403 4.5005
R19539 VSS.n2722 VSS.n2403 4.5005
R19540 VSS.n2723 VSS.n2403 4.5005
R19541 VSS.n2725 VSS.n2403 4.5005
R19542 VSS.n2793 VSS.n2403 4.5005
R19543 VSS.n2859 VSS.n2403 4.5005
R19544 VSS.n3051 VSS.n2429 4.5005
R19545 VSS.n2429 VSS.n2351 4.5005
R19546 VSS.n2483 VSS.n2429 4.5005
R19547 VSS.n2484 VSS.n2429 4.5005
R19548 VSS.n2486 VSS.n2429 4.5005
R19549 VSS.n2489 VSS.n2429 4.5005
R19550 VSS.n2491 VSS.n2429 4.5005
R19551 VSS.n2492 VSS.n2429 4.5005
R19552 VSS.n2494 VSS.n2429 4.5005
R19553 VSS.n2497 VSS.n2429 4.5005
R19554 VSS.n2499 VSS.n2429 4.5005
R19555 VSS.n2500 VSS.n2429 4.5005
R19556 VSS.n2502 VSS.n2429 4.5005
R19557 VSS.n2505 VSS.n2429 4.5005
R19558 VSS.n2507 VSS.n2429 4.5005
R19559 VSS.n2508 VSS.n2429 4.5005
R19560 VSS.n2510 VSS.n2429 4.5005
R19561 VSS.n2513 VSS.n2429 4.5005
R19562 VSS.n2515 VSS.n2429 4.5005
R19563 VSS.n2516 VSS.n2429 4.5005
R19564 VSS.n2518 VSS.n2429 4.5005
R19565 VSS.n2521 VSS.n2429 4.5005
R19566 VSS.n2523 VSS.n2429 4.5005
R19567 VSS.n2524 VSS.n2429 4.5005
R19568 VSS.n2526 VSS.n2429 4.5005
R19569 VSS.n2529 VSS.n2429 4.5005
R19570 VSS.n2531 VSS.n2429 4.5005
R19571 VSS.n2532 VSS.n2429 4.5005
R19572 VSS.n2534 VSS.n2429 4.5005
R19573 VSS.n2537 VSS.n2429 4.5005
R19574 VSS.n2539 VSS.n2429 4.5005
R19575 VSS.n2540 VSS.n2429 4.5005
R19576 VSS.n2542 VSS.n2429 4.5005
R19577 VSS.n2545 VSS.n2429 4.5005
R19578 VSS.n2547 VSS.n2429 4.5005
R19579 VSS.n2548 VSS.n2429 4.5005
R19580 VSS.n2550 VSS.n2429 4.5005
R19581 VSS.n2553 VSS.n2429 4.5005
R19582 VSS.n2555 VSS.n2429 4.5005
R19583 VSS.n2556 VSS.n2429 4.5005
R19584 VSS.n2558 VSS.n2429 4.5005
R19585 VSS.n2561 VSS.n2429 4.5005
R19586 VSS.n2563 VSS.n2429 4.5005
R19587 VSS.n2564 VSS.n2429 4.5005
R19588 VSS.n2566 VSS.n2429 4.5005
R19589 VSS.n2569 VSS.n2429 4.5005
R19590 VSS.n2571 VSS.n2429 4.5005
R19591 VSS.n2572 VSS.n2429 4.5005
R19592 VSS.n2574 VSS.n2429 4.5005
R19593 VSS.n2577 VSS.n2429 4.5005
R19594 VSS.n2579 VSS.n2429 4.5005
R19595 VSS.n2580 VSS.n2429 4.5005
R19596 VSS.n2582 VSS.n2429 4.5005
R19597 VSS.n2585 VSS.n2429 4.5005
R19598 VSS.n2587 VSS.n2429 4.5005
R19599 VSS.n2588 VSS.n2429 4.5005
R19600 VSS.n2590 VSS.n2429 4.5005
R19601 VSS.n2593 VSS.n2429 4.5005
R19602 VSS.n2595 VSS.n2429 4.5005
R19603 VSS.n2596 VSS.n2429 4.5005
R19604 VSS.n2598 VSS.n2429 4.5005
R19605 VSS.n2601 VSS.n2429 4.5005
R19606 VSS.n2603 VSS.n2429 4.5005
R19607 VSS.n2604 VSS.n2429 4.5005
R19608 VSS.n2606 VSS.n2429 4.5005
R19609 VSS.n2609 VSS.n2429 4.5005
R19610 VSS.n2611 VSS.n2429 4.5005
R19611 VSS.n2612 VSS.n2429 4.5005
R19612 VSS.n2614 VSS.n2429 4.5005
R19613 VSS.n2617 VSS.n2429 4.5005
R19614 VSS.n2619 VSS.n2429 4.5005
R19615 VSS.n2620 VSS.n2429 4.5005
R19616 VSS.n2622 VSS.n2429 4.5005
R19617 VSS.n2625 VSS.n2429 4.5005
R19618 VSS.n2627 VSS.n2429 4.5005
R19619 VSS.n2628 VSS.n2429 4.5005
R19620 VSS.n2630 VSS.n2429 4.5005
R19621 VSS.n2633 VSS.n2429 4.5005
R19622 VSS.n2635 VSS.n2429 4.5005
R19623 VSS.n2636 VSS.n2429 4.5005
R19624 VSS.n2638 VSS.n2429 4.5005
R19625 VSS.n2640 VSS.n2429 4.5005
R19626 VSS.n2642 VSS.n2429 4.5005
R19627 VSS.n2643 VSS.n2429 4.5005
R19628 VSS.n2645 VSS.n2429 4.5005
R19629 VSS.n2648 VSS.n2429 4.5005
R19630 VSS.n2650 VSS.n2429 4.5005
R19631 VSS.n2651 VSS.n2429 4.5005
R19632 VSS.n2653 VSS.n2429 4.5005
R19633 VSS.n2656 VSS.n2429 4.5005
R19634 VSS.n2658 VSS.n2429 4.5005
R19635 VSS.n2659 VSS.n2429 4.5005
R19636 VSS.n2661 VSS.n2429 4.5005
R19637 VSS.n2664 VSS.n2429 4.5005
R19638 VSS.n2666 VSS.n2429 4.5005
R19639 VSS.n2667 VSS.n2429 4.5005
R19640 VSS.n2669 VSS.n2429 4.5005
R19641 VSS.n2672 VSS.n2429 4.5005
R19642 VSS.n2674 VSS.n2429 4.5005
R19643 VSS.n2675 VSS.n2429 4.5005
R19644 VSS.n2677 VSS.n2429 4.5005
R19645 VSS.n2680 VSS.n2429 4.5005
R19646 VSS.n2682 VSS.n2429 4.5005
R19647 VSS.n2683 VSS.n2429 4.5005
R19648 VSS.n2685 VSS.n2429 4.5005
R19649 VSS.n2688 VSS.n2429 4.5005
R19650 VSS.n2690 VSS.n2429 4.5005
R19651 VSS.n2691 VSS.n2429 4.5005
R19652 VSS.n2693 VSS.n2429 4.5005
R19653 VSS.n2696 VSS.n2429 4.5005
R19654 VSS.n2698 VSS.n2429 4.5005
R19655 VSS.n2699 VSS.n2429 4.5005
R19656 VSS.n2701 VSS.n2429 4.5005
R19657 VSS.n2704 VSS.n2429 4.5005
R19658 VSS.n2706 VSS.n2429 4.5005
R19659 VSS.n2707 VSS.n2429 4.5005
R19660 VSS.n2709 VSS.n2429 4.5005
R19661 VSS.n2712 VSS.n2429 4.5005
R19662 VSS.n2714 VSS.n2429 4.5005
R19663 VSS.n2715 VSS.n2429 4.5005
R19664 VSS.n2717 VSS.n2429 4.5005
R19665 VSS.n2720 VSS.n2429 4.5005
R19666 VSS.n2722 VSS.n2429 4.5005
R19667 VSS.n2723 VSS.n2429 4.5005
R19668 VSS.n2725 VSS.n2429 4.5005
R19669 VSS.n2793 VSS.n2429 4.5005
R19670 VSS.n2859 VSS.n2429 4.5005
R19671 VSS.n3051 VSS.n2402 4.5005
R19672 VSS.n2402 VSS.n2351 4.5005
R19673 VSS.n2483 VSS.n2402 4.5005
R19674 VSS.n2484 VSS.n2402 4.5005
R19675 VSS.n2486 VSS.n2402 4.5005
R19676 VSS.n2489 VSS.n2402 4.5005
R19677 VSS.n2491 VSS.n2402 4.5005
R19678 VSS.n2492 VSS.n2402 4.5005
R19679 VSS.n2494 VSS.n2402 4.5005
R19680 VSS.n2497 VSS.n2402 4.5005
R19681 VSS.n2499 VSS.n2402 4.5005
R19682 VSS.n2500 VSS.n2402 4.5005
R19683 VSS.n2502 VSS.n2402 4.5005
R19684 VSS.n2505 VSS.n2402 4.5005
R19685 VSS.n2507 VSS.n2402 4.5005
R19686 VSS.n2508 VSS.n2402 4.5005
R19687 VSS.n2510 VSS.n2402 4.5005
R19688 VSS.n2513 VSS.n2402 4.5005
R19689 VSS.n2515 VSS.n2402 4.5005
R19690 VSS.n2516 VSS.n2402 4.5005
R19691 VSS.n2518 VSS.n2402 4.5005
R19692 VSS.n2521 VSS.n2402 4.5005
R19693 VSS.n2523 VSS.n2402 4.5005
R19694 VSS.n2524 VSS.n2402 4.5005
R19695 VSS.n2526 VSS.n2402 4.5005
R19696 VSS.n2529 VSS.n2402 4.5005
R19697 VSS.n2531 VSS.n2402 4.5005
R19698 VSS.n2532 VSS.n2402 4.5005
R19699 VSS.n2534 VSS.n2402 4.5005
R19700 VSS.n2537 VSS.n2402 4.5005
R19701 VSS.n2539 VSS.n2402 4.5005
R19702 VSS.n2540 VSS.n2402 4.5005
R19703 VSS.n2542 VSS.n2402 4.5005
R19704 VSS.n2545 VSS.n2402 4.5005
R19705 VSS.n2547 VSS.n2402 4.5005
R19706 VSS.n2548 VSS.n2402 4.5005
R19707 VSS.n2550 VSS.n2402 4.5005
R19708 VSS.n2553 VSS.n2402 4.5005
R19709 VSS.n2555 VSS.n2402 4.5005
R19710 VSS.n2556 VSS.n2402 4.5005
R19711 VSS.n2558 VSS.n2402 4.5005
R19712 VSS.n2561 VSS.n2402 4.5005
R19713 VSS.n2563 VSS.n2402 4.5005
R19714 VSS.n2564 VSS.n2402 4.5005
R19715 VSS.n2566 VSS.n2402 4.5005
R19716 VSS.n2569 VSS.n2402 4.5005
R19717 VSS.n2571 VSS.n2402 4.5005
R19718 VSS.n2572 VSS.n2402 4.5005
R19719 VSS.n2574 VSS.n2402 4.5005
R19720 VSS.n2577 VSS.n2402 4.5005
R19721 VSS.n2579 VSS.n2402 4.5005
R19722 VSS.n2580 VSS.n2402 4.5005
R19723 VSS.n2582 VSS.n2402 4.5005
R19724 VSS.n2585 VSS.n2402 4.5005
R19725 VSS.n2587 VSS.n2402 4.5005
R19726 VSS.n2588 VSS.n2402 4.5005
R19727 VSS.n2590 VSS.n2402 4.5005
R19728 VSS.n2593 VSS.n2402 4.5005
R19729 VSS.n2595 VSS.n2402 4.5005
R19730 VSS.n2596 VSS.n2402 4.5005
R19731 VSS.n2598 VSS.n2402 4.5005
R19732 VSS.n2601 VSS.n2402 4.5005
R19733 VSS.n2603 VSS.n2402 4.5005
R19734 VSS.n2604 VSS.n2402 4.5005
R19735 VSS.n2606 VSS.n2402 4.5005
R19736 VSS.n2609 VSS.n2402 4.5005
R19737 VSS.n2611 VSS.n2402 4.5005
R19738 VSS.n2612 VSS.n2402 4.5005
R19739 VSS.n2614 VSS.n2402 4.5005
R19740 VSS.n2617 VSS.n2402 4.5005
R19741 VSS.n2619 VSS.n2402 4.5005
R19742 VSS.n2620 VSS.n2402 4.5005
R19743 VSS.n2622 VSS.n2402 4.5005
R19744 VSS.n2625 VSS.n2402 4.5005
R19745 VSS.n2627 VSS.n2402 4.5005
R19746 VSS.n2628 VSS.n2402 4.5005
R19747 VSS.n2630 VSS.n2402 4.5005
R19748 VSS.n2633 VSS.n2402 4.5005
R19749 VSS.n2635 VSS.n2402 4.5005
R19750 VSS.n2636 VSS.n2402 4.5005
R19751 VSS.n2638 VSS.n2402 4.5005
R19752 VSS.n2640 VSS.n2402 4.5005
R19753 VSS.n2642 VSS.n2402 4.5005
R19754 VSS.n2643 VSS.n2402 4.5005
R19755 VSS.n2645 VSS.n2402 4.5005
R19756 VSS.n2648 VSS.n2402 4.5005
R19757 VSS.n2650 VSS.n2402 4.5005
R19758 VSS.n2651 VSS.n2402 4.5005
R19759 VSS.n2653 VSS.n2402 4.5005
R19760 VSS.n2656 VSS.n2402 4.5005
R19761 VSS.n2658 VSS.n2402 4.5005
R19762 VSS.n2659 VSS.n2402 4.5005
R19763 VSS.n2661 VSS.n2402 4.5005
R19764 VSS.n2664 VSS.n2402 4.5005
R19765 VSS.n2666 VSS.n2402 4.5005
R19766 VSS.n2667 VSS.n2402 4.5005
R19767 VSS.n2669 VSS.n2402 4.5005
R19768 VSS.n2672 VSS.n2402 4.5005
R19769 VSS.n2674 VSS.n2402 4.5005
R19770 VSS.n2675 VSS.n2402 4.5005
R19771 VSS.n2677 VSS.n2402 4.5005
R19772 VSS.n2680 VSS.n2402 4.5005
R19773 VSS.n2682 VSS.n2402 4.5005
R19774 VSS.n2683 VSS.n2402 4.5005
R19775 VSS.n2685 VSS.n2402 4.5005
R19776 VSS.n2688 VSS.n2402 4.5005
R19777 VSS.n2690 VSS.n2402 4.5005
R19778 VSS.n2691 VSS.n2402 4.5005
R19779 VSS.n2693 VSS.n2402 4.5005
R19780 VSS.n2696 VSS.n2402 4.5005
R19781 VSS.n2698 VSS.n2402 4.5005
R19782 VSS.n2699 VSS.n2402 4.5005
R19783 VSS.n2701 VSS.n2402 4.5005
R19784 VSS.n2704 VSS.n2402 4.5005
R19785 VSS.n2706 VSS.n2402 4.5005
R19786 VSS.n2707 VSS.n2402 4.5005
R19787 VSS.n2709 VSS.n2402 4.5005
R19788 VSS.n2712 VSS.n2402 4.5005
R19789 VSS.n2714 VSS.n2402 4.5005
R19790 VSS.n2715 VSS.n2402 4.5005
R19791 VSS.n2717 VSS.n2402 4.5005
R19792 VSS.n2720 VSS.n2402 4.5005
R19793 VSS.n2722 VSS.n2402 4.5005
R19794 VSS.n2723 VSS.n2402 4.5005
R19795 VSS.n2725 VSS.n2402 4.5005
R19796 VSS.n2793 VSS.n2402 4.5005
R19797 VSS.n2859 VSS.n2402 4.5005
R19798 VSS.n3051 VSS.n2430 4.5005
R19799 VSS.n2430 VSS.n2351 4.5005
R19800 VSS.n2483 VSS.n2430 4.5005
R19801 VSS.n2484 VSS.n2430 4.5005
R19802 VSS.n2486 VSS.n2430 4.5005
R19803 VSS.n2489 VSS.n2430 4.5005
R19804 VSS.n2491 VSS.n2430 4.5005
R19805 VSS.n2492 VSS.n2430 4.5005
R19806 VSS.n2494 VSS.n2430 4.5005
R19807 VSS.n2497 VSS.n2430 4.5005
R19808 VSS.n2499 VSS.n2430 4.5005
R19809 VSS.n2500 VSS.n2430 4.5005
R19810 VSS.n2502 VSS.n2430 4.5005
R19811 VSS.n2505 VSS.n2430 4.5005
R19812 VSS.n2507 VSS.n2430 4.5005
R19813 VSS.n2508 VSS.n2430 4.5005
R19814 VSS.n2510 VSS.n2430 4.5005
R19815 VSS.n2513 VSS.n2430 4.5005
R19816 VSS.n2515 VSS.n2430 4.5005
R19817 VSS.n2516 VSS.n2430 4.5005
R19818 VSS.n2518 VSS.n2430 4.5005
R19819 VSS.n2521 VSS.n2430 4.5005
R19820 VSS.n2523 VSS.n2430 4.5005
R19821 VSS.n2524 VSS.n2430 4.5005
R19822 VSS.n2526 VSS.n2430 4.5005
R19823 VSS.n2529 VSS.n2430 4.5005
R19824 VSS.n2531 VSS.n2430 4.5005
R19825 VSS.n2532 VSS.n2430 4.5005
R19826 VSS.n2534 VSS.n2430 4.5005
R19827 VSS.n2537 VSS.n2430 4.5005
R19828 VSS.n2539 VSS.n2430 4.5005
R19829 VSS.n2540 VSS.n2430 4.5005
R19830 VSS.n2542 VSS.n2430 4.5005
R19831 VSS.n2545 VSS.n2430 4.5005
R19832 VSS.n2547 VSS.n2430 4.5005
R19833 VSS.n2548 VSS.n2430 4.5005
R19834 VSS.n2550 VSS.n2430 4.5005
R19835 VSS.n2553 VSS.n2430 4.5005
R19836 VSS.n2555 VSS.n2430 4.5005
R19837 VSS.n2556 VSS.n2430 4.5005
R19838 VSS.n2558 VSS.n2430 4.5005
R19839 VSS.n2561 VSS.n2430 4.5005
R19840 VSS.n2563 VSS.n2430 4.5005
R19841 VSS.n2564 VSS.n2430 4.5005
R19842 VSS.n2566 VSS.n2430 4.5005
R19843 VSS.n2569 VSS.n2430 4.5005
R19844 VSS.n2571 VSS.n2430 4.5005
R19845 VSS.n2572 VSS.n2430 4.5005
R19846 VSS.n2574 VSS.n2430 4.5005
R19847 VSS.n2577 VSS.n2430 4.5005
R19848 VSS.n2579 VSS.n2430 4.5005
R19849 VSS.n2580 VSS.n2430 4.5005
R19850 VSS.n2582 VSS.n2430 4.5005
R19851 VSS.n2585 VSS.n2430 4.5005
R19852 VSS.n2587 VSS.n2430 4.5005
R19853 VSS.n2588 VSS.n2430 4.5005
R19854 VSS.n2590 VSS.n2430 4.5005
R19855 VSS.n2593 VSS.n2430 4.5005
R19856 VSS.n2595 VSS.n2430 4.5005
R19857 VSS.n2596 VSS.n2430 4.5005
R19858 VSS.n2598 VSS.n2430 4.5005
R19859 VSS.n2601 VSS.n2430 4.5005
R19860 VSS.n2603 VSS.n2430 4.5005
R19861 VSS.n2604 VSS.n2430 4.5005
R19862 VSS.n2606 VSS.n2430 4.5005
R19863 VSS.n2609 VSS.n2430 4.5005
R19864 VSS.n2611 VSS.n2430 4.5005
R19865 VSS.n2612 VSS.n2430 4.5005
R19866 VSS.n2614 VSS.n2430 4.5005
R19867 VSS.n2617 VSS.n2430 4.5005
R19868 VSS.n2619 VSS.n2430 4.5005
R19869 VSS.n2620 VSS.n2430 4.5005
R19870 VSS.n2622 VSS.n2430 4.5005
R19871 VSS.n2625 VSS.n2430 4.5005
R19872 VSS.n2627 VSS.n2430 4.5005
R19873 VSS.n2628 VSS.n2430 4.5005
R19874 VSS.n2630 VSS.n2430 4.5005
R19875 VSS.n2633 VSS.n2430 4.5005
R19876 VSS.n2635 VSS.n2430 4.5005
R19877 VSS.n2636 VSS.n2430 4.5005
R19878 VSS.n2638 VSS.n2430 4.5005
R19879 VSS.n2640 VSS.n2430 4.5005
R19880 VSS.n2642 VSS.n2430 4.5005
R19881 VSS.n2643 VSS.n2430 4.5005
R19882 VSS.n2645 VSS.n2430 4.5005
R19883 VSS.n2648 VSS.n2430 4.5005
R19884 VSS.n2650 VSS.n2430 4.5005
R19885 VSS.n2651 VSS.n2430 4.5005
R19886 VSS.n2653 VSS.n2430 4.5005
R19887 VSS.n2656 VSS.n2430 4.5005
R19888 VSS.n2658 VSS.n2430 4.5005
R19889 VSS.n2659 VSS.n2430 4.5005
R19890 VSS.n2661 VSS.n2430 4.5005
R19891 VSS.n2664 VSS.n2430 4.5005
R19892 VSS.n2666 VSS.n2430 4.5005
R19893 VSS.n2667 VSS.n2430 4.5005
R19894 VSS.n2669 VSS.n2430 4.5005
R19895 VSS.n2672 VSS.n2430 4.5005
R19896 VSS.n2674 VSS.n2430 4.5005
R19897 VSS.n2675 VSS.n2430 4.5005
R19898 VSS.n2677 VSS.n2430 4.5005
R19899 VSS.n2680 VSS.n2430 4.5005
R19900 VSS.n2682 VSS.n2430 4.5005
R19901 VSS.n2683 VSS.n2430 4.5005
R19902 VSS.n2685 VSS.n2430 4.5005
R19903 VSS.n2688 VSS.n2430 4.5005
R19904 VSS.n2690 VSS.n2430 4.5005
R19905 VSS.n2691 VSS.n2430 4.5005
R19906 VSS.n2693 VSS.n2430 4.5005
R19907 VSS.n2696 VSS.n2430 4.5005
R19908 VSS.n2698 VSS.n2430 4.5005
R19909 VSS.n2699 VSS.n2430 4.5005
R19910 VSS.n2701 VSS.n2430 4.5005
R19911 VSS.n2704 VSS.n2430 4.5005
R19912 VSS.n2706 VSS.n2430 4.5005
R19913 VSS.n2707 VSS.n2430 4.5005
R19914 VSS.n2709 VSS.n2430 4.5005
R19915 VSS.n2712 VSS.n2430 4.5005
R19916 VSS.n2714 VSS.n2430 4.5005
R19917 VSS.n2715 VSS.n2430 4.5005
R19918 VSS.n2717 VSS.n2430 4.5005
R19919 VSS.n2720 VSS.n2430 4.5005
R19920 VSS.n2722 VSS.n2430 4.5005
R19921 VSS.n2723 VSS.n2430 4.5005
R19922 VSS.n2725 VSS.n2430 4.5005
R19923 VSS.n2793 VSS.n2430 4.5005
R19924 VSS.n2859 VSS.n2430 4.5005
R19925 VSS.n3051 VSS.n2401 4.5005
R19926 VSS.n2401 VSS.n2351 4.5005
R19927 VSS.n2483 VSS.n2401 4.5005
R19928 VSS.n2484 VSS.n2401 4.5005
R19929 VSS.n2486 VSS.n2401 4.5005
R19930 VSS.n2489 VSS.n2401 4.5005
R19931 VSS.n2491 VSS.n2401 4.5005
R19932 VSS.n2492 VSS.n2401 4.5005
R19933 VSS.n2494 VSS.n2401 4.5005
R19934 VSS.n2497 VSS.n2401 4.5005
R19935 VSS.n2499 VSS.n2401 4.5005
R19936 VSS.n2500 VSS.n2401 4.5005
R19937 VSS.n2502 VSS.n2401 4.5005
R19938 VSS.n2505 VSS.n2401 4.5005
R19939 VSS.n2507 VSS.n2401 4.5005
R19940 VSS.n2508 VSS.n2401 4.5005
R19941 VSS.n2510 VSS.n2401 4.5005
R19942 VSS.n2513 VSS.n2401 4.5005
R19943 VSS.n2515 VSS.n2401 4.5005
R19944 VSS.n2516 VSS.n2401 4.5005
R19945 VSS.n2518 VSS.n2401 4.5005
R19946 VSS.n2521 VSS.n2401 4.5005
R19947 VSS.n2523 VSS.n2401 4.5005
R19948 VSS.n2524 VSS.n2401 4.5005
R19949 VSS.n2526 VSS.n2401 4.5005
R19950 VSS.n2529 VSS.n2401 4.5005
R19951 VSS.n2531 VSS.n2401 4.5005
R19952 VSS.n2532 VSS.n2401 4.5005
R19953 VSS.n2534 VSS.n2401 4.5005
R19954 VSS.n2537 VSS.n2401 4.5005
R19955 VSS.n2539 VSS.n2401 4.5005
R19956 VSS.n2540 VSS.n2401 4.5005
R19957 VSS.n2542 VSS.n2401 4.5005
R19958 VSS.n2545 VSS.n2401 4.5005
R19959 VSS.n2547 VSS.n2401 4.5005
R19960 VSS.n2548 VSS.n2401 4.5005
R19961 VSS.n2550 VSS.n2401 4.5005
R19962 VSS.n2553 VSS.n2401 4.5005
R19963 VSS.n2555 VSS.n2401 4.5005
R19964 VSS.n2556 VSS.n2401 4.5005
R19965 VSS.n2558 VSS.n2401 4.5005
R19966 VSS.n2561 VSS.n2401 4.5005
R19967 VSS.n2563 VSS.n2401 4.5005
R19968 VSS.n2564 VSS.n2401 4.5005
R19969 VSS.n2566 VSS.n2401 4.5005
R19970 VSS.n2569 VSS.n2401 4.5005
R19971 VSS.n2571 VSS.n2401 4.5005
R19972 VSS.n2572 VSS.n2401 4.5005
R19973 VSS.n2574 VSS.n2401 4.5005
R19974 VSS.n2577 VSS.n2401 4.5005
R19975 VSS.n2579 VSS.n2401 4.5005
R19976 VSS.n2580 VSS.n2401 4.5005
R19977 VSS.n2582 VSS.n2401 4.5005
R19978 VSS.n2585 VSS.n2401 4.5005
R19979 VSS.n2587 VSS.n2401 4.5005
R19980 VSS.n2588 VSS.n2401 4.5005
R19981 VSS.n2590 VSS.n2401 4.5005
R19982 VSS.n2593 VSS.n2401 4.5005
R19983 VSS.n2595 VSS.n2401 4.5005
R19984 VSS.n2596 VSS.n2401 4.5005
R19985 VSS.n2598 VSS.n2401 4.5005
R19986 VSS.n2601 VSS.n2401 4.5005
R19987 VSS.n2603 VSS.n2401 4.5005
R19988 VSS.n2604 VSS.n2401 4.5005
R19989 VSS.n2606 VSS.n2401 4.5005
R19990 VSS.n2609 VSS.n2401 4.5005
R19991 VSS.n2611 VSS.n2401 4.5005
R19992 VSS.n2612 VSS.n2401 4.5005
R19993 VSS.n2614 VSS.n2401 4.5005
R19994 VSS.n2617 VSS.n2401 4.5005
R19995 VSS.n2619 VSS.n2401 4.5005
R19996 VSS.n2620 VSS.n2401 4.5005
R19997 VSS.n2622 VSS.n2401 4.5005
R19998 VSS.n2625 VSS.n2401 4.5005
R19999 VSS.n2627 VSS.n2401 4.5005
R20000 VSS.n2628 VSS.n2401 4.5005
R20001 VSS.n2630 VSS.n2401 4.5005
R20002 VSS.n2633 VSS.n2401 4.5005
R20003 VSS.n2635 VSS.n2401 4.5005
R20004 VSS.n2636 VSS.n2401 4.5005
R20005 VSS.n2638 VSS.n2401 4.5005
R20006 VSS.n2640 VSS.n2401 4.5005
R20007 VSS.n2642 VSS.n2401 4.5005
R20008 VSS.n2643 VSS.n2401 4.5005
R20009 VSS.n2645 VSS.n2401 4.5005
R20010 VSS.n2648 VSS.n2401 4.5005
R20011 VSS.n2650 VSS.n2401 4.5005
R20012 VSS.n2651 VSS.n2401 4.5005
R20013 VSS.n2653 VSS.n2401 4.5005
R20014 VSS.n2656 VSS.n2401 4.5005
R20015 VSS.n2658 VSS.n2401 4.5005
R20016 VSS.n2659 VSS.n2401 4.5005
R20017 VSS.n2661 VSS.n2401 4.5005
R20018 VSS.n2664 VSS.n2401 4.5005
R20019 VSS.n2666 VSS.n2401 4.5005
R20020 VSS.n2667 VSS.n2401 4.5005
R20021 VSS.n2669 VSS.n2401 4.5005
R20022 VSS.n2672 VSS.n2401 4.5005
R20023 VSS.n2674 VSS.n2401 4.5005
R20024 VSS.n2675 VSS.n2401 4.5005
R20025 VSS.n2677 VSS.n2401 4.5005
R20026 VSS.n2680 VSS.n2401 4.5005
R20027 VSS.n2682 VSS.n2401 4.5005
R20028 VSS.n2683 VSS.n2401 4.5005
R20029 VSS.n2685 VSS.n2401 4.5005
R20030 VSS.n2688 VSS.n2401 4.5005
R20031 VSS.n2690 VSS.n2401 4.5005
R20032 VSS.n2691 VSS.n2401 4.5005
R20033 VSS.n2693 VSS.n2401 4.5005
R20034 VSS.n2696 VSS.n2401 4.5005
R20035 VSS.n2698 VSS.n2401 4.5005
R20036 VSS.n2699 VSS.n2401 4.5005
R20037 VSS.n2701 VSS.n2401 4.5005
R20038 VSS.n2704 VSS.n2401 4.5005
R20039 VSS.n2706 VSS.n2401 4.5005
R20040 VSS.n2707 VSS.n2401 4.5005
R20041 VSS.n2709 VSS.n2401 4.5005
R20042 VSS.n2712 VSS.n2401 4.5005
R20043 VSS.n2714 VSS.n2401 4.5005
R20044 VSS.n2715 VSS.n2401 4.5005
R20045 VSS.n2717 VSS.n2401 4.5005
R20046 VSS.n2720 VSS.n2401 4.5005
R20047 VSS.n2722 VSS.n2401 4.5005
R20048 VSS.n2723 VSS.n2401 4.5005
R20049 VSS.n2725 VSS.n2401 4.5005
R20050 VSS.n2793 VSS.n2401 4.5005
R20051 VSS.n2859 VSS.n2401 4.5005
R20052 VSS.n3051 VSS.n2431 4.5005
R20053 VSS.n2431 VSS.n2351 4.5005
R20054 VSS.n2483 VSS.n2431 4.5005
R20055 VSS.n2484 VSS.n2431 4.5005
R20056 VSS.n2486 VSS.n2431 4.5005
R20057 VSS.n2489 VSS.n2431 4.5005
R20058 VSS.n2491 VSS.n2431 4.5005
R20059 VSS.n2492 VSS.n2431 4.5005
R20060 VSS.n2494 VSS.n2431 4.5005
R20061 VSS.n2497 VSS.n2431 4.5005
R20062 VSS.n2499 VSS.n2431 4.5005
R20063 VSS.n2500 VSS.n2431 4.5005
R20064 VSS.n2502 VSS.n2431 4.5005
R20065 VSS.n2505 VSS.n2431 4.5005
R20066 VSS.n2507 VSS.n2431 4.5005
R20067 VSS.n2508 VSS.n2431 4.5005
R20068 VSS.n2510 VSS.n2431 4.5005
R20069 VSS.n2513 VSS.n2431 4.5005
R20070 VSS.n2515 VSS.n2431 4.5005
R20071 VSS.n2516 VSS.n2431 4.5005
R20072 VSS.n2518 VSS.n2431 4.5005
R20073 VSS.n2521 VSS.n2431 4.5005
R20074 VSS.n2523 VSS.n2431 4.5005
R20075 VSS.n2524 VSS.n2431 4.5005
R20076 VSS.n2526 VSS.n2431 4.5005
R20077 VSS.n2529 VSS.n2431 4.5005
R20078 VSS.n2531 VSS.n2431 4.5005
R20079 VSS.n2532 VSS.n2431 4.5005
R20080 VSS.n2534 VSS.n2431 4.5005
R20081 VSS.n2537 VSS.n2431 4.5005
R20082 VSS.n2539 VSS.n2431 4.5005
R20083 VSS.n2540 VSS.n2431 4.5005
R20084 VSS.n2542 VSS.n2431 4.5005
R20085 VSS.n2545 VSS.n2431 4.5005
R20086 VSS.n2547 VSS.n2431 4.5005
R20087 VSS.n2548 VSS.n2431 4.5005
R20088 VSS.n2550 VSS.n2431 4.5005
R20089 VSS.n2553 VSS.n2431 4.5005
R20090 VSS.n2555 VSS.n2431 4.5005
R20091 VSS.n2556 VSS.n2431 4.5005
R20092 VSS.n2558 VSS.n2431 4.5005
R20093 VSS.n2561 VSS.n2431 4.5005
R20094 VSS.n2563 VSS.n2431 4.5005
R20095 VSS.n2564 VSS.n2431 4.5005
R20096 VSS.n2566 VSS.n2431 4.5005
R20097 VSS.n2569 VSS.n2431 4.5005
R20098 VSS.n2571 VSS.n2431 4.5005
R20099 VSS.n2572 VSS.n2431 4.5005
R20100 VSS.n2574 VSS.n2431 4.5005
R20101 VSS.n2577 VSS.n2431 4.5005
R20102 VSS.n2579 VSS.n2431 4.5005
R20103 VSS.n2580 VSS.n2431 4.5005
R20104 VSS.n2582 VSS.n2431 4.5005
R20105 VSS.n2585 VSS.n2431 4.5005
R20106 VSS.n2587 VSS.n2431 4.5005
R20107 VSS.n2588 VSS.n2431 4.5005
R20108 VSS.n2590 VSS.n2431 4.5005
R20109 VSS.n2593 VSS.n2431 4.5005
R20110 VSS.n2595 VSS.n2431 4.5005
R20111 VSS.n2596 VSS.n2431 4.5005
R20112 VSS.n2598 VSS.n2431 4.5005
R20113 VSS.n2601 VSS.n2431 4.5005
R20114 VSS.n2603 VSS.n2431 4.5005
R20115 VSS.n2604 VSS.n2431 4.5005
R20116 VSS.n2606 VSS.n2431 4.5005
R20117 VSS.n2609 VSS.n2431 4.5005
R20118 VSS.n2611 VSS.n2431 4.5005
R20119 VSS.n2612 VSS.n2431 4.5005
R20120 VSS.n2614 VSS.n2431 4.5005
R20121 VSS.n2617 VSS.n2431 4.5005
R20122 VSS.n2619 VSS.n2431 4.5005
R20123 VSS.n2620 VSS.n2431 4.5005
R20124 VSS.n2622 VSS.n2431 4.5005
R20125 VSS.n2625 VSS.n2431 4.5005
R20126 VSS.n2627 VSS.n2431 4.5005
R20127 VSS.n2628 VSS.n2431 4.5005
R20128 VSS.n2630 VSS.n2431 4.5005
R20129 VSS.n2633 VSS.n2431 4.5005
R20130 VSS.n2635 VSS.n2431 4.5005
R20131 VSS.n2636 VSS.n2431 4.5005
R20132 VSS.n2638 VSS.n2431 4.5005
R20133 VSS.n2640 VSS.n2431 4.5005
R20134 VSS.n2642 VSS.n2431 4.5005
R20135 VSS.n2643 VSS.n2431 4.5005
R20136 VSS.n2645 VSS.n2431 4.5005
R20137 VSS.n2648 VSS.n2431 4.5005
R20138 VSS.n2650 VSS.n2431 4.5005
R20139 VSS.n2651 VSS.n2431 4.5005
R20140 VSS.n2653 VSS.n2431 4.5005
R20141 VSS.n2656 VSS.n2431 4.5005
R20142 VSS.n2658 VSS.n2431 4.5005
R20143 VSS.n2659 VSS.n2431 4.5005
R20144 VSS.n2661 VSS.n2431 4.5005
R20145 VSS.n2664 VSS.n2431 4.5005
R20146 VSS.n2666 VSS.n2431 4.5005
R20147 VSS.n2667 VSS.n2431 4.5005
R20148 VSS.n2669 VSS.n2431 4.5005
R20149 VSS.n2672 VSS.n2431 4.5005
R20150 VSS.n2674 VSS.n2431 4.5005
R20151 VSS.n2675 VSS.n2431 4.5005
R20152 VSS.n2677 VSS.n2431 4.5005
R20153 VSS.n2680 VSS.n2431 4.5005
R20154 VSS.n2682 VSS.n2431 4.5005
R20155 VSS.n2683 VSS.n2431 4.5005
R20156 VSS.n2685 VSS.n2431 4.5005
R20157 VSS.n2688 VSS.n2431 4.5005
R20158 VSS.n2690 VSS.n2431 4.5005
R20159 VSS.n2691 VSS.n2431 4.5005
R20160 VSS.n2693 VSS.n2431 4.5005
R20161 VSS.n2696 VSS.n2431 4.5005
R20162 VSS.n2698 VSS.n2431 4.5005
R20163 VSS.n2699 VSS.n2431 4.5005
R20164 VSS.n2701 VSS.n2431 4.5005
R20165 VSS.n2704 VSS.n2431 4.5005
R20166 VSS.n2706 VSS.n2431 4.5005
R20167 VSS.n2707 VSS.n2431 4.5005
R20168 VSS.n2709 VSS.n2431 4.5005
R20169 VSS.n2712 VSS.n2431 4.5005
R20170 VSS.n2714 VSS.n2431 4.5005
R20171 VSS.n2715 VSS.n2431 4.5005
R20172 VSS.n2717 VSS.n2431 4.5005
R20173 VSS.n2720 VSS.n2431 4.5005
R20174 VSS.n2722 VSS.n2431 4.5005
R20175 VSS.n2723 VSS.n2431 4.5005
R20176 VSS.n2725 VSS.n2431 4.5005
R20177 VSS.n2793 VSS.n2431 4.5005
R20178 VSS.n2859 VSS.n2431 4.5005
R20179 VSS.n3051 VSS.n2400 4.5005
R20180 VSS.n2400 VSS.n2351 4.5005
R20181 VSS.n2483 VSS.n2400 4.5005
R20182 VSS.n2484 VSS.n2400 4.5005
R20183 VSS.n2486 VSS.n2400 4.5005
R20184 VSS.n2489 VSS.n2400 4.5005
R20185 VSS.n2491 VSS.n2400 4.5005
R20186 VSS.n2492 VSS.n2400 4.5005
R20187 VSS.n2494 VSS.n2400 4.5005
R20188 VSS.n2497 VSS.n2400 4.5005
R20189 VSS.n2499 VSS.n2400 4.5005
R20190 VSS.n2500 VSS.n2400 4.5005
R20191 VSS.n2502 VSS.n2400 4.5005
R20192 VSS.n2505 VSS.n2400 4.5005
R20193 VSS.n2507 VSS.n2400 4.5005
R20194 VSS.n2508 VSS.n2400 4.5005
R20195 VSS.n2510 VSS.n2400 4.5005
R20196 VSS.n2513 VSS.n2400 4.5005
R20197 VSS.n2515 VSS.n2400 4.5005
R20198 VSS.n2516 VSS.n2400 4.5005
R20199 VSS.n2518 VSS.n2400 4.5005
R20200 VSS.n2521 VSS.n2400 4.5005
R20201 VSS.n2523 VSS.n2400 4.5005
R20202 VSS.n2524 VSS.n2400 4.5005
R20203 VSS.n2526 VSS.n2400 4.5005
R20204 VSS.n2529 VSS.n2400 4.5005
R20205 VSS.n2531 VSS.n2400 4.5005
R20206 VSS.n2532 VSS.n2400 4.5005
R20207 VSS.n2534 VSS.n2400 4.5005
R20208 VSS.n2537 VSS.n2400 4.5005
R20209 VSS.n2539 VSS.n2400 4.5005
R20210 VSS.n2540 VSS.n2400 4.5005
R20211 VSS.n2542 VSS.n2400 4.5005
R20212 VSS.n2545 VSS.n2400 4.5005
R20213 VSS.n2547 VSS.n2400 4.5005
R20214 VSS.n2548 VSS.n2400 4.5005
R20215 VSS.n2550 VSS.n2400 4.5005
R20216 VSS.n2553 VSS.n2400 4.5005
R20217 VSS.n2555 VSS.n2400 4.5005
R20218 VSS.n2556 VSS.n2400 4.5005
R20219 VSS.n2558 VSS.n2400 4.5005
R20220 VSS.n2561 VSS.n2400 4.5005
R20221 VSS.n2563 VSS.n2400 4.5005
R20222 VSS.n2564 VSS.n2400 4.5005
R20223 VSS.n2566 VSS.n2400 4.5005
R20224 VSS.n2569 VSS.n2400 4.5005
R20225 VSS.n2571 VSS.n2400 4.5005
R20226 VSS.n2572 VSS.n2400 4.5005
R20227 VSS.n2574 VSS.n2400 4.5005
R20228 VSS.n2577 VSS.n2400 4.5005
R20229 VSS.n2579 VSS.n2400 4.5005
R20230 VSS.n2580 VSS.n2400 4.5005
R20231 VSS.n2582 VSS.n2400 4.5005
R20232 VSS.n2585 VSS.n2400 4.5005
R20233 VSS.n2587 VSS.n2400 4.5005
R20234 VSS.n2588 VSS.n2400 4.5005
R20235 VSS.n2590 VSS.n2400 4.5005
R20236 VSS.n2593 VSS.n2400 4.5005
R20237 VSS.n2595 VSS.n2400 4.5005
R20238 VSS.n2596 VSS.n2400 4.5005
R20239 VSS.n2598 VSS.n2400 4.5005
R20240 VSS.n2601 VSS.n2400 4.5005
R20241 VSS.n2603 VSS.n2400 4.5005
R20242 VSS.n2604 VSS.n2400 4.5005
R20243 VSS.n2606 VSS.n2400 4.5005
R20244 VSS.n2609 VSS.n2400 4.5005
R20245 VSS.n2611 VSS.n2400 4.5005
R20246 VSS.n2612 VSS.n2400 4.5005
R20247 VSS.n2614 VSS.n2400 4.5005
R20248 VSS.n2617 VSS.n2400 4.5005
R20249 VSS.n2619 VSS.n2400 4.5005
R20250 VSS.n2620 VSS.n2400 4.5005
R20251 VSS.n2622 VSS.n2400 4.5005
R20252 VSS.n2625 VSS.n2400 4.5005
R20253 VSS.n2627 VSS.n2400 4.5005
R20254 VSS.n2628 VSS.n2400 4.5005
R20255 VSS.n2630 VSS.n2400 4.5005
R20256 VSS.n2633 VSS.n2400 4.5005
R20257 VSS.n2635 VSS.n2400 4.5005
R20258 VSS.n2636 VSS.n2400 4.5005
R20259 VSS.n2638 VSS.n2400 4.5005
R20260 VSS.n2640 VSS.n2400 4.5005
R20261 VSS.n2642 VSS.n2400 4.5005
R20262 VSS.n2643 VSS.n2400 4.5005
R20263 VSS.n2645 VSS.n2400 4.5005
R20264 VSS.n2648 VSS.n2400 4.5005
R20265 VSS.n2650 VSS.n2400 4.5005
R20266 VSS.n2651 VSS.n2400 4.5005
R20267 VSS.n2653 VSS.n2400 4.5005
R20268 VSS.n2656 VSS.n2400 4.5005
R20269 VSS.n2658 VSS.n2400 4.5005
R20270 VSS.n2659 VSS.n2400 4.5005
R20271 VSS.n2661 VSS.n2400 4.5005
R20272 VSS.n2664 VSS.n2400 4.5005
R20273 VSS.n2666 VSS.n2400 4.5005
R20274 VSS.n2667 VSS.n2400 4.5005
R20275 VSS.n2669 VSS.n2400 4.5005
R20276 VSS.n2672 VSS.n2400 4.5005
R20277 VSS.n2674 VSS.n2400 4.5005
R20278 VSS.n2675 VSS.n2400 4.5005
R20279 VSS.n2677 VSS.n2400 4.5005
R20280 VSS.n2680 VSS.n2400 4.5005
R20281 VSS.n2682 VSS.n2400 4.5005
R20282 VSS.n2683 VSS.n2400 4.5005
R20283 VSS.n2685 VSS.n2400 4.5005
R20284 VSS.n2688 VSS.n2400 4.5005
R20285 VSS.n2690 VSS.n2400 4.5005
R20286 VSS.n2691 VSS.n2400 4.5005
R20287 VSS.n2693 VSS.n2400 4.5005
R20288 VSS.n2696 VSS.n2400 4.5005
R20289 VSS.n2698 VSS.n2400 4.5005
R20290 VSS.n2699 VSS.n2400 4.5005
R20291 VSS.n2701 VSS.n2400 4.5005
R20292 VSS.n2704 VSS.n2400 4.5005
R20293 VSS.n2706 VSS.n2400 4.5005
R20294 VSS.n2707 VSS.n2400 4.5005
R20295 VSS.n2709 VSS.n2400 4.5005
R20296 VSS.n2712 VSS.n2400 4.5005
R20297 VSS.n2714 VSS.n2400 4.5005
R20298 VSS.n2715 VSS.n2400 4.5005
R20299 VSS.n2717 VSS.n2400 4.5005
R20300 VSS.n2720 VSS.n2400 4.5005
R20301 VSS.n2722 VSS.n2400 4.5005
R20302 VSS.n2723 VSS.n2400 4.5005
R20303 VSS.n2725 VSS.n2400 4.5005
R20304 VSS.n2793 VSS.n2400 4.5005
R20305 VSS.n2859 VSS.n2400 4.5005
R20306 VSS.n3051 VSS.n2432 4.5005
R20307 VSS.n2432 VSS.n2351 4.5005
R20308 VSS.n2483 VSS.n2432 4.5005
R20309 VSS.n2484 VSS.n2432 4.5005
R20310 VSS.n2486 VSS.n2432 4.5005
R20311 VSS.n2489 VSS.n2432 4.5005
R20312 VSS.n2491 VSS.n2432 4.5005
R20313 VSS.n2492 VSS.n2432 4.5005
R20314 VSS.n2494 VSS.n2432 4.5005
R20315 VSS.n2497 VSS.n2432 4.5005
R20316 VSS.n2499 VSS.n2432 4.5005
R20317 VSS.n2500 VSS.n2432 4.5005
R20318 VSS.n2502 VSS.n2432 4.5005
R20319 VSS.n2505 VSS.n2432 4.5005
R20320 VSS.n2507 VSS.n2432 4.5005
R20321 VSS.n2508 VSS.n2432 4.5005
R20322 VSS.n2510 VSS.n2432 4.5005
R20323 VSS.n2513 VSS.n2432 4.5005
R20324 VSS.n2515 VSS.n2432 4.5005
R20325 VSS.n2516 VSS.n2432 4.5005
R20326 VSS.n2518 VSS.n2432 4.5005
R20327 VSS.n2521 VSS.n2432 4.5005
R20328 VSS.n2523 VSS.n2432 4.5005
R20329 VSS.n2524 VSS.n2432 4.5005
R20330 VSS.n2526 VSS.n2432 4.5005
R20331 VSS.n2529 VSS.n2432 4.5005
R20332 VSS.n2531 VSS.n2432 4.5005
R20333 VSS.n2532 VSS.n2432 4.5005
R20334 VSS.n2534 VSS.n2432 4.5005
R20335 VSS.n2537 VSS.n2432 4.5005
R20336 VSS.n2539 VSS.n2432 4.5005
R20337 VSS.n2540 VSS.n2432 4.5005
R20338 VSS.n2542 VSS.n2432 4.5005
R20339 VSS.n2545 VSS.n2432 4.5005
R20340 VSS.n2547 VSS.n2432 4.5005
R20341 VSS.n2548 VSS.n2432 4.5005
R20342 VSS.n2550 VSS.n2432 4.5005
R20343 VSS.n2553 VSS.n2432 4.5005
R20344 VSS.n2555 VSS.n2432 4.5005
R20345 VSS.n2556 VSS.n2432 4.5005
R20346 VSS.n2558 VSS.n2432 4.5005
R20347 VSS.n2561 VSS.n2432 4.5005
R20348 VSS.n2563 VSS.n2432 4.5005
R20349 VSS.n2564 VSS.n2432 4.5005
R20350 VSS.n2566 VSS.n2432 4.5005
R20351 VSS.n2569 VSS.n2432 4.5005
R20352 VSS.n2571 VSS.n2432 4.5005
R20353 VSS.n2572 VSS.n2432 4.5005
R20354 VSS.n2574 VSS.n2432 4.5005
R20355 VSS.n2577 VSS.n2432 4.5005
R20356 VSS.n2579 VSS.n2432 4.5005
R20357 VSS.n2580 VSS.n2432 4.5005
R20358 VSS.n2582 VSS.n2432 4.5005
R20359 VSS.n2585 VSS.n2432 4.5005
R20360 VSS.n2587 VSS.n2432 4.5005
R20361 VSS.n2588 VSS.n2432 4.5005
R20362 VSS.n2590 VSS.n2432 4.5005
R20363 VSS.n2593 VSS.n2432 4.5005
R20364 VSS.n2595 VSS.n2432 4.5005
R20365 VSS.n2596 VSS.n2432 4.5005
R20366 VSS.n2598 VSS.n2432 4.5005
R20367 VSS.n2601 VSS.n2432 4.5005
R20368 VSS.n2603 VSS.n2432 4.5005
R20369 VSS.n2604 VSS.n2432 4.5005
R20370 VSS.n2606 VSS.n2432 4.5005
R20371 VSS.n2609 VSS.n2432 4.5005
R20372 VSS.n2611 VSS.n2432 4.5005
R20373 VSS.n2612 VSS.n2432 4.5005
R20374 VSS.n2614 VSS.n2432 4.5005
R20375 VSS.n2617 VSS.n2432 4.5005
R20376 VSS.n2619 VSS.n2432 4.5005
R20377 VSS.n2620 VSS.n2432 4.5005
R20378 VSS.n2622 VSS.n2432 4.5005
R20379 VSS.n2625 VSS.n2432 4.5005
R20380 VSS.n2627 VSS.n2432 4.5005
R20381 VSS.n2628 VSS.n2432 4.5005
R20382 VSS.n2630 VSS.n2432 4.5005
R20383 VSS.n2633 VSS.n2432 4.5005
R20384 VSS.n2635 VSS.n2432 4.5005
R20385 VSS.n2636 VSS.n2432 4.5005
R20386 VSS.n2638 VSS.n2432 4.5005
R20387 VSS.n2640 VSS.n2432 4.5005
R20388 VSS.n2642 VSS.n2432 4.5005
R20389 VSS.n2643 VSS.n2432 4.5005
R20390 VSS.n2645 VSS.n2432 4.5005
R20391 VSS.n2648 VSS.n2432 4.5005
R20392 VSS.n2650 VSS.n2432 4.5005
R20393 VSS.n2651 VSS.n2432 4.5005
R20394 VSS.n2653 VSS.n2432 4.5005
R20395 VSS.n2656 VSS.n2432 4.5005
R20396 VSS.n2658 VSS.n2432 4.5005
R20397 VSS.n2659 VSS.n2432 4.5005
R20398 VSS.n2661 VSS.n2432 4.5005
R20399 VSS.n2664 VSS.n2432 4.5005
R20400 VSS.n2666 VSS.n2432 4.5005
R20401 VSS.n2667 VSS.n2432 4.5005
R20402 VSS.n2669 VSS.n2432 4.5005
R20403 VSS.n2672 VSS.n2432 4.5005
R20404 VSS.n2674 VSS.n2432 4.5005
R20405 VSS.n2675 VSS.n2432 4.5005
R20406 VSS.n2677 VSS.n2432 4.5005
R20407 VSS.n2680 VSS.n2432 4.5005
R20408 VSS.n2682 VSS.n2432 4.5005
R20409 VSS.n2683 VSS.n2432 4.5005
R20410 VSS.n2685 VSS.n2432 4.5005
R20411 VSS.n2688 VSS.n2432 4.5005
R20412 VSS.n2690 VSS.n2432 4.5005
R20413 VSS.n2691 VSS.n2432 4.5005
R20414 VSS.n2693 VSS.n2432 4.5005
R20415 VSS.n2696 VSS.n2432 4.5005
R20416 VSS.n2698 VSS.n2432 4.5005
R20417 VSS.n2699 VSS.n2432 4.5005
R20418 VSS.n2701 VSS.n2432 4.5005
R20419 VSS.n2704 VSS.n2432 4.5005
R20420 VSS.n2706 VSS.n2432 4.5005
R20421 VSS.n2707 VSS.n2432 4.5005
R20422 VSS.n2709 VSS.n2432 4.5005
R20423 VSS.n2712 VSS.n2432 4.5005
R20424 VSS.n2714 VSS.n2432 4.5005
R20425 VSS.n2715 VSS.n2432 4.5005
R20426 VSS.n2717 VSS.n2432 4.5005
R20427 VSS.n2720 VSS.n2432 4.5005
R20428 VSS.n2722 VSS.n2432 4.5005
R20429 VSS.n2723 VSS.n2432 4.5005
R20430 VSS.n2725 VSS.n2432 4.5005
R20431 VSS.n2793 VSS.n2432 4.5005
R20432 VSS.n2859 VSS.n2432 4.5005
R20433 VSS.n3051 VSS.n2399 4.5005
R20434 VSS.n2399 VSS.n2351 4.5005
R20435 VSS.n2483 VSS.n2399 4.5005
R20436 VSS.n2484 VSS.n2399 4.5005
R20437 VSS.n2486 VSS.n2399 4.5005
R20438 VSS.n2489 VSS.n2399 4.5005
R20439 VSS.n2491 VSS.n2399 4.5005
R20440 VSS.n2492 VSS.n2399 4.5005
R20441 VSS.n2494 VSS.n2399 4.5005
R20442 VSS.n2497 VSS.n2399 4.5005
R20443 VSS.n2499 VSS.n2399 4.5005
R20444 VSS.n2500 VSS.n2399 4.5005
R20445 VSS.n2502 VSS.n2399 4.5005
R20446 VSS.n2505 VSS.n2399 4.5005
R20447 VSS.n2507 VSS.n2399 4.5005
R20448 VSS.n2508 VSS.n2399 4.5005
R20449 VSS.n2510 VSS.n2399 4.5005
R20450 VSS.n2513 VSS.n2399 4.5005
R20451 VSS.n2515 VSS.n2399 4.5005
R20452 VSS.n2516 VSS.n2399 4.5005
R20453 VSS.n2518 VSS.n2399 4.5005
R20454 VSS.n2521 VSS.n2399 4.5005
R20455 VSS.n2523 VSS.n2399 4.5005
R20456 VSS.n2524 VSS.n2399 4.5005
R20457 VSS.n2526 VSS.n2399 4.5005
R20458 VSS.n2529 VSS.n2399 4.5005
R20459 VSS.n2531 VSS.n2399 4.5005
R20460 VSS.n2532 VSS.n2399 4.5005
R20461 VSS.n2534 VSS.n2399 4.5005
R20462 VSS.n2537 VSS.n2399 4.5005
R20463 VSS.n2539 VSS.n2399 4.5005
R20464 VSS.n2540 VSS.n2399 4.5005
R20465 VSS.n2542 VSS.n2399 4.5005
R20466 VSS.n2545 VSS.n2399 4.5005
R20467 VSS.n2547 VSS.n2399 4.5005
R20468 VSS.n2548 VSS.n2399 4.5005
R20469 VSS.n2550 VSS.n2399 4.5005
R20470 VSS.n2553 VSS.n2399 4.5005
R20471 VSS.n2555 VSS.n2399 4.5005
R20472 VSS.n2556 VSS.n2399 4.5005
R20473 VSS.n2558 VSS.n2399 4.5005
R20474 VSS.n2561 VSS.n2399 4.5005
R20475 VSS.n2563 VSS.n2399 4.5005
R20476 VSS.n2564 VSS.n2399 4.5005
R20477 VSS.n2566 VSS.n2399 4.5005
R20478 VSS.n2569 VSS.n2399 4.5005
R20479 VSS.n2571 VSS.n2399 4.5005
R20480 VSS.n2572 VSS.n2399 4.5005
R20481 VSS.n2574 VSS.n2399 4.5005
R20482 VSS.n2577 VSS.n2399 4.5005
R20483 VSS.n2579 VSS.n2399 4.5005
R20484 VSS.n2580 VSS.n2399 4.5005
R20485 VSS.n2582 VSS.n2399 4.5005
R20486 VSS.n2585 VSS.n2399 4.5005
R20487 VSS.n2587 VSS.n2399 4.5005
R20488 VSS.n2588 VSS.n2399 4.5005
R20489 VSS.n2590 VSS.n2399 4.5005
R20490 VSS.n2593 VSS.n2399 4.5005
R20491 VSS.n2595 VSS.n2399 4.5005
R20492 VSS.n2596 VSS.n2399 4.5005
R20493 VSS.n2598 VSS.n2399 4.5005
R20494 VSS.n2601 VSS.n2399 4.5005
R20495 VSS.n2603 VSS.n2399 4.5005
R20496 VSS.n2604 VSS.n2399 4.5005
R20497 VSS.n2606 VSS.n2399 4.5005
R20498 VSS.n2609 VSS.n2399 4.5005
R20499 VSS.n2611 VSS.n2399 4.5005
R20500 VSS.n2612 VSS.n2399 4.5005
R20501 VSS.n2614 VSS.n2399 4.5005
R20502 VSS.n2617 VSS.n2399 4.5005
R20503 VSS.n2619 VSS.n2399 4.5005
R20504 VSS.n2620 VSS.n2399 4.5005
R20505 VSS.n2622 VSS.n2399 4.5005
R20506 VSS.n2625 VSS.n2399 4.5005
R20507 VSS.n2627 VSS.n2399 4.5005
R20508 VSS.n2628 VSS.n2399 4.5005
R20509 VSS.n2630 VSS.n2399 4.5005
R20510 VSS.n2633 VSS.n2399 4.5005
R20511 VSS.n2635 VSS.n2399 4.5005
R20512 VSS.n2636 VSS.n2399 4.5005
R20513 VSS.n2638 VSS.n2399 4.5005
R20514 VSS.n2640 VSS.n2399 4.5005
R20515 VSS.n2642 VSS.n2399 4.5005
R20516 VSS.n2643 VSS.n2399 4.5005
R20517 VSS.n2645 VSS.n2399 4.5005
R20518 VSS.n2648 VSS.n2399 4.5005
R20519 VSS.n2650 VSS.n2399 4.5005
R20520 VSS.n2651 VSS.n2399 4.5005
R20521 VSS.n2653 VSS.n2399 4.5005
R20522 VSS.n2656 VSS.n2399 4.5005
R20523 VSS.n2658 VSS.n2399 4.5005
R20524 VSS.n2659 VSS.n2399 4.5005
R20525 VSS.n2661 VSS.n2399 4.5005
R20526 VSS.n2664 VSS.n2399 4.5005
R20527 VSS.n2666 VSS.n2399 4.5005
R20528 VSS.n2667 VSS.n2399 4.5005
R20529 VSS.n2669 VSS.n2399 4.5005
R20530 VSS.n2672 VSS.n2399 4.5005
R20531 VSS.n2674 VSS.n2399 4.5005
R20532 VSS.n2675 VSS.n2399 4.5005
R20533 VSS.n2677 VSS.n2399 4.5005
R20534 VSS.n2680 VSS.n2399 4.5005
R20535 VSS.n2682 VSS.n2399 4.5005
R20536 VSS.n2683 VSS.n2399 4.5005
R20537 VSS.n2685 VSS.n2399 4.5005
R20538 VSS.n2688 VSS.n2399 4.5005
R20539 VSS.n2690 VSS.n2399 4.5005
R20540 VSS.n2691 VSS.n2399 4.5005
R20541 VSS.n2693 VSS.n2399 4.5005
R20542 VSS.n2696 VSS.n2399 4.5005
R20543 VSS.n2698 VSS.n2399 4.5005
R20544 VSS.n2699 VSS.n2399 4.5005
R20545 VSS.n2701 VSS.n2399 4.5005
R20546 VSS.n2704 VSS.n2399 4.5005
R20547 VSS.n2706 VSS.n2399 4.5005
R20548 VSS.n2707 VSS.n2399 4.5005
R20549 VSS.n2709 VSS.n2399 4.5005
R20550 VSS.n2712 VSS.n2399 4.5005
R20551 VSS.n2714 VSS.n2399 4.5005
R20552 VSS.n2715 VSS.n2399 4.5005
R20553 VSS.n2717 VSS.n2399 4.5005
R20554 VSS.n2720 VSS.n2399 4.5005
R20555 VSS.n2722 VSS.n2399 4.5005
R20556 VSS.n2723 VSS.n2399 4.5005
R20557 VSS.n2725 VSS.n2399 4.5005
R20558 VSS.n2793 VSS.n2399 4.5005
R20559 VSS.n2859 VSS.n2399 4.5005
R20560 VSS.n3051 VSS.n2433 4.5005
R20561 VSS.n2433 VSS.n2351 4.5005
R20562 VSS.n2483 VSS.n2433 4.5005
R20563 VSS.n2484 VSS.n2433 4.5005
R20564 VSS.n2486 VSS.n2433 4.5005
R20565 VSS.n2489 VSS.n2433 4.5005
R20566 VSS.n2491 VSS.n2433 4.5005
R20567 VSS.n2492 VSS.n2433 4.5005
R20568 VSS.n2494 VSS.n2433 4.5005
R20569 VSS.n2497 VSS.n2433 4.5005
R20570 VSS.n2499 VSS.n2433 4.5005
R20571 VSS.n2500 VSS.n2433 4.5005
R20572 VSS.n2502 VSS.n2433 4.5005
R20573 VSS.n2505 VSS.n2433 4.5005
R20574 VSS.n2507 VSS.n2433 4.5005
R20575 VSS.n2508 VSS.n2433 4.5005
R20576 VSS.n2510 VSS.n2433 4.5005
R20577 VSS.n2513 VSS.n2433 4.5005
R20578 VSS.n2515 VSS.n2433 4.5005
R20579 VSS.n2516 VSS.n2433 4.5005
R20580 VSS.n2518 VSS.n2433 4.5005
R20581 VSS.n2521 VSS.n2433 4.5005
R20582 VSS.n2523 VSS.n2433 4.5005
R20583 VSS.n2524 VSS.n2433 4.5005
R20584 VSS.n2526 VSS.n2433 4.5005
R20585 VSS.n2529 VSS.n2433 4.5005
R20586 VSS.n2531 VSS.n2433 4.5005
R20587 VSS.n2532 VSS.n2433 4.5005
R20588 VSS.n2534 VSS.n2433 4.5005
R20589 VSS.n2537 VSS.n2433 4.5005
R20590 VSS.n2539 VSS.n2433 4.5005
R20591 VSS.n2540 VSS.n2433 4.5005
R20592 VSS.n2542 VSS.n2433 4.5005
R20593 VSS.n2545 VSS.n2433 4.5005
R20594 VSS.n2547 VSS.n2433 4.5005
R20595 VSS.n2548 VSS.n2433 4.5005
R20596 VSS.n2550 VSS.n2433 4.5005
R20597 VSS.n2553 VSS.n2433 4.5005
R20598 VSS.n2555 VSS.n2433 4.5005
R20599 VSS.n2556 VSS.n2433 4.5005
R20600 VSS.n2558 VSS.n2433 4.5005
R20601 VSS.n2561 VSS.n2433 4.5005
R20602 VSS.n2563 VSS.n2433 4.5005
R20603 VSS.n2564 VSS.n2433 4.5005
R20604 VSS.n2566 VSS.n2433 4.5005
R20605 VSS.n2569 VSS.n2433 4.5005
R20606 VSS.n2571 VSS.n2433 4.5005
R20607 VSS.n2572 VSS.n2433 4.5005
R20608 VSS.n2574 VSS.n2433 4.5005
R20609 VSS.n2577 VSS.n2433 4.5005
R20610 VSS.n2579 VSS.n2433 4.5005
R20611 VSS.n2580 VSS.n2433 4.5005
R20612 VSS.n2582 VSS.n2433 4.5005
R20613 VSS.n2585 VSS.n2433 4.5005
R20614 VSS.n2587 VSS.n2433 4.5005
R20615 VSS.n2588 VSS.n2433 4.5005
R20616 VSS.n2590 VSS.n2433 4.5005
R20617 VSS.n2593 VSS.n2433 4.5005
R20618 VSS.n2595 VSS.n2433 4.5005
R20619 VSS.n2596 VSS.n2433 4.5005
R20620 VSS.n2598 VSS.n2433 4.5005
R20621 VSS.n2601 VSS.n2433 4.5005
R20622 VSS.n2603 VSS.n2433 4.5005
R20623 VSS.n2604 VSS.n2433 4.5005
R20624 VSS.n2606 VSS.n2433 4.5005
R20625 VSS.n2609 VSS.n2433 4.5005
R20626 VSS.n2611 VSS.n2433 4.5005
R20627 VSS.n2612 VSS.n2433 4.5005
R20628 VSS.n2614 VSS.n2433 4.5005
R20629 VSS.n2617 VSS.n2433 4.5005
R20630 VSS.n2619 VSS.n2433 4.5005
R20631 VSS.n2620 VSS.n2433 4.5005
R20632 VSS.n2622 VSS.n2433 4.5005
R20633 VSS.n2625 VSS.n2433 4.5005
R20634 VSS.n2627 VSS.n2433 4.5005
R20635 VSS.n2628 VSS.n2433 4.5005
R20636 VSS.n2630 VSS.n2433 4.5005
R20637 VSS.n2633 VSS.n2433 4.5005
R20638 VSS.n2635 VSS.n2433 4.5005
R20639 VSS.n2636 VSS.n2433 4.5005
R20640 VSS.n2638 VSS.n2433 4.5005
R20641 VSS.n2640 VSS.n2433 4.5005
R20642 VSS.n2642 VSS.n2433 4.5005
R20643 VSS.n2643 VSS.n2433 4.5005
R20644 VSS.n2645 VSS.n2433 4.5005
R20645 VSS.n2648 VSS.n2433 4.5005
R20646 VSS.n2650 VSS.n2433 4.5005
R20647 VSS.n2651 VSS.n2433 4.5005
R20648 VSS.n2653 VSS.n2433 4.5005
R20649 VSS.n2656 VSS.n2433 4.5005
R20650 VSS.n2658 VSS.n2433 4.5005
R20651 VSS.n2659 VSS.n2433 4.5005
R20652 VSS.n2661 VSS.n2433 4.5005
R20653 VSS.n2664 VSS.n2433 4.5005
R20654 VSS.n2666 VSS.n2433 4.5005
R20655 VSS.n2667 VSS.n2433 4.5005
R20656 VSS.n2669 VSS.n2433 4.5005
R20657 VSS.n2672 VSS.n2433 4.5005
R20658 VSS.n2674 VSS.n2433 4.5005
R20659 VSS.n2675 VSS.n2433 4.5005
R20660 VSS.n2677 VSS.n2433 4.5005
R20661 VSS.n2680 VSS.n2433 4.5005
R20662 VSS.n2682 VSS.n2433 4.5005
R20663 VSS.n2683 VSS.n2433 4.5005
R20664 VSS.n2685 VSS.n2433 4.5005
R20665 VSS.n2688 VSS.n2433 4.5005
R20666 VSS.n2690 VSS.n2433 4.5005
R20667 VSS.n2691 VSS.n2433 4.5005
R20668 VSS.n2693 VSS.n2433 4.5005
R20669 VSS.n2696 VSS.n2433 4.5005
R20670 VSS.n2698 VSS.n2433 4.5005
R20671 VSS.n2699 VSS.n2433 4.5005
R20672 VSS.n2701 VSS.n2433 4.5005
R20673 VSS.n2704 VSS.n2433 4.5005
R20674 VSS.n2706 VSS.n2433 4.5005
R20675 VSS.n2707 VSS.n2433 4.5005
R20676 VSS.n2709 VSS.n2433 4.5005
R20677 VSS.n2712 VSS.n2433 4.5005
R20678 VSS.n2714 VSS.n2433 4.5005
R20679 VSS.n2715 VSS.n2433 4.5005
R20680 VSS.n2717 VSS.n2433 4.5005
R20681 VSS.n2720 VSS.n2433 4.5005
R20682 VSS.n2722 VSS.n2433 4.5005
R20683 VSS.n2723 VSS.n2433 4.5005
R20684 VSS.n2725 VSS.n2433 4.5005
R20685 VSS.n2793 VSS.n2433 4.5005
R20686 VSS.n2859 VSS.n2433 4.5005
R20687 VSS.n3051 VSS.n2398 4.5005
R20688 VSS.n2398 VSS.n2351 4.5005
R20689 VSS.n2483 VSS.n2398 4.5005
R20690 VSS.n2484 VSS.n2398 4.5005
R20691 VSS.n2486 VSS.n2398 4.5005
R20692 VSS.n2489 VSS.n2398 4.5005
R20693 VSS.n2491 VSS.n2398 4.5005
R20694 VSS.n2492 VSS.n2398 4.5005
R20695 VSS.n2494 VSS.n2398 4.5005
R20696 VSS.n2497 VSS.n2398 4.5005
R20697 VSS.n2499 VSS.n2398 4.5005
R20698 VSS.n2500 VSS.n2398 4.5005
R20699 VSS.n2502 VSS.n2398 4.5005
R20700 VSS.n2505 VSS.n2398 4.5005
R20701 VSS.n2507 VSS.n2398 4.5005
R20702 VSS.n2508 VSS.n2398 4.5005
R20703 VSS.n2510 VSS.n2398 4.5005
R20704 VSS.n2513 VSS.n2398 4.5005
R20705 VSS.n2515 VSS.n2398 4.5005
R20706 VSS.n2516 VSS.n2398 4.5005
R20707 VSS.n2518 VSS.n2398 4.5005
R20708 VSS.n2521 VSS.n2398 4.5005
R20709 VSS.n2523 VSS.n2398 4.5005
R20710 VSS.n2524 VSS.n2398 4.5005
R20711 VSS.n2526 VSS.n2398 4.5005
R20712 VSS.n2529 VSS.n2398 4.5005
R20713 VSS.n2531 VSS.n2398 4.5005
R20714 VSS.n2532 VSS.n2398 4.5005
R20715 VSS.n2534 VSS.n2398 4.5005
R20716 VSS.n2537 VSS.n2398 4.5005
R20717 VSS.n2539 VSS.n2398 4.5005
R20718 VSS.n2540 VSS.n2398 4.5005
R20719 VSS.n2542 VSS.n2398 4.5005
R20720 VSS.n2545 VSS.n2398 4.5005
R20721 VSS.n2547 VSS.n2398 4.5005
R20722 VSS.n2548 VSS.n2398 4.5005
R20723 VSS.n2550 VSS.n2398 4.5005
R20724 VSS.n2553 VSS.n2398 4.5005
R20725 VSS.n2555 VSS.n2398 4.5005
R20726 VSS.n2556 VSS.n2398 4.5005
R20727 VSS.n2558 VSS.n2398 4.5005
R20728 VSS.n2561 VSS.n2398 4.5005
R20729 VSS.n2563 VSS.n2398 4.5005
R20730 VSS.n2564 VSS.n2398 4.5005
R20731 VSS.n2566 VSS.n2398 4.5005
R20732 VSS.n2569 VSS.n2398 4.5005
R20733 VSS.n2571 VSS.n2398 4.5005
R20734 VSS.n2572 VSS.n2398 4.5005
R20735 VSS.n2574 VSS.n2398 4.5005
R20736 VSS.n2577 VSS.n2398 4.5005
R20737 VSS.n2579 VSS.n2398 4.5005
R20738 VSS.n2580 VSS.n2398 4.5005
R20739 VSS.n2582 VSS.n2398 4.5005
R20740 VSS.n2585 VSS.n2398 4.5005
R20741 VSS.n2587 VSS.n2398 4.5005
R20742 VSS.n2588 VSS.n2398 4.5005
R20743 VSS.n2590 VSS.n2398 4.5005
R20744 VSS.n2593 VSS.n2398 4.5005
R20745 VSS.n2595 VSS.n2398 4.5005
R20746 VSS.n2596 VSS.n2398 4.5005
R20747 VSS.n2598 VSS.n2398 4.5005
R20748 VSS.n2601 VSS.n2398 4.5005
R20749 VSS.n2603 VSS.n2398 4.5005
R20750 VSS.n2604 VSS.n2398 4.5005
R20751 VSS.n2606 VSS.n2398 4.5005
R20752 VSS.n2609 VSS.n2398 4.5005
R20753 VSS.n2611 VSS.n2398 4.5005
R20754 VSS.n2612 VSS.n2398 4.5005
R20755 VSS.n2614 VSS.n2398 4.5005
R20756 VSS.n2617 VSS.n2398 4.5005
R20757 VSS.n2619 VSS.n2398 4.5005
R20758 VSS.n2620 VSS.n2398 4.5005
R20759 VSS.n2622 VSS.n2398 4.5005
R20760 VSS.n2625 VSS.n2398 4.5005
R20761 VSS.n2627 VSS.n2398 4.5005
R20762 VSS.n2628 VSS.n2398 4.5005
R20763 VSS.n2630 VSS.n2398 4.5005
R20764 VSS.n2633 VSS.n2398 4.5005
R20765 VSS.n2635 VSS.n2398 4.5005
R20766 VSS.n2636 VSS.n2398 4.5005
R20767 VSS.n2638 VSS.n2398 4.5005
R20768 VSS.n2640 VSS.n2398 4.5005
R20769 VSS.n2642 VSS.n2398 4.5005
R20770 VSS.n2643 VSS.n2398 4.5005
R20771 VSS.n2645 VSS.n2398 4.5005
R20772 VSS.n2648 VSS.n2398 4.5005
R20773 VSS.n2650 VSS.n2398 4.5005
R20774 VSS.n2651 VSS.n2398 4.5005
R20775 VSS.n2653 VSS.n2398 4.5005
R20776 VSS.n2656 VSS.n2398 4.5005
R20777 VSS.n2658 VSS.n2398 4.5005
R20778 VSS.n2659 VSS.n2398 4.5005
R20779 VSS.n2661 VSS.n2398 4.5005
R20780 VSS.n2664 VSS.n2398 4.5005
R20781 VSS.n2666 VSS.n2398 4.5005
R20782 VSS.n2667 VSS.n2398 4.5005
R20783 VSS.n2669 VSS.n2398 4.5005
R20784 VSS.n2672 VSS.n2398 4.5005
R20785 VSS.n2674 VSS.n2398 4.5005
R20786 VSS.n2675 VSS.n2398 4.5005
R20787 VSS.n2677 VSS.n2398 4.5005
R20788 VSS.n2680 VSS.n2398 4.5005
R20789 VSS.n2682 VSS.n2398 4.5005
R20790 VSS.n2683 VSS.n2398 4.5005
R20791 VSS.n2685 VSS.n2398 4.5005
R20792 VSS.n2688 VSS.n2398 4.5005
R20793 VSS.n2690 VSS.n2398 4.5005
R20794 VSS.n2691 VSS.n2398 4.5005
R20795 VSS.n2693 VSS.n2398 4.5005
R20796 VSS.n2696 VSS.n2398 4.5005
R20797 VSS.n2698 VSS.n2398 4.5005
R20798 VSS.n2699 VSS.n2398 4.5005
R20799 VSS.n2701 VSS.n2398 4.5005
R20800 VSS.n2704 VSS.n2398 4.5005
R20801 VSS.n2706 VSS.n2398 4.5005
R20802 VSS.n2707 VSS.n2398 4.5005
R20803 VSS.n2709 VSS.n2398 4.5005
R20804 VSS.n2712 VSS.n2398 4.5005
R20805 VSS.n2714 VSS.n2398 4.5005
R20806 VSS.n2715 VSS.n2398 4.5005
R20807 VSS.n2717 VSS.n2398 4.5005
R20808 VSS.n2720 VSS.n2398 4.5005
R20809 VSS.n2722 VSS.n2398 4.5005
R20810 VSS.n2723 VSS.n2398 4.5005
R20811 VSS.n2725 VSS.n2398 4.5005
R20812 VSS.n2793 VSS.n2398 4.5005
R20813 VSS.n2859 VSS.n2398 4.5005
R20814 VSS.n3051 VSS.n2434 4.5005
R20815 VSS.n2434 VSS.n2351 4.5005
R20816 VSS.n2483 VSS.n2434 4.5005
R20817 VSS.n2484 VSS.n2434 4.5005
R20818 VSS.n2486 VSS.n2434 4.5005
R20819 VSS.n2489 VSS.n2434 4.5005
R20820 VSS.n2491 VSS.n2434 4.5005
R20821 VSS.n2492 VSS.n2434 4.5005
R20822 VSS.n2494 VSS.n2434 4.5005
R20823 VSS.n2497 VSS.n2434 4.5005
R20824 VSS.n2499 VSS.n2434 4.5005
R20825 VSS.n2500 VSS.n2434 4.5005
R20826 VSS.n2502 VSS.n2434 4.5005
R20827 VSS.n2505 VSS.n2434 4.5005
R20828 VSS.n2507 VSS.n2434 4.5005
R20829 VSS.n2508 VSS.n2434 4.5005
R20830 VSS.n2510 VSS.n2434 4.5005
R20831 VSS.n2513 VSS.n2434 4.5005
R20832 VSS.n2515 VSS.n2434 4.5005
R20833 VSS.n2516 VSS.n2434 4.5005
R20834 VSS.n2518 VSS.n2434 4.5005
R20835 VSS.n2521 VSS.n2434 4.5005
R20836 VSS.n2523 VSS.n2434 4.5005
R20837 VSS.n2524 VSS.n2434 4.5005
R20838 VSS.n2526 VSS.n2434 4.5005
R20839 VSS.n2529 VSS.n2434 4.5005
R20840 VSS.n2531 VSS.n2434 4.5005
R20841 VSS.n2532 VSS.n2434 4.5005
R20842 VSS.n2534 VSS.n2434 4.5005
R20843 VSS.n2537 VSS.n2434 4.5005
R20844 VSS.n2539 VSS.n2434 4.5005
R20845 VSS.n2540 VSS.n2434 4.5005
R20846 VSS.n2542 VSS.n2434 4.5005
R20847 VSS.n2545 VSS.n2434 4.5005
R20848 VSS.n2547 VSS.n2434 4.5005
R20849 VSS.n2548 VSS.n2434 4.5005
R20850 VSS.n2550 VSS.n2434 4.5005
R20851 VSS.n2553 VSS.n2434 4.5005
R20852 VSS.n2555 VSS.n2434 4.5005
R20853 VSS.n2556 VSS.n2434 4.5005
R20854 VSS.n2558 VSS.n2434 4.5005
R20855 VSS.n2561 VSS.n2434 4.5005
R20856 VSS.n2563 VSS.n2434 4.5005
R20857 VSS.n2564 VSS.n2434 4.5005
R20858 VSS.n2566 VSS.n2434 4.5005
R20859 VSS.n2569 VSS.n2434 4.5005
R20860 VSS.n2571 VSS.n2434 4.5005
R20861 VSS.n2572 VSS.n2434 4.5005
R20862 VSS.n2574 VSS.n2434 4.5005
R20863 VSS.n2577 VSS.n2434 4.5005
R20864 VSS.n2579 VSS.n2434 4.5005
R20865 VSS.n2580 VSS.n2434 4.5005
R20866 VSS.n2582 VSS.n2434 4.5005
R20867 VSS.n2585 VSS.n2434 4.5005
R20868 VSS.n2587 VSS.n2434 4.5005
R20869 VSS.n2588 VSS.n2434 4.5005
R20870 VSS.n2590 VSS.n2434 4.5005
R20871 VSS.n2593 VSS.n2434 4.5005
R20872 VSS.n2595 VSS.n2434 4.5005
R20873 VSS.n2596 VSS.n2434 4.5005
R20874 VSS.n2598 VSS.n2434 4.5005
R20875 VSS.n2601 VSS.n2434 4.5005
R20876 VSS.n2603 VSS.n2434 4.5005
R20877 VSS.n2604 VSS.n2434 4.5005
R20878 VSS.n2606 VSS.n2434 4.5005
R20879 VSS.n2609 VSS.n2434 4.5005
R20880 VSS.n2611 VSS.n2434 4.5005
R20881 VSS.n2612 VSS.n2434 4.5005
R20882 VSS.n2614 VSS.n2434 4.5005
R20883 VSS.n2617 VSS.n2434 4.5005
R20884 VSS.n2619 VSS.n2434 4.5005
R20885 VSS.n2620 VSS.n2434 4.5005
R20886 VSS.n2622 VSS.n2434 4.5005
R20887 VSS.n2625 VSS.n2434 4.5005
R20888 VSS.n2627 VSS.n2434 4.5005
R20889 VSS.n2628 VSS.n2434 4.5005
R20890 VSS.n2630 VSS.n2434 4.5005
R20891 VSS.n2633 VSS.n2434 4.5005
R20892 VSS.n2635 VSS.n2434 4.5005
R20893 VSS.n2636 VSS.n2434 4.5005
R20894 VSS.n2638 VSS.n2434 4.5005
R20895 VSS.n2640 VSS.n2434 4.5005
R20896 VSS.n2642 VSS.n2434 4.5005
R20897 VSS.n2643 VSS.n2434 4.5005
R20898 VSS.n2645 VSS.n2434 4.5005
R20899 VSS.n2648 VSS.n2434 4.5005
R20900 VSS.n2650 VSS.n2434 4.5005
R20901 VSS.n2651 VSS.n2434 4.5005
R20902 VSS.n2653 VSS.n2434 4.5005
R20903 VSS.n2656 VSS.n2434 4.5005
R20904 VSS.n2658 VSS.n2434 4.5005
R20905 VSS.n2659 VSS.n2434 4.5005
R20906 VSS.n2661 VSS.n2434 4.5005
R20907 VSS.n2664 VSS.n2434 4.5005
R20908 VSS.n2666 VSS.n2434 4.5005
R20909 VSS.n2667 VSS.n2434 4.5005
R20910 VSS.n2669 VSS.n2434 4.5005
R20911 VSS.n2672 VSS.n2434 4.5005
R20912 VSS.n2674 VSS.n2434 4.5005
R20913 VSS.n2675 VSS.n2434 4.5005
R20914 VSS.n2677 VSS.n2434 4.5005
R20915 VSS.n2680 VSS.n2434 4.5005
R20916 VSS.n2682 VSS.n2434 4.5005
R20917 VSS.n2683 VSS.n2434 4.5005
R20918 VSS.n2685 VSS.n2434 4.5005
R20919 VSS.n2688 VSS.n2434 4.5005
R20920 VSS.n2690 VSS.n2434 4.5005
R20921 VSS.n2691 VSS.n2434 4.5005
R20922 VSS.n2693 VSS.n2434 4.5005
R20923 VSS.n2696 VSS.n2434 4.5005
R20924 VSS.n2698 VSS.n2434 4.5005
R20925 VSS.n2699 VSS.n2434 4.5005
R20926 VSS.n2701 VSS.n2434 4.5005
R20927 VSS.n2704 VSS.n2434 4.5005
R20928 VSS.n2706 VSS.n2434 4.5005
R20929 VSS.n2707 VSS.n2434 4.5005
R20930 VSS.n2709 VSS.n2434 4.5005
R20931 VSS.n2712 VSS.n2434 4.5005
R20932 VSS.n2714 VSS.n2434 4.5005
R20933 VSS.n2715 VSS.n2434 4.5005
R20934 VSS.n2717 VSS.n2434 4.5005
R20935 VSS.n2720 VSS.n2434 4.5005
R20936 VSS.n2722 VSS.n2434 4.5005
R20937 VSS.n2723 VSS.n2434 4.5005
R20938 VSS.n2725 VSS.n2434 4.5005
R20939 VSS.n2793 VSS.n2434 4.5005
R20940 VSS.n2859 VSS.n2434 4.5005
R20941 VSS.n3051 VSS.n2397 4.5005
R20942 VSS.n2397 VSS.n2351 4.5005
R20943 VSS.n2483 VSS.n2397 4.5005
R20944 VSS.n2484 VSS.n2397 4.5005
R20945 VSS.n2486 VSS.n2397 4.5005
R20946 VSS.n2489 VSS.n2397 4.5005
R20947 VSS.n2491 VSS.n2397 4.5005
R20948 VSS.n2492 VSS.n2397 4.5005
R20949 VSS.n2494 VSS.n2397 4.5005
R20950 VSS.n2497 VSS.n2397 4.5005
R20951 VSS.n2499 VSS.n2397 4.5005
R20952 VSS.n2500 VSS.n2397 4.5005
R20953 VSS.n2502 VSS.n2397 4.5005
R20954 VSS.n2505 VSS.n2397 4.5005
R20955 VSS.n2507 VSS.n2397 4.5005
R20956 VSS.n2508 VSS.n2397 4.5005
R20957 VSS.n2510 VSS.n2397 4.5005
R20958 VSS.n2513 VSS.n2397 4.5005
R20959 VSS.n2515 VSS.n2397 4.5005
R20960 VSS.n2516 VSS.n2397 4.5005
R20961 VSS.n2518 VSS.n2397 4.5005
R20962 VSS.n2521 VSS.n2397 4.5005
R20963 VSS.n2523 VSS.n2397 4.5005
R20964 VSS.n2524 VSS.n2397 4.5005
R20965 VSS.n2526 VSS.n2397 4.5005
R20966 VSS.n2529 VSS.n2397 4.5005
R20967 VSS.n2531 VSS.n2397 4.5005
R20968 VSS.n2532 VSS.n2397 4.5005
R20969 VSS.n2534 VSS.n2397 4.5005
R20970 VSS.n2537 VSS.n2397 4.5005
R20971 VSS.n2539 VSS.n2397 4.5005
R20972 VSS.n2540 VSS.n2397 4.5005
R20973 VSS.n2542 VSS.n2397 4.5005
R20974 VSS.n2545 VSS.n2397 4.5005
R20975 VSS.n2547 VSS.n2397 4.5005
R20976 VSS.n2548 VSS.n2397 4.5005
R20977 VSS.n2550 VSS.n2397 4.5005
R20978 VSS.n2553 VSS.n2397 4.5005
R20979 VSS.n2555 VSS.n2397 4.5005
R20980 VSS.n2556 VSS.n2397 4.5005
R20981 VSS.n2558 VSS.n2397 4.5005
R20982 VSS.n2561 VSS.n2397 4.5005
R20983 VSS.n2563 VSS.n2397 4.5005
R20984 VSS.n2564 VSS.n2397 4.5005
R20985 VSS.n2566 VSS.n2397 4.5005
R20986 VSS.n2569 VSS.n2397 4.5005
R20987 VSS.n2571 VSS.n2397 4.5005
R20988 VSS.n2572 VSS.n2397 4.5005
R20989 VSS.n2574 VSS.n2397 4.5005
R20990 VSS.n2577 VSS.n2397 4.5005
R20991 VSS.n2579 VSS.n2397 4.5005
R20992 VSS.n2580 VSS.n2397 4.5005
R20993 VSS.n2582 VSS.n2397 4.5005
R20994 VSS.n2585 VSS.n2397 4.5005
R20995 VSS.n2587 VSS.n2397 4.5005
R20996 VSS.n2588 VSS.n2397 4.5005
R20997 VSS.n2590 VSS.n2397 4.5005
R20998 VSS.n2593 VSS.n2397 4.5005
R20999 VSS.n2595 VSS.n2397 4.5005
R21000 VSS.n2596 VSS.n2397 4.5005
R21001 VSS.n2598 VSS.n2397 4.5005
R21002 VSS.n2601 VSS.n2397 4.5005
R21003 VSS.n2603 VSS.n2397 4.5005
R21004 VSS.n2604 VSS.n2397 4.5005
R21005 VSS.n2606 VSS.n2397 4.5005
R21006 VSS.n2609 VSS.n2397 4.5005
R21007 VSS.n2611 VSS.n2397 4.5005
R21008 VSS.n2612 VSS.n2397 4.5005
R21009 VSS.n2614 VSS.n2397 4.5005
R21010 VSS.n2617 VSS.n2397 4.5005
R21011 VSS.n2619 VSS.n2397 4.5005
R21012 VSS.n2620 VSS.n2397 4.5005
R21013 VSS.n2622 VSS.n2397 4.5005
R21014 VSS.n2625 VSS.n2397 4.5005
R21015 VSS.n2627 VSS.n2397 4.5005
R21016 VSS.n2628 VSS.n2397 4.5005
R21017 VSS.n2630 VSS.n2397 4.5005
R21018 VSS.n2633 VSS.n2397 4.5005
R21019 VSS.n2635 VSS.n2397 4.5005
R21020 VSS.n2636 VSS.n2397 4.5005
R21021 VSS.n2638 VSS.n2397 4.5005
R21022 VSS.n2640 VSS.n2397 4.5005
R21023 VSS.n2642 VSS.n2397 4.5005
R21024 VSS.n2643 VSS.n2397 4.5005
R21025 VSS.n2645 VSS.n2397 4.5005
R21026 VSS.n2648 VSS.n2397 4.5005
R21027 VSS.n2650 VSS.n2397 4.5005
R21028 VSS.n2651 VSS.n2397 4.5005
R21029 VSS.n2653 VSS.n2397 4.5005
R21030 VSS.n2656 VSS.n2397 4.5005
R21031 VSS.n2658 VSS.n2397 4.5005
R21032 VSS.n2659 VSS.n2397 4.5005
R21033 VSS.n2661 VSS.n2397 4.5005
R21034 VSS.n2664 VSS.n2397 4.5005
R21035 VSS.n2666 VSS.n2397 4.5005
R21036 VSS.n2667 VSS.n2397 4.5005
R21037 VSS.n2669 VSS.n2397 4.5005
R21038 VSS.n2672 VSS.n2397 4.5005
R21039 VSS.n2674 VSS.n2397 4.5005
R21040 VSS.n2675 VSS.n2397 4.5005
R21041 VSS.n2677 VSS.n2397 4.5005
R21042 VSS.n2680 VSS.n2397 4.5005
R21043 VSS.n2682 VSS.n2397 4.5005
R21044 VSS.n2683 VSS.n2397 4.5005
R21045 VSS.n2685 VSS.n2397 4.5005
R21046 VSS.n2688 VSS.n2397 4.5005
R21047 VSS.n2690 VSS.n2397 4.5005
R21048 VSS.n2691 VSS.n2397 4.5005
R21049 VSS.n2693 VSS.n2397 4.5005
R21050 VSS.n2696 VSS.n2397 4.5005
R21051 VSS.n2698 VSS.n2397 4.5005
R21052 VSS.n2699 VSS.n2397 4.5005
R21053 VSS.n2701 VSS.n2397 4.5005
R21054 VSS.n2704 VSS.n2397 4.5005
R21055 VSS.n2706 VSS.n2397 4.5005
R21056 VSS.n2707 VSS.n2397 4.5005
R21057 VSS.n2709 VSS.n2397 4.5005
R21058 VSS.n2712 VSS.n2397 4.5005
R21059 VSS.n2714 VSS.n2397 4.5005
R21060 VSS.n2715 VSS.n2397 4.5005
R21061 VSS.n2717 VSS.n2397 4.5005
R21062 VSS.n2720 VSS.n2397 4.5005
R21063 VSS.n2722 VSS.n2397 4.5005
R21064 VSS.n2723 VSS.n2397 4.5005
R21065 VSS.n2725 VSS.n2397 4.5005
R21066 VSS.n2793 VSS.n2397 4.5005
R21067 VSS.n2859 VSS.n2397 4.5005
R21068 VSS.n3051 VSS.n2435 4.5005
R21069 VSS.n2435 VSS.n2351 4.5005
R21070 VSS.n2483 VSS.n2435 4.5005
R21071 VSS.n2484 VSS.n2435 4.5005
R21072 VSS.n2486 VSS.n2435 4.5005
R21073 VSS.n2489 VSS.n2435 4.5005
R21074 VSS.n2491 VSS.n2435 4.5005
R21075 VSS.n2492 VSS.n2435 4.5005
R21076 VSS.n2494 VSS.n2435 4.5005
R21077 VSS.n2497 VSS.n2435 4.5005
R21078 VSS.n2499 VSS.n2435 4.5005
R21079 VSS.n2500 VSS.n2435 4.5005
R21080 VSS.n2502 VSS.n2435 4.5005
R21081 VSS.n2505 VSS.n2435 4.5005
R21082 VSS.n2507 VSS.n2435 4.5005
R21083 VSS.n2508 VSS.n2435 4.5005
R21084 VSS.n2510 VSS.n2435 4.5005
R21085 VSS.n2513 VSS.n2435 4.5005
R21086 VSS.n2515 VSS.n2435 4.5005
R21087 VSS.n2516 VSS.n2435 4.5005
R21088 VSS.n2518 VSS.n2435 4.5005
R21089 VSS.n2521 VSS.n2435 4.5005
R21090 VSS.n2523 VSS.n2435 4.5005
R21091 VSS.n2524 VSS.n2435 4.5005
R21092 VSS.n2526 VSS.n2435 4.5005
R21093 VSS.n2529 VSS.n2435 4.5005
R21094 VSS.n2531 VSS.n2435 4.5005
R21095 VSS.n2532 VSS.n2435 4.5005
R21096 VSS.n2534 VSS.n2435 4.5005
R21097 VSS.n2537 VSS.n2435 4.5005
R21098 VSS.n2539 VSS.n2435 4.5005
R21099 VSS.n2540 VSS.n2435 4.5005
R21100 VSS.n2542 VSS.n2435 4.5005
R21101 VSS.n2545 VSS.n2435 4.5005
R21102 VSS.n2547 VSS.n2435 4.5005
R21103 VSS.n2548 VSS.n2435 4.5005
R21104 VSS.n2550 VSS.n2435 4.5005
R21105 VSS.n2553 VSS.n2435 4.5005
R21106 VSS.n2555 VSS.n2435 4.5005
R21107 VSS.n2556 VSS.n2435 4.5005
R21108 VSS.n2558 VSS.n2435 4.5005
R21109 VSS.n2561 VSS.n2435 4.5005
R21110 VSS.n2563 VSS.n2435 4.5005
R21111 VSS.n2564 VSS.n2435 4.5005
R21112 VSS.n2566 VSS.n2435 4.5005
R21113 VSS.n2569 VSS.n2435 4.5005
R21114 VSS.n2571 VSS.n2435 4.5005
R21115 VSS.n2572 VSS.n2435 4.5005
R21116 VSS.n2574 VSS.n2435 4.5005
R21117 VSS.n2577 VSS.n2435 4.5005
R21118 VSS.n2579 VSS.n2435 4.5005
R21119 VSS.n2580 VSS.n2435 4.5005
R21120 VSS.n2582 VSS.n2435 4.5005
R21121 VSS.n2585 VSS.n2435 4.5005
R21122 VSS.n2587 VSS.n2435 4.5005
R21123 VSS.n2588 VSS.n2435 4.5005
R21124 VSS.n2590 VSS.n2435 4.5005
R21125 VSS.n2593 VSS.n2435 4.5005
R21126 VSS.n2595 VSS.n2435 4.5005
R21127 VSS.n2596 VSS.n2435 4.5005
R21128 VSS.n2598 VSS.n2435 4.5005
R21129 VSS.n2601 VSS.n2435 4.5005
R21130 VSS.n2603 VSS.n2435 4.5005
R21131 VSS.n2604 VSS.n2435 4.5005
R21132 VSS.n2606 VSS.n2435 4.5005
R21133 VSS.n2609 VSS.n2435 4.5005
R21134 VSS.n2611 VSS.n2435 4.5005
R21135 VSS.n2612 VSS.n2435 4.5005
R21136 VSS.n2614 VSS.n2435 4.5005
R21137 VSS.n2617 VSS.n2435 4.5005
R21138 VSS.n2619 VSS.n2435 4.5005
R21139 VSS.n2620 VSS.n2435 4.5005
R21140 VSS.n2622 VSS.n2435 4.5005
R21141 VSS.n2625 VSS.n2435 4.5005
R21142 VSS.n2627 VSS.n2435 4.5005
R21143 VSS.n2628 VSS.n2435 4.5005
R21144 VSS.n2630 VSS.n2435 4.5005
R21145 VSS.n2633 VSS.n2435 4.5005
R21146 VSS.n2635 VSS.n2435 4.5005
R21147 VSS.n2636 VSS.n2435 4.5005
R21148 VSS.n2638 VSS.n2435 4.5005
R21149 VSS.n2640 VSS.n2435 4.5005
R21150 VSS.n2642 VSS.n2435 4.5005
R21151 VSS.n2643 VSS.n2435 4.5005
R21152 VSS.n2645 VSS.n2435 4.5005
R21153 VSS.n2648 VSS.n2435 4.5005
R21154 VSS.n2650 VSS.n2435 4.5005
R21155 VSS.n2651 VSS.n2435 4.5005
R21156 VSS.n2653 VSS.n2435 4.5005
R21157 VSS.n2656 VSS.n2435 4.5005
R21158 VSS.n2658 VSS.n2435 4.5005
R21159 VSS.n2659 VSS.n2435 4.5005
R21160 VSS.n2661 VSS.n2435 4.5005
R21161 VSS.n2664 VSS.n2435 4.5005
R21162 VSS.n2666 VSS.n2435 4.5005
R21163 VSS.n2667 VSS.n2435 4.5005
R21164 VSS.n2669 VSS.n2435 4.5005
R21165 VSS.n2672 VSS.n2435 4.5005
R21166 VSS.n2674 VSS.n2435 4.5005
R21167 VSS.n2675 VSS.n2435 4.5005
R21168 VSS.n2677 VSS.n2435 4.5005
R21169 VSS.n2680 VSS.n2435 4.5005
R21170 VSS.n2682 VSS.n2435 4.5005
R21171 VSS.n2683 VSS.n2435 4.5005
R21172 VSS.n2685 VSS.n2435 4.5005
R21173 VSS.n2688 VSS.n2435 4.5005
R21174 VSS.n2690 VSS.n2435 4.5005
R21175 VSS.n2691 VSS.n2435 4.5005
R21176 VSS.n2693 VSS.n2435 4.5005
R21177 VSS.n2696 VSS.n2435 4.5005
R21178 VSS.n2698 VSS.n2435 4.5005
R21179 VSS.n2699 VSS.n2435 4.5005
R21180 VSS.n2701 VSS.n2435 4.5005
R21181 VSS.n2704 VSS.n2435 4.5005
R21182 VSS.n2706 VSS.n2435 4.5005
R21183 VSS.n2707 VSS.n2435 4.5005
R21184 VSS.n2709 VSS.n2435 4.5005
R21185 VSS.n2712 VSS.n2435 4.5005
R21186 VSS.n2714 VSS.n2435 4.5005
R21187 VSS.n2715 VSS.n2435 4.5005
R21188 VSS.n2717 VSS.n2435 4.5005
R21189 VSS.n2720 VSS.n2435 4.5005
R21190 VSS.n2722 VSS.n2435 4.5005
R21191 VSS.n2723 VSS.n2435 4.5005
R21192 VSS.n2725 VSS.n2435 4.5005
R21193 VSS.n2793 VSS.n2435 4.5005
R21194 VSS.n2859 VSS.n2435 4.5005
R21195 VSS.n3051 VSS.n2396 4.5005
R21196 VSS.n2396 VSS.n2351 4.5005
R21197 VSS.n2483 VSS.n2396 4.5005
R21198 VSS.n2484 VSS.n2396 4.5005
R21199 VSS.n2486 VSS.n2396 4.5005
R21200 VSS.n2489 VSS.n2396 4.5005
R21201 VSS.n2491 VSS.n2396 4.5005
R21202 VSS.n2492 VSS.n2396 4.5005
R21203 VSS.n2494 VSS.n2396 4.5005
R21204 VSS.n2497 VSS.n2396 4.5005
R21205 VSS.n2499 VSS.n2396 4.5005
R21206 VSS.n2500 VSS.n2396 4.5005
R21207 VSS.n2502 VSS.n2396 4.5005
R21208 VSS.n2505 VSS.n2396 4.5005
R21209 VSS.n2507 VSS.n2396 4.5005
R21210 VSS.n2508 VSS.n2396 4.5005
R21211 VSS.n2510 VSS.n2396 4.5005
R21212 VSS.n2513 VSS.n2396 4.5005
R21213 VSS.n2515 VSS.n2396 4.5005
R21214 VSS.n2516 VSS.n2396 4.5005
R21215 VSS.n2518 VSS.n2396 4.5005
R21216 VSS.n2521 VSS.n2396 4.5005
R21217 VSS.n2523 VSS.n2396 4.5005
R21218 VSS.n2524 VSS.n2396 4.5005
R21219 VSS.n2526 VSS.n2396 4.5005
R21220 VSS.n2529 VSS.n2396 4.5005
R21221 VSS.n2531 VSS.n2396 4.5005
R21222 VSS.n2532 VSS.n2396 4.5005
R21223 VSS.n2534 VSS.n2396 4.5005
R21224 VSS.n2537 VSS.n2396 4.5005
R21225 VSS.n2539 VSS.n2396 4.5005
R21226 VSS.n2540 VSS.n2396 4.5005
R21227 VSS.n2542 VSS.n2396 4.5005
R21228 VSS.n2545 VSS.n2396 4.5005
R21229 VSS.n2547 VSS.n2396 4.5005
R21230 VSS.n2548 VSS.n2396 4.5005
R21231 VSS.n2550 VSS.n2396 4.5005
R21232 VSS.n2553 VSS.n2396 4.5005
R21233 VSS.n2555 VSS.n2396 4.5005
R21234 VSS.n2556 VSS.n2396 4.5005
R21235 VSS.n2558 VSS.n2396 4.5005
R21236 VSS.n2561 VSS.n2396 4.5005
R21237 VSS.n2563 VSS.n2396 4.5005
R21238 VSS.n2564 VSS.n2396 4.5005
R21239 VSS.n2566 VSS.n2396 4.5005
R21240 VSS.n2569 VSS.n2396 4.5005
R21241 VSS.n2571 VSS.n2396 4.5005
R21242 VSS.n2572 VSS.n2396 4.5005
R21243 VSS.n2574 VSS.n2396 4.5005
R21244 VSS.n2577 VSS.n2396 4.5005
R21245 VSS.n2579 VSS.n2396 4.5005
R21246 VSS.n2580 VSS.n2396 4.5005
R21247 VSS.n2582 VSS.n2396 4.5005
R21248 VSS.n2585 VSS.n2396 4.5005
R21249 VSS.n2587 VSS.n2396 4.5005
R21250 VSS.n2588 VSS.n2396 4.5005
R21251 VSS.n2590 VSS.n2396 4.5005
R21252 VSS.n2593 VSS.n2396 4.5005
R21253 VSS.n2595 VSS.n2396 4.5005
R21254 VSS.n2596 VSS.n2396 4.5005
R21255 VSS.n2598 VSS.n2396 4.5005
R21256 VSS.n2601 VSS.n2396 4.5005
R21257 VSS.n2603 VSS.n2396 4.5005
R21258 VSS.n2604 VSS.n2396 4.5005
R21259 VSS.n2606 VSS.n2396 4.5005
R21260 VSS.n2609 VSS.n2396 4.5005
R21261 VSS.n2611 VSS.n2396 4.5005
R21262 VSS.n2612 VSS.n2396 4.5005
R21263 VSS.n2614 VSS.n2396 4.5005
R21264 VSS.n2617 VSS.n2396 4.5005
R21265 VSS.n2619 VSS.n2396 4.5005
R21266 VSS.n2620 VSS.n2396 4.5005
R21267 VSS.n2622 VSS.n2396 4.5005
R21268 VSS.n2625 VSS.n2396 4.5005
R21269 VSS.n2627 VSS.n2396 4.5005
R21270 VSS.n2628 VSS.n2396 4.5005
R21271 VSS.n2630 VSS.n2396 4.5005
R21272 VSS.n2633 VSS.n2396 4.5005
R21273 VSS.n2635 VSS.n2396 4.5005
R21274 VSS.n2636 VSS.n2396 4.5005
R21275 VSS.n2638 VSS.n2396 4.5005
R21276 VSS.n2640 VSS.n2396 4.5005
R21277 VSS.n2642 VSS.n2396 4.5005
R21278 VSS.n2643 VSS.n2396 4.5005
R21279 VSS.n2645 VSS.n2396 4.5005
R21280 VSS.n2648 VSS.n2396 4.5005
R21281 VSS.n2650 VSS.n2396 4.5005
R21282 VSS.n2651 VSS.n2396 4.5005
R21283 VSS.n2653 VSS.n2396 4.5005
R21284 VSS.n2656 VSS.n2396 4.5005
R21285 VSS.n2658 VSS.n2396 4.5005
R21286 VSS.n2659 VSS.n2396 4.5005
R21287 VSS.n2661 VSS.n2396 4.5005
R21288 VSS.n2664 VSS.n2396 4.5005
R21289 VSS.n2666 VSS.n2396 4.5005
R21290 VSS.n2667 VSS.n2396 4.5005
R21291 VSS.n2669 VSS.n2396 4.5005
R21292 VSS.n2672 VSS.n2396 4.5005
R21293 VSS.n2674 VSS.n2396 4.5005
R21294 VSS.n2675 VSS.n2396 4.5005
R21295 VSS.n2677 VSS.n2396 4.5005
R21296 VSS.n2680 VSS.n2396 4.5005
R21297 VSS.n2682 VSS.n2396 4.5005
R21298 VSS.n2683 VSS.n2396 4.5005
R21299 VSS.n2685 VSS.n2396 4.5005
R21300 VSS.n2688 VSS.n2396 4.5005
R21301 VSS.n2690 VSS.n2396 4.5005
R21302 VSS.n2691 VSS.n2396 4.5005
R21303 VSS.n2693 VSS.n2396 4.5005
R21304 VSS.n2696 VSS.n2396 4.5005
R21305 VSS.n2698 VSS.n2396 4.5005
R21306 VSS.n2699 VSS.n2396 4.5005
R21307 VSS.n2701 VSS.n2396 4.5005
R21308 VSS.n2704 VSS.n2396 4.5005
R21309 VSS.n2706 VSS.n2396 4.5005
R21310 VSS.n2707 VSS.n2396 4.5005
R21311 VSS.n2709 VSS.n2396 4.5005
R21312 VSS.n2712 VSS.n2396 4.5005
R21313 VSS.n2714 VSS.n2396 4.5005
R21314 VSS.n2715 VSS.n2396 4.5005
R21315 VSS.n2717 VSS.n2396 4.5005
R21316 VSS.n2720 VSS.n2396 4.5005
R21317 VSS.n2722 VSS.n2396 4.5005
R21318 VSS.n2723 VSS.n2396 4.5005
R21319 VSS.n2725 VSS.n2396 4.5005
R21320 VSS.n2793 VSS.n2396 4.5005
R21321 VSS.n2859 VSS.n2396 4.5005
R21322 VSS.n3051 VSS.n2436 4.5005
R21323 VSS.n2436 VSS.n2351 4.5005
R21324 VSS.n2483 VSS.n2436 4.5005
R21325 VSS.n2484 VSS.n2436 4.5005
R21326 VSS.n2486 VSS.n2436 4.5005
R21327 VSS.n2489 VSS.n2436 4.5005
R21328 VSS.n2491 VSS.n2436 4.5005
R21329 VSS.n2492 VSS.n2436 4.5005
R21330 VSS.n2494 VSS.n2436 4.5005
R21331 VSS.n2497 VSS.n2436 4.5005
R21332 VSS.n2499 VSS.n2436 4.5005
R21333 VSS.n2500 VSS.n2436 4.5005
R21334 VSS.n2502 VSS.n2436 4.5005
R21335 VSS.n2505 VSS.n2436 4.5005
R21336 VSS.n2507 VSS.n2436 4.5005
R21337 VSS.n2508 VSS.n2436 4.5005
R21338 VSS.n2510 VSS.n2436 4.5005
R21339 VSS.n2513 VSS.n2436 4.5005
R21340 VSS.n2515 VSS.n2436 4.5005
R21341 VSS.n2516 VSS.n2436 4.5005
R21342 VSS.n2518 VSS.n2436 4.5005
R21343 VSS.n2521 VSS.n2436 4.5005
R21344 VSS.n2523 VSS.n2436 4.5005
R21345 VSS.n2524 VSS.n2436 4.5005
R21346 VSS.n2526 VSS.n2436 4.5005
R21347 VSS.n2529 VSS.n2436 4.5005
R21348 VSS.n2531 VSS.n2436 4.5005
R21349 VSS.n2532 VSS.n2436 4.5005
R21350 VSS.n2534 VSS.n2436 4.5005
R21351 VSS.n2537 VSS.n2436 4.5005
R21352 VSS.n2539 VSS.n2436 4.5005
R21353 VSS.n2540 VSS.n2436 4.5005
R21354 VSS.n2542 VSS.n2436 4.5005
R21355 VSS.n2545 VSS.n2436 4.5005
R21356 VSS.n2547 VSS.n2436 4.5005
R21357 VSS.n2548 VSS.n2436 4.5005
R21358 VSS.n2550 VSS.n2436 4.5005
R21359 VSS.n2553 VSS.n2436 4.5005
R21360 VSS.n2555 VSS.n2436 4.5005
R21361 VSS.n2556 VSS.n2436 4.5005
R21362 VSS.n2558 VSS.n2436 4.5005
R21363 VSS.n2561 VSS.n2436 4.5005
R21364 VSS.n2563 VSS.n2436 4.5005
R21365 VSS.n2564 VSS.n2436 4.5005
R21366 VSS.n2566 VSS.n2436 4.5005
R21367 VSS.n2569 VSS.n2436 4.5005
R21368 VSS.n2571 VSS.n2436 4.5005
R21369 VSS.n2572 VSS.n2436 4.5005
R21370 VSS.n2574 VSS.n2436 4.5005
R21371 VSS.n2577 VSS.n2436 4.5005
R21372 VSS.n2579 VSS.n2436 4.5005
R21373 VSS.n2580 VSS.n2436 4.5005
R21374 VSS.n2582 VSS.n2436 4.5005
R21375 VSS.n2585 VSS.n2436 4.5005
R21376 VSS.n2587 VSS.n2436 4.5005
R21377 VSS.n2588 VSS.n2436 4.5005
R21378 VSS.n2590 VSS.n2436 4.5005
R21379 VSS.n2593 VSS.n2436 4.5005
R21380 VSS.n2595 VSS.n2436 4.5005
R21381 VSS.n2596 VSS.n2436 4.5005
R21382 VSS.n2598 VSS.n2436 4.5005
R21383 VSS.n2601 VSS.n2436 4.5005
R21384 VSS.n2603 VSS.n2436 4.5005
R21385 VSS.n2604 VSS.n2436 4.5005
R21386 VSS.n2606 VSS.n2436 4.5005
R21387 VSS.n2609 VSS.n2436 4.5005
R21388 VSS.n2611 VSS.n2436 4.5005
R21389 VSS.n2612 VSS.n2436 4.5005
R21390 VSS.n2614 VSS.n2436 4.5005
R21391 VSS.n2617 VSS.n2436 4.5005
R21392 VSS.n2619 VSS.n2436 4.5005
R21393 VSS.n2620 VSS.n2436 4.5005
R21394 VSS.n2622 VSS.n2436 4.5005
R21395 VSS.n2625 VSS.n2436 4.5005
R21396 VSS.n2627 VSS.n2436 4.5005
R21397 VSS.n2628 VSS.n2436 4.5005
R21398 VSS.n2630 VSS.n2436 4.5005
R21399 VSS.n2633 VSS.n2436 4.5005
R21400 VSS.n2635 VSS.n2436 4.5005
R21401 VSS.n2636 VSS.n2436 4.5005
R21402 VSS.n2638 VSS.n2436 4.5005
R21403 VSS.n2640 VSS.n2436 4.5005
R21404 VSS.n2642 VSS.n2436 4.5005
R21405 VSS.n2643 VSS.n2436 4.5005
R21406 VSS.n2645 VSS.n2436 4.5005
R21407 VSS.n2648 VSS.n2436 4.5005
R21408 VSS.n2650 VSS.n2436 4.5005
R21409 VSS.n2651 VSS.n2436 4.5005
R21410 VSS.n2653 VSS.n2436 4.5005
R21411 VSS.n2656 VSS.n2436 4.5005
R21412 VSS.n2658 VSS.n2436 4.5005
R21413 VSS.n2659 VSS.n2436 4.5005
R21414 VSS.n2661 VSS.n2436 4.5005
R21415 VSS.n2664 VSS.n2436 4.5005
R21416 VSS.n2666 VSS.n2436 4.5005
R21417 VSS.n2667 VSS.n2436 4.5005
R21418 VSS.n2669 VSS.n2436 4.5005
R21419 VSS.n2672 VSS.n2436 4.5005
R21420 VSS.n2674 VSS.n2436 4.5005
R21421 VSS.n2675 VSS.n2436 4.5005
R21422 VSS.n2677 VSS.n2436 4.5005
R21423 VSS.n2680 VSS.n2436 4.5005
R21424 VSS.n2682 VSS.n2436 4.5005
R21425 VSS.n2683 VSS.n2436 4.5005
R21426 VSS.n2685 VSS.n2436 4.5005
R21427 VSS.n2688 VSS.n2436 4.5005
R21428 VSS.n2690 VSS.n2436 4.5005
R21429 VSS.n2691 VSS.n2436 4.5005
R21430 VSS.n2693 VSS.n2436 4.5005
R21431 VSS.n2696 VSS.n2436 4.5005
R21432 VSS.n2698 VSS.n2436 4.5005
R21433 VSS.n2699 VSS.n2436 4.5005
R21434 VSS.n2701 VSS.n2436 4.5005
R21435 VSS.n2704 VSS.n2436 4.5005
R21436 VSS.n2706 VSS.n2436 4.5005
R21437 VSS.n2707 VSS.n2436 4.5005
R21438 VSS.n2709 VSS.n2436 4.5005
R21439 VSS.n2712 VSS.n2436 4.5005
R21440 VSS.n2714 VSS.n2436 4.5005
R21441 VSS.n2715 VSS.n2436 4.5005
R21442 VSS.n2717 VSS.n2436 4.5005
R21443 VSS.n2720 VSS.n2436 4.5005
R21444 VSS.n2722 VSS.n2436 4.5005
R21445 VSS.n2723 VSS.n2436 4.5005
R21446 VSS.n2725 VSS.n2436 4.5005
R21447 VSS.n2793 VSS.n2436 4.5005
R21448 VSS.n2859 VSS.n2436 4.5005
R21449 VSS.n3051 VSS.n2395 4.5005
R21450 VSS.n2395 VSS.n2351 4.5005
R21451 VSS.n2483 VSS.n2395 4.5005
R21452 VSS.n2484 VSS.n2395 4.5005
R21453 VSS.n2486 VSS.n2395 4.5005
R21454 VSS.n2489 VSS.n2395 4.5005
R21455 VSS.n2491 VSS.n2395 4.5005
R21456 VSS.n2492 VSS.n2395 4.5005
R21457 VSS.n2494 VSS.n2395 4.5005
R21458 VSS.n2497 VSS.n2395 4.5005
R21459 VSS.n2499 VSS.n2395 4.5005
R21460 VSS.n2500 VSS.n2395 4.5005
R21461 VSS.n2502 VSS.n2395 4.5005
R21462 VSS.n2505 VSS.n2395 4.5005
R21463 VSS.n2507 VSS.n2395 4.5005
R21464 VSS.n2508 VSS.n2395 4.5005
R21465 VSS.n2510 VSS.n2395 4.5005
R21466 VSS.n2513 VSS.n2395 4.5005
R21467 VSS.n2515 VSS.n2395 4.5005
R21468 VSS.n2516 VSS.n2395 4.5005
R21469 VSS.n2518 VSS.n2395 4.5005
R21470 VSS.n2521 VSS.n2395 4.5005
R21471 VSS.n2523 VSS.n2395 4.5005
R21472 VSS.n2524 VSS.n2395 4.5005
R21473 VSS.n2526 VSS.n2395 4.5005
R21474 VSS.n2529 VSS.n2395 4.5005
R21475 VSS.n2531 VSS.n2395 4.5005
R21476 VSS.n2532 VSS.n2395 4.5005
R21477 VSS.n2534 VSS.n2395 4.5005
R21478 VSS.n2537 VSS.n2395 4.5005
R21479 VSS.n2539 VSS.n2395 4.5005
R21480 VSS.n2540 VSS.n2395 4.5005
R21481 VSS.n2542 VSS.n2395 4.5005
R21482 VSS.n2545 VSS.n2395 4.5005
R21483 VSS.n2547 VSS.n2395 4.5005
R21484 VSS.n2548 VSS.n2395 4.5005
R21485 VSS.n2550 VSS.n2395 4.5005
R21486 VSS.n2553 VSS.n2395 4.5005
R21487 VSS.n2555 VSS.n2395 4.5005
R21488 VSS.n2556 VSS.n2395 4.5005
R21489 VSS.n2558 VSS.n2395 4.5005
R21490 VSS.n2561 VSS.n2395 4.5005
R21491 VSS.n2563 VSS.n2395 4.5005
R21492 VSS.n2564 VSS.n2395 4.5005
R21493 VSS.n2566 VSS.n2395 4.5005
R21494 VSS.n2569 VSS.n2395 4.5005
R21495 VSS.n2571 VSS.n2395 4.5005
R21496 VSS.n2572 VSS.n2395 4.5005
R21497 VSS.n2574 VSS.n2395 4.5005
R21498 VSS.n2577 VSS.n2395 4.5005
R21499 VSS.n2579 VSS.n2395 4.5005
R21500 VSS.n2580 VSS.n2395 4.5005
R21501 VSS.n2582 VSS.n2395 4.5005
R21502 VSS.n2585 VSS.n2395 4.5005
R21503 VSS.n2587 VSS.n2395 4.5005
R21504 VSS.n2588 VSS.n2395 4.5005
R21505 VSS.n2590 VSS.n2395 4.5005
R21506 VSS.n2593 VSS.n2395 4.5005
R21507 VSS.n2595 VSS.n2395 4.5005
R21508 VSS.n2596 VSS.n2395 4.5005
R21509 VSS.n2598 VSS.n2395 4.5005
R21510 VSS.n2601 VSS.n2395 4.5005
R21511 VSS.n2603 VSS.n2395 4.5005
R21512 VSS.n2604 VSS.n2395 4.5005
R21513 VSS.n2606 VSS.n2395 4.5005
R21514 VSS.n2609 VSS.n2395 4.5005
R21515 VSS.n2611 VSS.n2395 4.5005
R21516 VSS.n2612 VSS.n2395 4.5005
R21517 VSS.n2614 VSS.n2395 4.5005
R21518 VSS.n2617 VSS.n2395 4.5005
R21519 VSS.n2619 VSS.n2395 4.5005
R21520 VSS.n2620 VSS.n2395 4.5005
R21521 VSS.n2622 VSS.n2395 4.5005
R21522 VSS.n2625 VSS.n2395 4.5005
R21523 VSS.n2627 VSS.n2395 4.5005
R21524 VSS.n2628 VSS.n2395 4.5005
R21525 VSS.n2630 VSS.n2395 4.5005
R21526 VSS.n2633 VSS.n2395 4.5005
R21527 VSS.n2635 VSS.n2395 4.5005
R21528 VSS.n2636 VSS.n2395 4.5005
R21529 VSS.n2638 VSS.n2395 4.5005
R21530 VSS.n2640 VSS.n2395 4.5005
R21531 VSS.n2642 VSS.n2395 4.5005
R21532 VSS.n2643 VSS.n2395 4.5005
R21533 VSS.n2645 VSS.n2395 4.5005
R21534 VSS.n2648 VSS.n2395 4.5005
R21535 VSS.n2650 VSS.n2395 4.5005
R21536 VSS.n2651 VSS.n2395 4.5005
R21537 VSS.n2653 VSS.n2395 4.5005
R21538 VSS.n2656 VSS.n2395 4.5005
R21539 VSS.n2658 VSS.n2395 4.5005
R21540 VSS.n2659 VSS.n2395 4.5005
R21541 VSS.n2661 VSS.n2395 4.5005
R21542 VSS.n2664 VSS.n2395 4.5005
R21543 VSS.n2666 VSS.n2395 4.5005
R21544 VSS.n2667 VSS.n2395 4.5005
R21545 VSS.n2669 VSS.n2395 4.5005
R21546 VSS.n2672 VSS.n2395 4.5005
R21547 VSS.n2674 VSS.n2395 4.5005
R21548 VSS.n2675 VSS.n2395 4.5005
R21549 VSS.n2677 VSS.n2395 4.5005
R21550 VSS.n2680 VSS.n2395 4.5005
R21551 VSS.n2682 VSS.n2395 4.5005
R21552 VSS.n2683 VSS.n2395 4.5005
R21553 VSS.n2685 VSS.n2395 4.5005
R21554 VSS.n2688 VSS.n2395 4.5005
R21555 VSS.n2690 VSS.n2395 4.5005
R21556 VSS.n2691 VSS.n2395 4.5005
R21557 VSS.n2693 VSS.n2395 4.5005
R21558 VSS.n2696 VSS.n2395 4.5005
R21559 VSS.n2698 VSS.n2395 4.5005
R21560 VSS.n2699 VSS.n2395 4.5005
R21561 VSS.n2701 VSS.n2395 4.5005
R21562 VSS.n2704 VSS.n2395 4.5005
R21563 VSS.n2706 VSS.n2395 4.5005
R21564 VSS.n2707 VSS.n2395 4.5005
R21565 VSS.n2709 VSS.n2395 4.5005
R21566 VSS.n2712 VSS.n2395 4.5005
R21567 VSS.n2714 VSS.n2395 4.5005
R21568 VSS.n2715 VSS.n2395 4.5005
R21569 VSS.n2717 VSS.n2395 4.5005
R21570 VSS.n2720 VSS.n2395 4.5005
R21571 VSS.n2722 VSS.n2395 4.5005
R21572 VSS.n2723 VSS.n2395 4.5005
R21573 VSS.n2725 VSS.n2395 4.5005
R21574 VSS.n2793 VSS.n2395 4.5005
R21575 VSS.n2859 VSS.n2395 4.5005
R21576 VSS.n3051 VSS.n2437 4.5005
R21577 VSS.n2437 VSS.n2351 4.5005
R21578 VSS.n2483 VSS.n2437 4.5005
R21579 VSS.n2484 VSS.n2437 4.5005
R21580 VSS.n2486 VSS.n2437 4.5005
R21581 VSS.n2489 VSS.n2437 4.5005
R21582 VSS.n2491 VSS.n2437 4.5005
R21583 VSS.n2492 VSS.n2437 4.5005
R21584 VSS.n2494 VSS.n2437 4.5005
R21585 VSS.n2497 VSS.n2437 4.5005
R21586 VSS.n2499 VSS.n2437 4.5005
R21587 VSS.n2500 VSS.n2437 4.5005
R21588 VSS.n2502 VSS.n2437 4.5005
R21589 VSS.n2505 VSS.n2437 4.5005
R21590 VSS.n2507 VSS.n2437 4.5005
R21591 VSS.n2508 VSS.n2437 4.5005
R21592 VSS.n2510 VSS.n2437 4.5005
R21593 VSS.n2513 VSS.n2437 4.5005
R21594 VSS.n2515 VSS.n2437 4.5005
R21595 VSS.n2516 VSS.n2437 4.5005
R21596 VSS.n2518 VSS.n2437 4.5005
R21597 VSS.n2521 VSS.n2437 4.5005
R21598 VSS.n2523 VSS.n2437 4.5005
R21599 VSS.n2524 VSS.n2437 4.5005
R21600 VSS.n2526 VSS.n2437 4.5005
R21601 VSS.n2529 VSS.n2437 4.5005
R21602 VSS.n2531 VSS.n2437 4.5005
R21603 VSS.n2532 VSS.n2437 4.5005
R21604 VSS.n2534 VSS.n2437 4.5005
R21605 VSS.n2537 VSS.n2437 4.5005
R21606 VSS.n2539 VSS.n2437 4.5005
R21607 VSS.n2540 VSS.n2437 4.5005
R21608 VSS.n2542 VSS.n2437 4.5005
R21609 VSS.n2545 VSS.n2437 4.5005
R21610 VSS.n2547 VSS.n2437 4.5005
R21611 VSS.n2548 VSS.n2437 4.5005
R21612 VSS.n2550 VSS.n2437 4.5005
R21613 VSS.n2553 VSS.n2437 4.5005
R21614 VSS.n2555 VSS.n2437 4.5005
R21615 VSS.n2556 VSS.n2437 4.5005
R21616 VSS.n2558 VSS.n2437 4.5005
R21617 VSS.n2561 VSS.n2437 4.5005
R21618 VSS.n2563 VSS.n2437 4.5005
R21619 VSS.n2564 VSS.n2437 4.5005
R21620 VSS.n2566 VSS.n2437 4.5005
R21621 VSS.n2569 VSS.n2437 4.5005
R21622 VSS.n2571 VSS.n2437 4.5005
R21623 VSS.n2572 VSS.n2437 4.5005
R21624 VSS.n2574 VSS.n2437 4.5005
R21625 VSS.n2577 VSS.n2437 4.5005
R21626 VSS.n2579 VSS.n2437 4.5005
R21627 VSS.n2580 VSS.n2437 4.5005
R21628 VSS.n2582 VSS.n2437 4.5005
R21629 VSS.n2585 VSS.n2437 4.5005
R21630 VSS.n2587 VSS.n2437 4.5005
R21631 VSS.n2588 VSS.n2437 4.5005
R21632 VSS.n2590 VSS.n2437 4.5005
R21633 VSS.n2593 VSS.n2437 4.5005
R21634 VSS.n2595 VSS.n2437 4.5005
R21635 VSS.n2596 VSS.n2437 4.5005
R21636 VSS.n2598 VSS.n2437 4.5005
R21637 VSS.n2601 VSS.n2437 4.5005
R21638 VSS.n2603 VSS.n2437 4.5005
R21639 VSS.n2604 VSS.n2437 4.5005
R21640 VSS.n2606 VSS.n2437 4.5005
R21641 VSS.n2609 VSS.n2437 4.5005
R21642 VSS.n2611 VSS.n2437 4.5005
R21643 VSS.n2612 VSS.n2437 4.5005
R21644 VSS.n2614 VSS.n2437 4.5005
R21645 VSS.n2617 VSS.n2437 4.5005
R21646 VSS.n2619 VSS.n2437 4.5005
R21647 VSS.n2620 VSS.n2437 4.5005
R21648 VSS.n2622 VSS.n2437 4.5005
R21649 VSS.n2625 VSS.n2437 4.5005
R21650 VSS.n2627 VSS.n2437 4.5005
R21651 VSS.n2628 VSS.n2437 4.5005
R21652 VSS.n2630 VSS.n2437 4.5005
R21653 VSS.n2633 VSS.n2437 4.5005
R21654 VSS.n2635 VSS.n2437 4.5005
R21655 VSS.n2636 VSS.n2437 4.5005
R21656 VSS.n2638 VSS.n2437 4.5005
R21657 VSS.n2640 VSS.n2437 4.5005
R21658 VSS.n2642 VSS.n2437 4.5005
R21659 VSS.n2643 VSS.n2437 4.5005
R21660 VSS.n2645 VSS.n2437 4.5005
R21661 VSS.n2648 VSS.n2437 4.5005
R21662 VSS.n2650 VSS.n2437 4.5005
R21663 VSS.n2651 VSS.n2437 4.5005
R21664 VSS.n2653 VSS.n2437 4.5005
R21665 VSS.n2656 VSS.n2437 4.5005
R21666 VSS.n2658 VSS.n2437 4.5005
R21667 VSS.n2659 VSS.n2437 4.5005
R21668 VSS.n2661 VSS.n2437 4.5005
R21669 VSS.n2664 VSS.n2437 4.5005
R21670 VSS.n2666 VSS.n2437 4.5005
R21671 VSS.n2667 VSS.n2437 4.5005
R21672 VSS.n2669 VSS.n2437 4.5005
R21673 VSS.n2672 VSS.n2437 4.5005
R21674 VSS.n2674 VSS.n2437 4.5005
R21675 VSS.n2675 VSS.n2437 4.5005
R21676 VSS.n2677 VSS.n2437 4.5005
R21677 VSS.n2680 VSS.n2437 4.5005
R21678 VSS.n2682 VSS.n2437 4.5005
R21679 VSS.n2683 VSS.n2437 4.5005
R21680 VSS.n2685 VSS.n2437 4.5005
R21681 VSS.n2688 VSS.n2437 4.5005
R21682 VSS.n2690 VSS.n2437 4.5005
R21683 VSS.n2691 VSS.n2437 4.5005
R21684 VSS.n2693 VSS.n2437 4.5005
R21685 VSS.n2696 VSS.n2437 4.5005
R21686 VSS.n2698 VSS.n2437 4.5005
R21687 VSS.n2699 VSS.n2437 4.5005
R21688 VSS.n2701 VSS.n2437 4.5005
R21689 VSS.n2704 VSS.n2437 4.5005
R21690 VSS.n2706 VSS.n2437 4.5005
R21691 VSS.n2707 VSS.n2437 4.5005
R21692 VSS.n2709 VSS.n2437 4.5005
R21693 VSS.n2712 VSS.n2437 4.5005
R21694 VSS.n2714 VSS.n2437 4.5005
R21695 VSS.n2715 VSS.n2437 4.5005
R21696 VSS.n2717 VSS.n2437 4.5005
R21697 VSS.n2720 VSS.n2437 4.5005
R21698 VSS.n2722 VSS.n2437 4.5005
R21699 VSS.n2723 VSS.n2437 4.5005
R21700 VSS.n2725 VSS.n2437 4.5005
R21701 VSS.n2793 VSS.n2437 4.5005
R21702 VSS.n2859 VSS.n2437 4.5005
R21703 VSS.n3051 VSS.n2394 4.5005
R21704 VSS.n2394 VSS.n2351 4.5005
R21705 VSS.n2483 VSS.n2394 4.5005
R21706 VSS.n2484 VSS.n2394 4.5005
R21707 VSS.n2486 VSS.n2394 4.5005
R21708 VSS.n2489 VSS.n2394 4.5005
R21709 VSS.n2491 VSS.n2394 4.5005
R21710 VSS.n2492 VSS.n2394 4.5005
R21711 VSS.n2494 VSS.n2394 4.5005
R21712 VSS.n2497 VSS.n2394 4.5005
R21713 VSS.n2499 VSS.n2394 4.5005
R21714 VSS.n2500 VSS.n2394 4.5005
R21715 VSS.n2502 VSS.n2394 4.5005
R21716 VSS.n2505 VSS.n2394 4.5005
R21717 VSS.n2507 VSS.n2394 4.5005
R21718 VSS.n2508 VSS.n2394 4.5005
R21719 VSS.n2510 VSS.n2394 4.5005
R21720 VSS.n2513 VSS.n2394 4.5005
R21721 VSS.n2515 VSS.n2394 4.5005
R21722 VSS.n2516 VSS.n2394 4.5005
R21723 VSS.n2518 VSS.n2394 4.5005
R21724 VSS.n2521 VSS.n2394 4.5005
R21725 VSS.n2523 VSS.n2394 4.5005
R21726 VSS.n2524 VSS.n2394 4.5005
R21727 VSS.n2526 VSS.n2394 4.5005
R21728 VSS.n2529 VSS.n2394 4.5005
R21729 VSS.n2531 VSS.n2394 4.5005
R21730 VSS.n2532 VSS.n2394 4.5005
R21731 VSS.n2534 VSS.n2394 4.5005
R21732 VSS.n2537 VSS.n2394 4.5005
R21733 VSS.n2539 VSS.n2394 4.5005
R21734 VSS.n2540 VSS.n2394 4.5005
R21735 VSS.n2542 VSS.n2394 4.5005
R21736 VSS.n2545 VSS.n2394 4.5005
R21737 VSS.n2547 VSS.n2394 4.5005
R21738 VSS.n2548 VSS.n2394 4.5005
R21739 VSS.n2550 VSS.n2394 4.5005
R21740 VSS.n2553 VSS.n2394 4.5005
R21741 VSS.n2555 VSS.n2394 4.5005
R21742 VSS.n2556 VSS.n2394 4.5005
R21743 VSS.n2558 VSS.n2394 4.5005
R21744 VSS.n2561 VSS.n2394 4.5005
R21745 VSS.n2563 VSS.n2394 4.5005
R21746 VSS.n2564 VSS.n2394 4.5005
R21747 VSS.n2566 VSS.n2394 4.5005
R21748 VSS.n2569 VSS.n2394 4.5005
R21749 VSS.n2571 VSS.n2394 4.5005
R21750 VSS.n2572 VSS.n2394 4.5005
R21751 VSS.n2574 VSS.n2394 4.5005
R21752 VSS.n2577 VSS.n2394 4.5005
R21753 VSS.n2579 VSS.n2394 4.5005
R21754 VSS.n2580 VSS.n2394 4.5005
R21755 VSS.n2582 VSS.n2394 4.5005
R21756 VSS.n2585 VSS.n2394 4.5005
R21757 VSS.n2587 VSS.n2394 4.5005
R21758 VSS.n2588 VSS.n2394 4.5005
R21759 VSS.n2590 VSS.n2394 4.5005
R21760 VSS.n2593 VSS.n2394 4.5005
R21761 VSS.n2595 VSS.n2394 4.5005
R21762 VSS.n2596 VSS.n2394 4.5005
R21763 VSS.n2598 VSS.n2394 4.5005
R21764 VSS.n2601 VSS.n2394 4.5005
R21765 VSS.n2603 VSS.n2394 4.5005
R21766 VSS.n2604 VSS.n2394 4.5005
R21767 VSS.n2606 VSS.n2394 4.5005
R21768 VSS.n2609 VSS.n2394 4.5005
R21769 VSS.n2611 VSS.n2394 4.5005
R21770 VSS.n2612 VSS.n2394 4.5005
R21771 VSS.n2614 VSS.n2394 4.5005
R21772 VSS.n2617 VSS.n2394 4.5005
R21773 VSS.n2619 VSS.n2394 4.5005
R21774 VSS.n2620 VSS.n2394 4.5005
R21775 VSS.n2622 VSS.n2394 4.5005
R21776 VSS.n2625 VSS.n2394 4.5005
R21777 VSS.n2627 VSS.n2394 4.5005
R21778 VSS.n2628 VSS.n2394 4.5005
R21779 VSS.n2630 VSS.n2394 4.5005
R21780 VSS.n2633 VSS.n2394 4.5005
R21781 VSS.n2635 VSS.n2394 4.5005
R21782 VSS.n2636 VSS.n2394 4.5005
R21783 VSS.n2638 VSS.n2394 4.5005
R21784 VSS.n2640 VSS.n2394 4.5005
R21785 VSS.n2642 VSS.n2394 4.5005
R21786 VSS.n2643 VSS.n2394 4.5005
R21787 VSS.n2645 VSS.n2394 4.5005
R21788 VSS.n2648 VSS.n2394 4.5005
R21789 VSS.n2650 VSS.n2394 4.5005
R21790 VSS.n2651 VSS.n2394 4.5005
R21791 VSS.n2653 VSS.n2394 4.5005
R21792 VSS.n2656 VSS.n2394 4.5005
R21793 VSS.n2658 VSS.n2394 4.5005
R21794 VSS.n2659 VSS.n2394 4.5005
R21795 VSS.n2661 VSS.n2394 4.5005
R21796 VSS.n2664 VSS.n2394 4.5005
R21797 VSS.n2666 VSS.n2394 4.5005
R21798 VSS.n2667 VSS.n2394 4.5005
R21799 VSS.n2669 VSS.n2394 4.5005
R21800 VSS.n2672 VSS.n2394 4.5005
R21801 VSS.n2674 VSS.n2394 4.5005
R21802 VSS.n2675 VSS.n2394 4.5005
R21803 VSS.n2677 VSS.n2394 4.5005
R21804 VSS.n2680 VSS.n2394 4.5005
R21805 VSS.n2682 VSS.n2394 4.5005
R21806 VSS.n2683 VSS.n2394 4.5005
R21807 VSS.n2685 VSS.n2394 4.5005
R21808 VSS.n2688 VSS.n2394 4.5005
R21809 VSS.n2690 VSS.n2394 4.5005
R21810 VSS.n2691 VSS.n2394 4.5005
R21811 VSS.n2693 VSS.n2394 4.5005
R21812 VSS.n2696 VSS.n2394 4.5005
R21813 VSS.n2698 VSS.n2394 4.5005
R21814 VSS.n2699 VSS.n2394 4.5005
R21815 VSS.n2701 VSS.n2394 4.5005
R21816 VSS.n2704 VSS.n2394 4.5005
R21817 VSS.n2706 VSS.n2394 4.5005
R21818 VSS.n2707 VSS.n2394 4.5005
R21819 VSS.n2709 VSS.n2394 4.5005
R21820 VSS.n2712 VSS.n2394 4.5005
R21821 VSS.n2714 VSS.n2394 4.5005
R21822 VSS.n2715 VSS.n2394 4.5005
R21823 VSS.n2717 VSS.n2394 4.5005
R21824 VSS.n2720 VSS.n2394 4.5005
R21825 VSS.n2722 VSS.n2394 4.5005
R21826 VSS.n2723 VSS.n2394 4.5005
R21827 VSS.n2725 VSS.n2394 4.5005
R21828 VSS.n2793 VSS.n2394 4.5005
R21829 VSS.n2859 VSS.n2394 4.5005
R21830 VSS.n3051 VSS.n2438 4.5005
R21831 VSS.n2438 VSS.n2351 4.5005
R21832 VSS.n2483 VSS.n2438 4.5005
R21833 VSS.n2484 VSS.n2438 4.5005
R21834 VSS.n2486 VSS.n2438 4.5005
R21835 VSS.n2489 VSS.n2438 4.5005
R21836 VSS.n2491 VSS.n2438 4.5005
R21837 VSS.n2492 VSS.n2438 4.5005
R21838 VSS.n2494 VSS.n2438 4.5005
R21839 VSS.n2497 VSS.n2438 4.5005
R21840 VSS.n2499 VSS.n2438 4.5005
R21841 VSS.n2500 VSS.n2438 4.5005
R21842 VSS.n2502 VSS.n2438 4.5005
R21843 VSS.n2505 VSS.n2438 4.5005
R21844 VSS.n2507 VSS.n2438 4.5005
R21845 VSS.n2508 VSS.n2438 4.5005
R21846 VSS.n2510 VSS.n2438 4.5005
R21847 VSS.n2513 VSS.n2438 4.5005
R21848 VSS.n2515 VSS.n2438 4.5005
R21849 VSS.n2516 VSS.n2438 4.5005
R21850 VSS.n2518 VSS.n2438 4.5005
R21851 VSS.n2521 VSS.n2438 4.5005
R21852 VSS.n2523 VSS.n2438 4.5005
R21853 VSS.n2524 VSS.n2438 4.5005
R21854 VSS.n2526 VSS.n2438 4.5005
R21855 VSS.n2529 VSS.n2438 4.5005
R21856 VSS.n2531 VSS.n2438 4.5005
R21857 VSS.n2532 VSS.n2438 4.5005
R21858 VSS.n2534 VSS.n2438 4.5005
R21859 VSS.n2537 VSS.n2438 4.5005
R21860 VSS.n2539 VSS.n2438 4.5005
R21861 VSS.n2540 VSS.n2438 4.5005
R21862 VSS.n2542 VSS.n2438 4.5005
R21863 VSS.n2545 VSS.n2438 4.5005
R21864 VSS.n2547 VSS.n2438 4.5005
R21865 VSS.n2548 VSS.n2438 4.5005
R21866 VSS.n2550 VSS.n2438 4.5005
R21867 VSS.n2553 VSS.n2438 4.5005
R21868 VSS.n2555 VSS.n2438 4.5005
R21869 VSS.n2556 VSS.n2438 4.5005
R21870 VSS.n2558 VSS.n2438 4.5005
R21871 VSS.n2561 VSS.n2438 4.5005
R21872 VSS.n2563 VSS.n2438 4.5005
R21873 VSS.n2564 VSS.n2438 4.5005
R21874 VSS.n2566 VSS.n2438 4.5005
R21875 VSS.n2569 VSS.n2438 4.5005
R21876 VSS.n2571 VSS.n2438 4.5005
R21877 VSS.n2572 VSS.n2438 4.5005
R21878 VSS.n2574 VSS.n2438 4.5005
R21879 VSS.n2577 VSS.n2438 4.5005
R21880 VSS.n2579 VSS.n2438 4.5005
R21881 VSS.n2580 VSS.n2438 4.5005
R21882 VSS.n2582 VSS.n2438 4.5005
R21883 VSS.n2585 VSS.n2438 4.5005
R21884 VSS.n2587 VSS.n2438 4.5005
R21885 VSS.n2588 VSS.n2438 4.5005
R21886 VSS.n2590 VSS.n2438 4.5005
R21887 VSS.n2593 VSS.n2438 4.5005
R21888 VSS.n2595 VSS.n2438 4.5005
R21889 VSS.n2596 VSS.n2438 4.5005
R21890 VSS.n2598 VSS.n2438 4.5005
R21891 VSS.n2601 VSS.n2438 4.5005
R21892 VSS.n2603 VSS.n2438 4.5005
R21893 VSS.n2604 VSS.n2438 4.5005
R21894 VSS.n2606 VSS.n2438 4.5005
R21895 VSS.n2609 VSS.n2438 4.5005
R21896 VSS.n2611 VSS.n2438 4.5005
R21897 VSS.n2612 VSS.n2438 4.5005
R21898 VSS.n2614 VSS.n2438 4.5005
R21899 VSS.n2617 VSS.n2438 4.5005
R21900 VSS.n2619 VSS.n2438 4.5005
R21901 VSS.n2620 VSS.n2438 4.5005
R21902 VSS.n2622 VSS.n2438 4.5005
R21903 VSS.n2625 VSS.n2438 4.5005
R21904 VSS.n2627 VSS.n2438 4.5005
R21905 VSS.n2628 VSS.n2438 4.5005
R21906 VSS.n2630 VSS.n2438 4.5005
R21907 VSS.n2633 VSS.n2438 4.5005
R21908 VSS.n2635 VSS.n2438 4.5005
R21909 VSS.n2636 VSS.n2438 4.5005
R21910 VSS.n2638 VSS.n2438 4.5005
R21911 VSS.n2640 VSS.n2438 4.5005
R21912 VSS.n2642 VSS.n2438 4.5005
R21913 VSS.n2643 VSS.n2438 4.5005
R21914 VSS.n2645 VSS.n2438 4.5005
R21915 VSS.n2648 VSS.n2438 4.5005
R21916 VSS.n2650 VSS.n2438 4.5005
R21917 VSS.n2651 VSS.n2438 4.5005
R21918 VSS.n2653 VSS.n2438 4.5005
R21919 VSS.n2656 VSS.n2438 4.5005
R21920 VSS.n2658 VSS.n2438 4.5005
R21921 VSS.n2659 VSS.n2438 4.5005
R21922 VSS.n2661 VSS.n2438 4.5005
R21923 VSS.n2664 VSS.n2438 4.5005
R21924 VSS.n2666 VSS.n2438 4.5005
R21925 VSS.n2667 VSS.n2438 4.5005
R21926 VSS.n2669 VSS.n2438 4.5005
R21927 VSS.n2672 VSS.n2438 4.5005
R21928 VSS.n2674 VSS.n2438 4.5005
R21929 VSS.n2675 VSS.n2438 4.5005
R21930 VSS.n2677 VSS.n2438 4.5005
R21931 VSS.n2680 VSS.n2438 4.5005
R21932 VSS.n2682 VSS.n2438 4.5005
R21933 VSS.n2683 VSS.n2438 4.5005
R21934 VSS.n2685 VSS.n2438 4.5005
R21935 VSS.n2688 VSS.n2438 4.5005
R21936 VSS.n2690 VSS.n2438 4.5005
R21937 VSS.n2691 VSS.n2438 4.5005
R21938 VSS.n2693 VSS.n2438 4.5005
R21939 VSS.n2696 VSS.n2438 4.5005
R21940 VSS.n2698 VSS.n2438 4.5005
R21941 VSS.n2699 VSS.n2438 4.5005
R21942 VSS.n2701 VSS.n2438 4.5005
R21943 VSS.n2704 VSS.n2438 4.5005
R21944 VSS.n2706 VSS.n2438 4.5005
R21945 VSS.n2707 VSS.n2438 4.5005
R21946 VSS.n2709 VSS.n2438 4.5005
R21947 VSS.n2712 VSS.n2438 4.5005
R21948 VSS.n2714 VSS.n2438 4.5005
R21949 VSS.n2715 VSS.n2438 4.5005
R21950 VSS.n2717 VSS.n2438 4.5005
R21951 VSS.n2720 VSS.n2438 4.5005
R21952 VSS.n2722 VSS.n2438 4.5005
R21953 VSS.n2723 VSS.n2438 4.5005
R21954 VSS.n2725 VSS.n2438 4.5005
R21955 VSS.n2793 VSS.n2438 4.5005
R21956 VSS.n2859 VSS.n2438 4.5005
R21957 VSS.n3051 VSS.n2393 4.5005
R21958 VSS.n2393 VSS.n2351 4.5005
R21959 VSS.n2483 VSS.n2393 4.5005
R21960 VSS.n2484 VSS.n2393 4.5005
R21961 VSS.n2486 VSS.n2393 4.5005
R21962 VSS.n2489 VSS.n2393 4.5005
R21963 VSS.n2491 VSS.n2393 4.5005
R21964 VSS.n2492 VSS.n2393 4.5005
R21965 VSS.n2494 VSS.n2393 4.5005
R21966 VSS.n2497 VSS.n2393 4.5005
R21967 VSS.n2499 VSS.n2393 4.5005
R21968 VSS.n2500 VSS.n2393 4.5005
R21969 VSS.n2502 VSS.n2393 4.5005
R21970 VSS.n2505 VSS.n2393 4.5005
R21971 VSS.n2507 VSS.n2393 4.5005
R21972 VSS.n2508 VSS.n2393 4.5005
R21973 VSS.n2510 VSS.n2393 4.5005
R21974 VSS.n2513 VSS.n2393 4.5005
R21975 VSS.n2515 VSS.n2393 4.5005
R21976 VSS.n2516 VSS.n2393 4.5005
R21977 VSS.n2518 VSS.n2393 4.5005
R21978 VSS.n2521 VSS.n2393 4.5005
R21979 VSS.n2523 VSS.n2393 4.5005
R21980 VSS.n2524 VSS.n2393 4.5005
R21981 VSS.n2526 VSS.n2393 4.5005
R21982 VSS.n2529 VSS.n2393 4.5005
R21983 VSS.n2531 VSS.n2393 4.5005
R21984 VSS.n2532 VSS.n2393 4.5005
R21985 VSS.n2534 VSS.n2393 4.5005
R21986 VSS.n2537 VSS.n2393 4.5005
R21987 VSS.n2539 VSS.n2393 4.5005
R21988 VSS.n2540 VSS.n2393 4.5005
R21989 VSS.n2542 VSS.n2393 4.5005
R21990 VSS.n2545 VSS.n2393 4.5005
R21991 VSS.n2547 VSS.n2393 4.5005
R21992 VSS.n2548 VSS.n2393 4.5005
R21993 VSS.n2550 VSS.n2393 4.5005
R21994 VSS.n2553 VSS.n2393 4.5005
R21995 VSS.n2555 VSS.n2393 4.5005
R21996 VSS.n2556 VSS.n2393 4.5005
R21997 VSS.n2558 VSS.n2393 4.5005
R21998 VSS.n2561 VSS.n2393 4.5005
R21999 VSS.n2563 VSS.n2393 4.5005
R22000 VSS.n2564 VSS.n2393 4.5005
R22001 VSS.n2566 VSS.n2393 4.5005
R22002 VSS.n2569 VSS.n2393 4.5005
R22003 VSS.n2571 VSS.n2393 4.5005
R22004 VSS.n2572 VSS.n2393 4.5005
R22005 VSS.n2574 VSS.n2393 4.5005
R22006 VSS.n2577 VSS.n2393 4.5005
R22007 VSS.n2579 VSS.n2393 4.5005
R22008 VSS.n2580 VSS.n2393 4.5005
R22009 VSS.n2582 VSS.n2393 4.5005
R22010 VSS.n2585 VSS.n2393 4.5005
R22011 VSS.n2587 VSS.n2393 4.5005
R22012 VSS.n2588 VSS.n2393 4.5005
R22013 VSS.n2590 VSS.n2393 4.5005
R22014 VSS.n2593 VSS.n2393 4.5005
R22015 VSS.n2595 VSS.n2393 4.5005
R22016 VSS.n2596 VSS.n2393 4.5005
R22017 VSS.n2598 VSS.n2393 4.5005
R22018 VSS.n2601 VSS.n2393 4.5005
R22019 VSS.n2603 VSS.n2393 4.5005
R22020 VSS.n2604 VSS.n2393 4.5005
R22021 VSS.n2606 VSS.n2393 4.5005
R22022 VSS.n2609 VSS.n2393 4.5005
R22023 VSS.n2611 VSS.n2393 4.5005
R22024 VSS.n2612 VSS.n2393 4.5005
R22025 VSS.n2614 VSS.n2393 4.5005
R22026 VSS.n2617 VSS.n2393 4.5005
R22027 VSS.n2619 VSS.n2393 4.5005
R22028 VSS.n2620 VSS.n2393 4.5005
R22029 VSS.n2622 VSS.n2393 4.5005
R22030 VSS.n2625 VSS.n2393 4.5005
R22031 VSS.n2627 VSS.n2393 4.5005
R22032 VSS.n2628 VSS.n2393 4.5005
R22033 VSS.n2630 VSS.n2393 4.5005
R22034 VSS.n2633 VSS.n2393 4.5005
R22035 VSS.n2635 VSS.n2393 4.5005
R22036 VSS.n2636 VSS.n2393 4.5005
R22037 VSS.n2638 VSS.n2393 4.5005
R22038 VSS.n2640 VSS.n2393 4.5005
R22039 VSS.n2642 VSS.n2393 4.5005
R22040 VSS.n2643 VSS.n2393 4.5005
R22041 VSS.n2645 VSS.n2393 4.5005
R22042 VSS.n2648 VSS.n2393 4.5005
R22043 VSS.n2650 VSS.n2393 4.5005
R22044 VSS.n2651 VSS.n2393 4.5005
R22045 VSS.n2653 VSS.n2393 4.5005
R22046 VSS.n2656 VSS.n2393 4.5005
R22047 VSS.n2658 VSS.n2393 4.5005
R22048 VSS.n2659 VSS.n2393 4.5005
R22049 VSS.n2661 VSS.n2393 4.5005
R22050 VSS.n2664 VSS.n2393 4.5005
R22051 VSS.n2666 VSS.n2393 4.5005
R22052 VSS.n2667 VSS.n2393 4.5005
R22053 VSS.n2669 VSS.n2393 4.5005
R22054 VSS.n2672 VSS.n2393 4.5005
R22055 VSS.n2674 VSS.n2393 4.5005
R22056 VSS.n2675 VSS.n2393 4.5005
R22057 VSS.n2677 VSS.n2393 4.5005
R22058 VSS.n2680 VSS.n2393 4.5005
R22059 VSS.n2682 VSS.n2393 4.5005
R22060 VSS.n2683 VSS.n2393 4.5005
R22061 VSS.n2685 VSS.n2393 4.5005
R22062 VSS.n2688 VSS.n2393 4.5005
R22063 VSS.n2690 VSS.n2393 4.5005
R22064 VSS.n2691 VSS.n2393 4.5005
R22065 VSS.n2693 VSS.n2393 4.5005
R22066 VSS.n2696 VSS.n2393 4.5005
R22067 VSS.n2698 VSS.n2393 4.5005
R22068 VSS.n2699 VSS.n2393 4.5005
R22069 VSS.n2701 VSS.n2393 4.5005
R22070 VSS.n2704 VSS.n2393 4.5005
R22071 VSS.n2706 VSS.n2393 4.5005
R22072 VSS.n2707 VSS.n2393 4.5005
R22073 VSS.n2709 VSS.n2393 4.5005
R22074 VSS.n2712 VSS.n2393 4.5005
R22075 VSS.n2714 VSS.n2393 4.5005
R22076 VSS.n2715 VSS.n2393 4.5005
R22077 VSS.n2717 VSS.n2393 4.5005
R22078 VSS.n2720 VSS.n2393 4.5005
R22079 VSS.n2722 VSS.n2393 4.5005
R22080 VSS.n2723 VSS.n2393 4.5005
R22081 VSS.n2725 VSS.n2393 4.5005
R22082 VSS.n2793 VSS.n2393 4.5005
R22083 VSS.n2859 VSS.n2393 4.5005
R22084 VSS.n3051 VSS.n2439 4.5005
R22085 VSS.n2439 VSS.n2351 4.5005
R22086 VSS.n2483 VSS.n2439 4.5005
R22087 VSS.n2484 VSS.n2439 4.5005
R22088 VSS.n2486 VSS.n2439 4.5005
R22089 VSS.n2489 VSS.n2439 4.5005
R22090 VSS.n2491 VSS.n2439 4.5005
R22091 VSS.n2492 VSS.n2439 4.5005
R22092 VSS.n2494 VSS.n2439 4.5005
R22093 VSS.n2497 VSS.n2439 4.5005
R22094 VSS.n2499 VSS.n2439 4.5005
R22095 VSS.n2500 VSS.n2439 4.5005
R22096 VSS.n2502 VSS.n2439 4.5005
R22097 VSS.n2505 VSS.n2439 4.5005
R22098 VSS.n2507 VSS.n2439 4.5005
R22099 VSS.n2508 VSS.n2439 4.5005
R22100 VSS.n2510 VSS.n2439 4.5005
R22101 VSS.n2513 VSS.n2439 4.5005
R22102 VSS.n2515 VSS.n2439 4.5005
R22103 VSS.n2516 VSS.n2439 4.5005
R22104 VSS.n2518 VSS.n2439 4.5005
R22105 VSS.n2521 VSS.n2439 4.5005
R22106 VSS.n2523 VSS.n2439 4.5005
R22107 VSS.n2524 VSS.n2439 4.5005
R22108 VSS.n2526 VSS.n2439 4.5005
R22109 VSS.n2529 VSS.n2439 4.5005
R22110 VSS.n2531 VSS.n2439 4.5005
R22111 VSS.n2532 VSS.n2439 4.5005
R22112 VSS.n2534 VSS.n2439 4.5005
R22113 VSS.n2537 VSS.n2439 4.5005
R22114 VSS.n2539 VSS.n2439 4.5005
R22115 VSS.n2540 VSS.n2439 4.5005
R22116 VSS.n2542 VSS.n2439 4.5005
R22117 VSS.n2545 VSS.n2439 4.5005
R22118 VSS.n2547 VSS.n2439 4.5005
R22119 VSS.n2548 VSS.n2439 4.5005
R22120 VSS.n2550 VSS.n2439 4.5005
R22121 VSS.n2553 VSS.n2439 4.5005
R22122 VSS.n2555 VSS.n2439 4.5005
R22123 VSS.n2556 VSS.n2439 4.5005
R22124 VSS.n2558 VSS.n2439 4.5005
R22125 VSS.n2561 VSS.n2439 4.5005
R22126 VSS.n2563 VSS.n2439 4.5005
R22127 VSS.n2564 VSS.n2439 4.5005
R22128 VSS.n2566 VSS.n2439 4.5005
R22129 VSS.n2569 VSS.n2439 4.5005
R22130 VSS.n2571 VSS.n2439 4.5005
R22131 VSS.n2572 VSS.n2439 4.5005
R22132 VSS.n2574 VSS.n2439 4.5005
R22133 VSS.n2577 VSS.n2439 4.5005
R22134 VSS.n2579 VSS.n2439 4.5005
R22135 VSS.n2580 VSS.n2439 4.5005
R22136 VSS.n2582 VSS.n2439 4.5005
R22137 VSS.n2585 VSS.n2439 4.5005
R22138 VSS.n2587 VSS.n2439 4.5005
R22139 VSS.n2588 VSS.n2439 4.5005
R22140 VSS.n2590 VSS.n2439 4.5005
R22141 VSS.n2593 VSS.n2439 4.5005
R22142 VSS.n2595 VSS.n2439 4.5005
R22143 VSS.n2596 VSS.n2439 4.5005
R22144 VSS.n2598 VSS.n2439 4.5005
R22145 VSS.n2601 VSS.n2439 4.5005
R22146 VSS.n2603 VSS.n2439 4.5005
R22147 VSS.n2604 VSS.n2439 4.5005
R22148 VSS.n2606 VSS.n2439 4.5005
R22149 VSS.n2609 VSS.n2439 4.5005
R22150 VSS.n2611 VSS.n2439 4.5005
R22151 VSS.n2612 VSS.n2439 4.5005
R22152 VSS.n2614 VSS.n2439 4.5005
R22153 VSS.n2617 VSS.n2439 4.5005
R22154 VSS.n2619 VSS.n2439 4.5005
R22155 VSS.n2620 VSS.n2439 4.5005
R22156 VSS.n2622 VSS.n2439 4.5005
R22157 VSS.n2625 VSS.n2439 4.5005
R22158 VSS.n2627 VSS.n2439 4.5005
R22159 VSS.n2628 VSS.n2439 4.5005
R22160 VSS.n2630 VSS.n2439 4.5005
R22161 VSS.n2633 VSS.n2439 4.5005
R22162 VSS.n2635 VSS.n2439 4.5005
R22163 VSS.n2636 VSS.n2439 4.5005
R22164 VSS.n2638 VSS.n2439 4.5005
R22165 VSS.n2640 VSS.n2439 4.5005
R22166 VSS.n2642 VSS.n2439 4.5005
R22167 VSS.n2643 VSS.n2439 4.5005
R22168 VSS.n2645 VSS.n2439 4.5005
R22169 VSS.n2648 VSS.n2439 4.5005
R22170 VSS.n2650 VSS.n2439 4.5005
R22171 VSS.n2651 VSS.n2439 4.5005
R22172 VSS.n2653 VSS.n2439 4.5005
R22173 VSS.n2656 VSS.n2439 4.5005
R22174 VSS.n2658 VSS.n2439 4.5005
R22175 VSS.n2659 VSS.n2439 4.5005
R22176 VSS.n2661 VSS.n2439 4.5005
R22177 VSS.n2664 VSS.n2439 4.5005
R22178 VSS.n2666 VSS.n2439 4.5005
R22179 VSS.n2667 VSS.n2439 4.5005
R22180 VSS.n2669 VSS.n2439 4.5005
R22181 VSS.n2672 VSS.n2439 4.5005
R22182 VSS.n2674 VSS.n2439 4.5005
R22183 VSS.n2675 VSS.n2439 4.5005
R22184 VSS.n2677 VSS.n2439 4.5005
R22185 VSS.n2680 VSS.n2439 4.5005
R22186 VSS.n2682 VSS.n2439 4.5005
R22187 VSS.n2683 VSS.n2439 4.5005
R22188 VSS.n2685 VSS.n2439 4.5005
R22189 VSS.n2688 VSS.n2439 4.5005
R22190 VSS.n2690 VSS.n2439 4.5005
R22191 VSS.n2691 VSS.n2439 4.5005
R22192 VSS.n2693 VSS.n2439 4.5005
R22193 VSS.n2696 VSS.n2439 4.5005
R22194 VSS.n2698 VSS.n2439 4.5005
R22195 VSS.n2699 VSS.n2439 4.5005
R22196 VSS.n2701 VSS.n2439 4.5005
R22197 VSS.n2704 VSS.n2439 4.5005
R22198 VSS.n2706 VSS.n2439 4.5005
R22199 VSS.n2707 VSS.n2439 4.5005
R22200 VSS.n2709 VSS.n2439 4.5005
R22201 VSS.n2712 VSS.n2439 4.5005
R22202 VSS.n2714 VSS.n2439 4.5005
R22203 VSS.n2715 VSS.n2439 4.5005
R22204 VSS.n2717 VSS.n2439 4.5005
R22205 VSS.n2720 VSS.n2439 4.5005
R22206 VSS.n2722 VSS.n2439 4.5005
R22207 VSS.n2723 VSS.n2439 4.5005
R22208 VSS.n2725 VSS.n2439 4.5005
R22209 VSS.n2793 VSS.n2439 4.5005
R22210 VSS.n2859 VSS.n2439 4.5005
R22211 VSS.n3051 VSS.n2392 4.5005
R22212 VSS.n2392 VSS.n2351 4.5005
R22213 VSS.n2483 VSS.n2392 4.5005
R22214 VSS.n2484 VSS.n2392 4.5005
R22215 VSS.n2486 VSS.n2392 4.5005
R22216 VSS.n2489 VSS.n2392 4.5005
R22217 VSS.n2491 VSS.n2392 4.5005
R22218 VSS.n2492 VSS.n2392 4.5005
R22219 VSS.n2494 VSS.n2392 4.5005
R22220 VSS.n2497 VSS.n2392 4.5005
R22221 VSS.n2499 VSS.n2392 4.5005
R22222 VSS.n2500 VSS.n2392 4.5005
R22223 VSS.n2502 VSS.n2392 4.5005
R22224 VSS.n2505 VSS.n2392 4.5005
R22225 VSS.n2507 VSS.n2392 4.5005
R22226 VSS.n2508 VSS.n2392 4.5005
R22227 VSS.n2510 VSS.n2392 4.5005
R22228 VSS.n2513 VSS.n2392 4.5005
R22229 VSS.n2515 VSS.n2392 4.5005
R22230 VSS.n2516 VSS.n2392 4.5005
R22231 VSS.n2518 VSS.n2392 4.5005
R22232 VSS.n2521 VSS.n2392 4.5005
R22233 VSS.n2523 VSS.n2392 4.5005
R22234 VSS.n2524 VSS.n2392 4.5005
R22235 VSS.n2526 VSS.n2392 4.5005
R22236 VSS.n2529 VSS.n2392 4.5005
R22237 VSS.n2531 VSS.n2392 4.5005
R22238 VSS.n2532 VSS.n2392 4.5005
R22239 VSS.n2534 VSS.n2392 4.5005
R22240 VSS.n2537 VSS.n2392 4.5005
R22241 VSS.n2539 VSS.n2392 4.5005
R22242 VSS.n2540 VSS.n2392 4.5005
R22243 VSS.n2542 VSS.n2392 4.5005
R22244 VSS.n2545 VSS.n2392 4.5005
R22245 VSS.n2547 VSS.n2392 4.5005
R22246 VSS.n2548 VSS.n2392 4.5005
R22247 VSS.n2550 VSS.n2392 4.5005
R22248 VSS.n2553 VSS.n2392 4.5005
R22249 VSS.n2555 VSS.n2392 4.5005
R22250 VSS.n2556 VSS.n2392 4.5005
R22251 VSS.n2558 VSS.n2392 4.5005
R22252 VSS.n2561 VSS.n2392 4.5005
R22253 VSS.n2563 VSS.n2392 4.5005
R22254 VSS.n2564 VSS.n2392 4.5005
R22255 VSS.n2566 VSS.n2392 4.5005
R22256 VSS.n2569 VSS.n2392 4.5005
R22257 VSS.n2571 VSS.n2392 4.5005
R22258 VSS.n2572 VSS.n2392 4.5005
R22259 VSS.n2574 VSS.n2392 4.5005
R22260 VSS.n2577 VSS.n2392 4.5005
R22261 VSS.n2579 VSS.n2392 4.5005
R22262 VSS.n2580 VSS.n2392 4.5005
R22263 VSS.n2582 VSS.n2392 4.5005
R22264 VSS.n2585 VSS.n2392 4.5005
R22265 VSS.n2587 VSS.n2392 4.5005
R22266 VSS.n2588 VSS.n2392 4.5005
R22267 VSS.n2590 VSS.n2392 4.5005
R22268 VSS.n2593 VSS.n2392 4.5005
R22269 VSS.n2595 VSS.n2392 4.5005
R22270 VSS.n2596 VSS.n2392 4.5005
R22271 VSS.n2598 VSS.n2392 4.5005
R22272 VSS.n2601 VSS.n2392 4.5005
R22273 VSS.n2603 VSS.n2392 4.5005
R22274 VSS.n2604 VSS.n2392 4.5005
R22275 VSS.n2606 VSS.n2392 4.5005
R22276 VSS.n2609 VSS.n2392 4.5005
R22277 VSS.n2611 VSS.n2392 4.5005
R22278 VSS.n2612 VSS.n2392 4.5005
R22279 VSS.n2614 VSS.n2392 4.5005
R22280 VSS.n2617 VSS.n2392 4.5005
R22281 VSS.n2619 VSS.n2392 4.5005
R22282 VSS.n2620 VSS.n2392 4.5005
R22283 VSS.n2622 VSS.n2392 4.5005
R22284 VSS.n2625 VSS.n2392 4.5005
R22285 VSS.n2627 VSS.n2392 4.5005
R22286 VSS.n2628 VSS.n2392 4.5005
R22287 VSS.n2630 VSS.n2392 4.5005
R22288 VSS.n2633 VSS.n2392 4.5005
R22289 VSS.n2635 VSS.n2392 4.5005
R22290 VSS.n2636 VSS.n2392 4.5005
R22291 VSS.n2638 VSS.n2392 4.5005
R22292 VSS.n2640 VSS.n2392 4.5005
R22293 VSS.n2642 VSS.n2392 4.5005
R22294 VSS.n2643 VSS.n2392 4.5005
R22295 VSS.n2645 VSS.n2392 4.5005
R22296 VSS.n2648 VSS.n2392 4.5005
R22297 VSS.n2650 VSS.n2392 4.5005
R22298 VSS.n2651 VSS.n2392 4.5005
R22299 VSS.n2653 VSS.n2392 4.5005
R22300 VSS.n2656 VSS.n2392 4.5005
R22301 VSS.n2658 VSS.n2392 4.5005
R22302 VSS.n2659 VSS.n2392 4.5005
R22303 VSS.n2661 VSS.n2392 4.5005
R22304 VSS.n2664 VSS.n2392 4.5005
R22305 VSS.n2666 VSS.n2392 4.5005
R22306 VSS.n2667 VSS.n2392 4.5005
R22307 VSS.n2669 VSS.n2392 4.5005
R22308 VSS.n2672 VSS.n2392 4.5005
R22309 VSS.n2674 VSS.n2392 4.5005
R22310 VSS.n2675 VSS.n2392 4.5005
R22311 VSS.n2677 VSS.n2392 4.5005
R22312 VSS.n2680 VSS.n2392 4.5005
R22313 VSS.n2682 VSS.n2392 4.5005
R22314 VSS.n2683 VSS.n2392 4.5005
R22315 VSS.n2685 VSS.n2392 4.5005
R22316 VSS.n2688 VSS.n2392 4.5005
R22317 VSS.n2690 VSS.n2392 4.5005
R22318 VSS.n2691 VSS.n2392 4.5005
R22319 VSS.n2693 VSS.n2392 4.5005
R22320 VSS.n2696 VSS.n2392 4.5005
R22321 VSS.n2698 VSS.n2392 4.5005
R22322 VSS.n2699 VSS.n2392 4.5005
R22323 VSS.n2701 VSS.n2392 4.5005
R22324 VSS.n2704 VSS.n2392 4.5005
R22325 VSS.n2706 VSS.n2392 4.5005
R22326 VSS.n2707 VSS.n2392 4.5005
R22327 VSS.n2709 VSS.n2392 4.5005
R22328 VSS.n2712 VSS.n2392 4.5005
R22329 VSS.n2714 VSS.n2392 4.5005
R22330 VSS.n2715 VSS.n2392 4.5005
R22331 VSS.n2717 VSS.n2392 4.5005
R22332 VSS.n2720 VSS.n2392 4.5005
R22333 VSS.n2722 VSS.n2392 4.5005
R22334 VSS.n2723 VSS.n2392 4.5005
R22335 VSS.n2725 VSS.n2392 4.5005
R22336 VSS.n2793 VSS.n2392 4.5005
R22337 VSS.n2859 VSS.n2392 4.5005
R22338 VSS.n3051 VSS.n2440 4.5005
R22339 VSS.n2440 VSS.n2351 4.5005
R22340 VSS.n2483 VSS.n2440 4.5005
R22341 VSS.n2484 VSS.n2440 4.5005
R22342 VSS.n2486 VSS.n2440 4.5005
R22343 VSS.n2489 VSS.n2440 4.5005
R22344 VSS.n2491 VSS.n2440 4.5005
R22345 VSS.n2492 VSS.n2440 4.5005
R22346 VSS.n2494 VSS.n2440 4.5005
R22347 VSS.n2497 VSS.n2440 4.5005
R22348 VSS.n2499 VSS.n2440 4.5005
R22349 VSS.n2500 VSS.n2440 4.5005
R22350 VSS.n2502 VSS.n2440 4.5005
R22351 VSS.n2505 VSS.n2440 4.5005
R22352 VSS.n2507 VSS.n2440 4.5005
R22353 VSS.n2508 VSS.n2440 4.5005
R22354 VSS.n2510 VSS.n2440 4.5005
R22355 VSS.n2513 VSS.n2440 4.5005
R22356 VSS.n2515 VSS.n2440 4.5005
R22357 VSS.n2516 VSS.n2440 4.5005
R22358 VSS.n2518 VSS.n2440 4.5005
R22359 VSS.n2521 VSS.n2440 4.5005
R22360 VSS.n2523 VSS.n2440 4.5005
R22361 VSS.n2524 VSS.n2440 4.5005
R22362 VSS.n2526 VSS.n2440 4.5005
R22363 VSS.n2529 VSS.n2440 4.5005
R22364 VSS.n2531 VSS.n2440 4.5005
R22365 VSS.n2532 VSS.n2440 4.5005
R22366 VSS.n2534 VSS.n2440 4.5005
R22367 VSS.n2537 VSS.n2440 4.5005
R22368 VSS.n2539 VSS.n2440 4.5005
R22369 VSS.n2540 VSS.n2440 4.5005
R22370 VSS.n2542 VSS.n2440 4.5005
R22371 VSS.n2545 VSS.n2440 4.5005
R22372 VSS.n2547 VSS.n2440 4.5005
R22373 VSS.n2548 VSS.n2440 4.5005
R22374 VSS.n2550 VSS.n2440 4.5005
R22375 VSS.n2553 VSS.n2440 4.5005
R22376 VSS.n2555 VSS.n2440 4.5005
R22377 VSS.n2556 VSS.n2440 4.5005
R22378 VSS.n2558 VSS.n2440 4.5005
R22379 VSS.n2561 VSS.n2440 4.5005
R22380 VSS.n2563 VSS.n2440 4.5005
R22381 VSS.n2564 VSS.n2440 4.5005
R22382 VSS.n2566 VSS.n2440 4.5005
R22383 VSS.n2569 VSS.n2440 4.5005
R22384 VSS.n2571 VSS.n2440 4.5005
R22385 VSS.n2572 VSS.n2440 4.5005
R22386 VSS.n2574 VSS.n2440 4.5005
R22387 VSS.n2577 VSS.n2440 4.5005
R22388 VSS.n2579 VSS.n2440 4.5005
R22389 VSS.n2580 VSS.n2440 4.5005
R22390 VSS.n2582 VSS.n2440 4.5005
R22391 VSS.n2585 VSS.n2440 4.5005
R22392 VSS.n2587 VSS.n2440 4.5005
R22393 VSS.n2588 VSS.n2440 4.5005
R22394 VSS.n2590 VSS.n2440 4.5005
R22395 VSS.n2593 VSS.n2440 4.5005
R22396 VSS.n2595 VSS.n2440 4.5005
R22397 VSS.n2596 VSS.n2440 4.5005
R22398 VSS.n2598 VSS.n2440 4.5005
R22399 VSS.n2601 VSS.n2440 4.5005
R22400 VSS.n2603 VSS.n2440 4.5005
R22401 VSS.n2604 VSS.n2440 4.5005
R22402 VSS.n2606 VSS.n2440 4.5005
R22403 VSS.n2609 VSS.n2440 4.5005
R22404 VSS.n2611 VSS.n2440 4.5005
R22405 VSS.n2612 VSS.n2440 4.5005
R22406 VSS.n2614 VSS.n2440 4.5005
R22407 VSS.n2617 VSS.n2440 4.5005
R22408 VSS.n2619 VSS.n2440 4.5005
R22409 VSS.n2620 VSS.n2440 4.5005
R22410 VSS.n2622 VSS.n2440 4.5005
R22411 VSS.n2625 VSS.n2440 4.5005
R22412 VSS.n2627 VSS.n2440 4.5005
R22413 VSS.n2628 VSS.n2440 4.5005
R22414 VSS.n2630 VSS.n2440 4.5005
R22415 VSS.n2633 VSS.n2440 4.5005
R22416 VSS.n2635 VSS.n2440 4.5005
R22417 VSS.n2636 VSS.n2440 4.5005
R22418 VSS.n2638 VSS.n2440 4.5005
R22419 VSS.n2640 VSS.n2440 4.5005
R22420 VSS.n2642 VSS.n2440 4.5005
R22421 VSS.n2643 VSS.n2440 4.5005
R22422 VSS.n2645 VSS.n2440 4.5005
R22423 VSS.n2648 VSS.n2440 4.5005
R22424 VSS.n2650 VSS.n2440 4.5005
R22425 VSS.n2651 VSS.n2440 4.5005
R22426 VSS.n2653 VSS.n2440 4.5005
R22427 VSS.n2656 VSS.n2440 4.5005
R22428 VSS.n2658 VSS.n2440 4.5005
R22429 VSS.n2659 VSS.n2440 4.5005
R22430 VSS.n2661 VSS.n2440 4.5005
R22431 VSS.n2664 VSS.n2440 4.5005
R22432 VSS.n2666 VSS.n2440 4.5005
R22433 VSS.n2667 VSS.n2440 4.5005
R22434 VSS.n2669 VSS.n2440 4.5005
R22435 VSS.n2672 VSS.n2440 4.5005
R22436 VSS.n2674 VSS.n2440 4.5005
R22437 VSS.n2675 VSS.n2440 4.5005
R22438 VSS.n2677 VSS.n2440 4.5005
R22439 VSS.n2680 VSS.n2440 4.5005
R22440 VSS.n2682 VSS.n2440 4.5005
R22441 VSS.n2683 VSS.n2440 4.5005
R22442 VSS.n2685 VSS.n2440 4.5005
R22443 VSS.n2688 VSS.n2440 4.5005
R22444 VSS.n2690 VSS.n2440 4.5005
R22445 VSS.n2691 VSS.n2440 4.5005
R22446 VSS.n2693 VSS.n2440 4.5005
R22447 VSS.n2696 VSS.n2440 4.5005
R22448 VSS.n2698 VSS.n2440 4.5005
R22449 VSS.n2699 VSS.n2440 4.5005
R22450 VSS.n2701 VSS.n2440 4.5005
R22451 VSS.n2704 VSS.n2440 4.5005
R22452 VSS.n2706 VSS.n2440 4.5005
R22453 VSS.n2707 VSS.n2440 4.5005
R22454 VSS.n2709 VSS.n2440 4.5005
R22455 VSS.n2712 VSS.n2440 4.5005
R22456 VSS.n2714 VSS.n2440 4.5005
R22457 VSS.n2715 VSS.n2440 4.5005
R22458 VSS.n2717 VSS.n2440 4.5005
R22459 VSS.n2720 VSS.n2440 4.5005
R22460 VSS.n2722 VSS.n2440 4.5005
R22461 VSS.n2723 VSS.n2440 4.5005
R22462 VSS.n2725 VSS.n2440 4.5005
R22463 VSS.n2793 VSS.n2440 4.5005
R22464 VSS.n2859 VSS.n2440 4.5005
R22465 VSS.n3051 VSS.n2391 4.5005
R22466 VSS.n2391 VSS.n2351 4.5005
R22467 VSS.n2483 VSS.n2391 4.5005
R22468 VSS.n2484 VSS.n2391 4.5005
R22469 VSS.n2486 VSS.n2391 4.5005
R22470 VSS.n2489 VSS.n2391 4.5005
R22471 VSS.n2491 VSS.n2391 4.5005
R22472 VSS.n2492 VSS.n2391 4.5005
R22473 VSS.n2494 VSS.n2391 4.5005
R22474 VSS.n2497 VSS.n2391 4.5005
R22475 VSS.n2499 VSS.n2391 4.5005
R22476 VSS.n2500 VSS.n2391 4.5005
R22477 VSS.n2502 VSS.n2391 4.5005
R22478 VSS.n2505 VSS.n2391 4.5005
R22479 VSS.n2507 VSS.n2391 4.5005
R22480 VSS.n2508 VSS.n2391 4.5005
R22481 VSS.n2510 VSS.n2391 4.5005
R22482 VSS.n2513 VSS.n2391 4.5005
R22483 VSS.n2515 VSS.n2391 4.5005
R22484 VSS.n2516 VSS.n2391 4.5005
R22485 VSS.n2518 VSS.n2391 4.5005
R22486 VSS.n2521 VSS.n2391 4.5005
R22487 VSS.n2523 VSS.n2391 4.5005
R22488 VSS.n2524 VSS.n2391 4.5005
R22489 VSS.n2526 VSS.n2391 4.5005
R22490 VSS.n2529 VSS.n2391 4.5005
R22491 VSS.n2531 VSS.n2391 4.5005
R22492 VSS.n2532 VSS.n2391 4.5005
R22493 VSS.n2534 VSS.n2391 4.5005
R22494 VSS.n2537 VSS.n2391 4.5005
R22495 VSS.n2539 VSS.n2391 4.5005
R22496 VSS.n2540 VSS.n2391 4.5005
R22497 VSS.n2542 VSS.n2391 4.5005
R22498 VSS.n2545 VSS.n2391 4.5005
R22499 VSS.n2547 VSS.n2391 4.5005
R22500 VSS.n2548 VSS.n2391 4.5005
R22501 VSS.n2550 VSS.n2391 4.5005
R22502 VSS.n2553 VSS.n2391 4.5005
R22503 VSS.n2555 VSS.n2391 4.5005
R22504 VSS.n2556 VSS.n2391 4.5005
R22505 VSS.n2558 VSS.n2391 4.5005
R22506 VSS.n2561 VSS.n2391 4.5005
R22507 VSS.n2563 VSS.n2391 4.5005
R22508 VSS.n2564 VSS.n2391 4.5005
R22509 VSS.n2566 VSS.n2391 4.5005
R22510 VSS.n2569 VSS.n2391 4.5005
R22511 VSS.n2571 VSS.n2391 4.5005
R22512 VSS.n2572 VSS.n2391 4.5005
R22513 VSS.n2574 VSS.n2391 4.5005
R22514 VSS.n2577 VSS.n2391 4.5005
R22515 VSS.n2579 VSS.n2391 4.5005
R22516 VSS.n2580 VSS.n2391 4.5005
R22517 VSS.n2582 VSS.n2391 4.5005
R22518 VSS.n2585 VSS.n2391 4.5005
R22519 VSS.n2587 VSS.n2391 4.5005
R22520 VSS.n2588 VSS.n2391 4.5005
R22521 VSS.n2590 VSS.n2391 4.5005
R22522 VSS.n2593 VSS.n2391 4.5005
R22523 VSS.n2595 VSS.n2391 4.5005
R22524 VSS.n2596 VSS.n2391 4.5005
R22525 VSS.n2598 VSS.n2391 4.5005
R22526 VSS.n2601 VSS.n2391 4.5005
R22527 VSS.n2603 VSS.n2391 4.5005
R22528 VSS.n2604 VSS.n2391 4.5005
R22529 VSS.n2606 VSS.n2391 4.5005
R22530 VSS.n2609 VSS.n2391 4.5005
R22531 VSS.n2611 VSS.n2391 4.5005
R22532 VSS.n2612 VSS.n2391 4.5005
R22533 VSS.n2614 VSS.n2391 4.5005
R22534 VSS.n2617 VSS.n2391 4.5005
R22535 VSS.n2619 VSS.n2391 4.5005
R22536 VSS.n2620 VSS.n2391 4.5005
R22537 VSS.n2622 VSS.n2391 4.5005
R22538 VSS.n2625 VSS.n2391 4.5005
R22539 VSS.n2627 VSS.n2391 4.5005
R22540 VSS.n2628 VSS.n2391 4.5005
R22541 VSS.n2630 VSS.n2391 4.5005
R22542 VSS.n2633 VSS.n2391 4.5005
R22543 VSS.n2635 VSS.n2391 4.5005
R22544 VSS.n2636 VSS.n2391 4.5005
R22545 VSS.n2638 VSS.n2391 4.5005
R22546 VSS.n2640 VSS.n2391 4.5005
R22547 VSS.n2642 VSS.n2391 4.5005
R22548 VSS.n2643 VSS.n2391 4.5005
R22549 VSS.n2645 VSS.n2391 4.5005
R22550 VSS.n2648 VSS.n2391 4.5005
R22551 VSS.n2650 VSS.n2391 4.5005
R22552 VSS.n2651 VSS.n2391 4.5005
R22553 VSS.n2653 VSS.n2391 4.5005
R22554 VSS.n2656 VSS.n2391 4.5005
R22555 VSS.n2658 VSS.n2391 4.5005
R22556 VSS.n2659 VSS.n2391 4.5005
R22557 VSS.n2661 VSS.n2391 4.5005
R22558 VSS.n2664 VSS.n2391 4.5005
R22559 VSS.n2666 VSS.n2391 4.5005
R22560 VSS.n2667 VSS.n2391 4.5005
R22561 VSS.n2669 VSS.n2391 4.5005
R22562 VSS.n2672 VSS.n2391 4.5005
R22563 VSS.n2674 VSS.n2391 4.5005
R22564 VSS.n2675 VSS.n2391 4.5005
R22565 VSS.n2677 VSS.n2391 4.5005
R22566 VSS.n2680 VSS.n2391 4.5005
R22567 VSS.n2682 VSS.n2391 4.5005
R22568 VSS.n2683 VSS.n2391 4.5005
R22569 VSS.n2685 VSS.n2391 4.5005
R22570 VSS.n2688 VSS.n2391 4.5005
R22571 VSS.n2690 VSS.n2391 4.5005
R22572 VSS.n2691 VSS.n2391 4.5005
R22573 VSS.n2693 VSS.n2391 4.5005
R22574 VSS.n2696 VSS.n2391 4.5005
R22575 VSS.n2698 VSS.n2391 4.5005
R22576 VSS.n2699 VSS.n2391 4.5005
R22577 VSS.n2701 VSS.n2391 4.5005
R22578 VSS.n2704 VSS.n2391 4.5005
R22579 VSS.n2706 VSS.n2391 4.5005
R22580 VSS.n2707 VSS.n2391 4.5005
R22581 VSS.n2709 VSS.n2391 4.5005
R22582 VSS.n2712 VSS.n2391 4.5005
R22583 VSS.n2714 VSS.n2391 4.5005
R22584 VSS.n2715 VSS.n2391 4.5005
R22585 VSS.n2717 VSS.n2391 4.5005
R22586 VSS.n2720 VSS.n2391 4.5005
R22587 VSS.n2722 VSS.n2391 4.5005
R22588 VSS.n2723 VSS.n2391 4.5005
R22589 VSS.n2725 VSS.n2391 4.5005
R22590 VSS.n2793 VSS.n2391 4.5005
R22591 VSS.n2859 VSS.n2391 4.5005
R22592 VSS.n3051 VSS.n2441 4.5005
R22593 VSS.n2441 VSS.n2351 4.5005
R22594 VSS.n2483 VSS.n2441 4.5005
R22595 VSS.n2484 VSS.n2441 4.5005
R22596 VSS.n2486 VSS.n2441 4.5005
R22597 VSS.n2489 VSS.n2441 4.5005
R22598 VSS.n2491 VSS.n2441 4.5005
R22599 VSS.n2492 VSS.n2441 4.5005
R22600 VSS.n2494 VSS.n2441 4.5005
R22601 VSS.n2497 VSS.n2441 4.5005
R22602 VSS.n2499 VSS.n2441 4.5005
R22603 VSS.n2500 VSS.n2441 4.5005
R22604 VSS.n2502 VSS.n2441 4.5005
R22605 VSS.n2505 VSS.n2441 4.5005
R22606 VSS.n2507 VSS.n2441 4.5005
R22607 VSS.n2508 VSS.n2441 4.5005
R22608 VSS.n2510 VSS.n2441 4.5005
R22609 VSS.n2513 VSS.n2441 4.5005
R22610 VSS.n2515 VSS.n2441 4.5005
R22611 VSS.n2516 VSS.n2441 4.5005
R22612 VSS.n2518 VSS.n2441 4.5005
R22613 VSS.n2521 VSS.n2441 4.5005
R22614 VSS.n2523 VSS.n2441 4.5005
R22615 VSS.n2524 VSS.n2441 4.5005
R22616 VSS.n2526 VSS.n2441 4.5005
R22617 VSS.n2529 VSS.n2441 4.5005
R22618 VSS.n2531 VSS.n2441 4.5005
R22619 VSS.n2532 VSS.n2441 4.5005
R22620 VSS.n2534 VSS.n2441 4.5005
R22621 VSS.n2537 VSS.n2441 4.5005
R22622 VSS.n2539 VSS.n2441 4.5005
R22623 VSS.n2540 VSS.n2441 4.5005
R22624 VSS.n2542 VSS.n2441 4.5005
R22625 VSS.n2545 VSS.n2441 4.5005
R22626 VSS.n2547 VSS.n2441 4.5005
R22627 VSS.n2548 VSS.n2441 4.5005
R22628 VSS.n2550 VSS.n2441 4.5005
R22629 VSS.n2553 VSS.n2441 4.5005
R22630 VSS.n2555 VSS.n2441 4.5005
R22631 VSS.n2556 VSS.n2441 4.5005
R22632 VSS.n2558 VSS.n2441 4.5005
R22633 VSS.n2561 VSS.n2441 4.5005
R22634 VSS.n2563 VSS.n2441 4.5005
R22635 VSS.n2564 VSS.n2441 4.5005
R22636 VSS.n2566 VSS.n2441 4.5005
R22637 VSS.n2569 VSS.n2441 4.5005
R22638 VSS.n2571 VSS.n2441 4.5005
R22639 VSS.n2572 VSS.n2441 4.5005
R22640 VSS.n2574 VSS.n2441 4.5005
R22641 VSS.n2577 VSS.n2441 4.5005
R22642 VSS.n2579 VSS.n2441 4.5005
R22643 VSS.n2580 VSS.n2441 4.5005
R22644 VSS.n2582 VSS.n2441 4.5005
R22645 VSS.n2585 VSS.n2441 4.5005
R22646 VSS.n2587 VSS.n2441 4.5005
R22647 VSS.n2588 VSS.n2441 4.5005
R22648 VSS.n2590 VSS.n2441 4.5005
R22649 VSS.n2593 VSS.n2441 4.5005
R22650 VSS.n2595 VSS.n2441 4.5005
R22651 VSS.n2596 VSS.n2441 4.5005
R22652 VSS.n2598 VSS.n2441 4.5005
R22653 VSS.n2601 VSS.n2441 4.5005
R22654 VSS.n2603 VSS.n2441 4.5005
R22655 VSS.n2604 VSS.n2441 4.5005
R22656 VSS.n2606 VSS.n2441 4.5005
R22657 VSS.n2609 VSS.n2441 4.5005
R22658 VSS.n2611 VSS.n2441 4.5005
R22659 VSS.n2612 VSS.n2441 4.5005
R22660 VSS.n2614 VSS.n2441 4.5005
R22661 VSS.n2617 VSS.n2441 4.5005
R22662 VSS.n2619 VSS.n2441 4.5005
R22663 VSS.n2620 VSS.n2441 4.5005
R22664 VSS.n2622 VSS.n2441 4.5005
R22665 VSS.n2625 VSS.n2441 4.5005
R22666 VSS.n2627 VSS.n2441 4.5005
R22667 VSS.n2628 VSS.n2441 4.5005
R22668 VSS.n2630 VSS.n2441 4.5005
R22669 VSS.n2633 VSS.n2441 4.5005
R22670 VSS.n2635 VSS.n2441 4.5005
R22671 VSS.n2636 VSS.n2441 4.5005
R22672 VSS.n2638 VSS.n2441 4.5005
R22673 VSS.n2640 VSS.n2441 4.5005
R22674 VSS.n2642 VSS.n2441 4.5005
R22675 VSS.n2643 VSS.n2441 4.5005
R22676 VSS.n2645 VSS.n2441 4.5005
R22677 VSS.n2648 VSS.n2441 4.5005
R22678 VSS.n2650 VSS.n2441 4.5005
R22679 VSS.n2651 VSS.n2441 4.5005
R22680 VSS.n2653 VSS.n2441 4.5005
R22681 VSS.n2656 VSS.n2441 4.5005
R22682 VSS.n2658 VSS.n2441 4.5005
R22683 VSS.n2659 VSS.n2441 4.5005
R22684 VSS.n2661 VSS.n2441 4.5005
R22685 VSS.n2664 VSS.n2441 4.5005
R22686 VSS.n2666 VSS.n2441 4.5005
R22687 VSS.n2667 VSS.n2441 4.5005
R22688 VSS.n2669 VSS.n2441 4.5005
R22689 VSS.n2672 VSS.n2441 4.5005
R22690 VSS.n2674 VSS.n2441 4.5005
R22691 VSS.n2675 VSS.n2441 4.5005
R22692 VSS.n2677 VSS.n2441 4.5005
R22693 VSS.n2680 VSS.n2441 4.5005
R22694 VSS.n2682 VSS.n2441 4.5005
R22695 VSS.n2683 VSS.n2441 4.5005
R22696 VSS.n2685 VSS.n2441 4.5005
R22697 VSS.n2688 VSS.n2441 4.5005
R22698 VSS.n2690 VSS.n2441 4.5005
R22699 VSS.n2691 VSS.n2441 4.5005
R22700 VSS.n2693 VSS.n2441 4.5005
R22701 VSS.n2696 VSS.n2441 4.5005
R22702 VSS.n2698 VSS.n2441 4.5005
R22703 VSS.n2699 VSS.n2441 4.5005
R22704 VSS.n2701 VSS.n2441 4.5005
R22705 VSS.n2704 VSS.n2441 4.5005
R22706 VSS.n2706 VSS.n2441 4.5005
R22707 VSS.n2707 VSS.n2441 4.5005
R22708 VSS.n2709 VSS.n2441 4.5005
R22709 VSS.n2712 VSS.n2441 4.5005
R22710 VSS.n2714 VSS.n2441 4.5005
R22711 VSS.n2715 VSS.n2441 4.5005
R22712 VSS.n2717 VSS.n2441 4.5005
R22713 VSS.n2720 VSS.n2441 4.5005
R22714 VSS.n2722 VSS.n2441 4.5005
R22715 VSS.n2723 VSS.n2441 4.5005
R22716 VSS.n2725 VSS.n2441 4.5005
R22717 VSS.n2793 VSS.n2441 4.5005
R22718 VSS.n2859 VSS.n2441 4.5005
R22719 VSS.n3051 VSS.n2390 4.5005
R22720 VSS.n2390 VSS.n2351 4.5005
R22721 VSS.n2483 VSS.n2390 4.5005
R22722 VSS.n2484 VSS.n2390 4.5005
R22723 VSS.n2486 VSS.n2390 4.5005
R22724 VSS.n2489 VSS.n2390 4.5005
R22725 VSS.n2491 VSS.n2390 4.5005
R22726 VSS.n2492 VSS.n2390 4.5005
R22727 VSS.n2494 VSS.n2390 4.5005
R22728 VSS.n2497 VSS.n2390 4.5005
R22729 VSS.n2499 VSS.n2390 4.5005
R22730 VSS.n2500 VSS.n2390 4.5005
R22731 VSS.n2502 VSS.n2390 4.5005
R22732 VSS.n2505 VSS.n2390 4.5005
R22733 VSS.n2507 VSS.n2390 4.5005
R22734 VSS.n2508 VSS.n2390 4.5005
R22735 VSS.n2510 VSS.n2390 4.5005
R22736 VSS.n2513 VSS.n2390 4.5005
R22737 VSS.n2515 VSS.n2390 4.5005
R22738 VSS.n2516 VSS.n2390 4.5005
R22739 VSS.n2518 VSS.n2390 4.5005
R22740 VSS.n2521 VSS.n2390 4.5005
R22741 VSS.n2523 VSS.n2390 4.5005
R22742 VSS.n2524 VSS.n2390 4.5005
R22743 VSS.n2526 VSS.n2390 4.5005
R22744 VSS.n2529 VSS.n2390 4.5005
R22745 VSS.n2531 VSS.n2390 4.5005
R22746 VSS.n2532 VSS.n2390 4.5005
R22747 VSS.n2534 VSS.n2390 4.5005
R22748 VSS.n2537 VSS.n2390 4.5005
R22749 VSS.n2539 VSS.n2390 4.5005
R22750 VSS.n2540 VSS.n2390 4.5005
R22751 VSS.n2542 VSS.n2390 4.5005
R22752 VSS.n2545 VSS.n2390 4.5005
R22753 VSS.n2547 VSS.n2390 4.5005
R22754 VSS.n2548 VSS.n2390 4.5005
R22755 VSS.n2550 VSS.n2390 4.5005
R22756 VSS.n2553 VSS.n2390 4.5005
R22757 VSS.n2555 VSS.n2390 4.5005
R22758 VSS.n2556 VSS.n2390 4.5005
R22759 VSS.n2558 VSS.n2390 4.5005
R22760 VSS.n2561 VSS.n2390 4.5005
R22761 VSS.n2563 VSS.n2390 4.5005
R22762 VSS.n2564 VSS.n2390 4.5005
R22763 VSS.n2566 VSS.n2390 4.5005
R22764 VSS.n2569 VSS.n2390 4.5005
R22765 VSS.n2571 VSS.n2390 4.5005
R22766 VSS.n2572 VSS.n2390 4.5005
R22767 VSS.n2574 VSS.n2390 4.5005
R22768 VSS.n2577 VSS.n2390 4.5005
R22769 VSS.n2579 VSS.n2390 4.5005
R22770 VSS.n2580 VSS.n2390 4.5005
R22771 VSS.n2582 VSS.n2390 4.5005
R22772 VSS.n2585 VSS.n2390 4.5005
R22773 VSS.n2587 VSS.n2390 4.5005
R22774 VSS.n2588 VSS.n2390 4.5005
R22775 VSS.n2590 VSS.n2390 4.5005
R22776 VSS.n2593 VSS.n2390 4.5005
R22777 VSS.n2595 VSS.n2390 4.5005
R22778 VSS.n2596 VSS.n2390 4.5005
R22779 VSS.n2598 VSS.n2390 4.5005
R22780 VSS.n2601 VSS.n2390 4.5005
R22781 VSS.n2603 VSS.n2390 4.5005
R22782 VSS.n2604 VSS.n2390 4.5005
R22783 VSS.n2606 VSS.n2390 4.5005
R22784 VSS.n2609 VSS.n2390 4.5005
R22785 VSS.n2611 VSS.n2390 4.5005
R22786 VSS.n2612 VSS.n2390 4.5005
R22787 VSS.n2614 VSS.n2390 4.5005
R22788 VSS.n2617 VSS.n2390 4.5005
R22789 VSS.n2619 VSS.n2390 4.5005
R22790 VSS.n2620 VSS.n2390 4.5005
R22791 VSS.n2622 VSS.n2390 4.5005
R22792 VSS.n2625 VSS.n2390 4.5005
R22793 VSS.n2627 VSS.n2390 4.5005
R22794 VSS.n2628 VSS.n2390 4.5005
R22795 VSS.n2630 VSS.n2390 4.5005
R22796 VSS.n2633 VSS.n2390 4.5005
R22797 VSS.n2635 VSS.n2390 4.5005
R22798 VSS.n2636 VSS.n2390 4.5005
R22799 VSS.n2638 VSS.n2390 4.5005
R22800 VSS.n2640 VSS.n2390 4.5005
R22801 VSS.n2642 VSS.n2390 4.5005
R22802 VSS.n2643 VSS.n2390 4.5005
R22803 VSS.n2645 VSS.n2390 4.5005
R22804 VSS.n2648 VSS.n2390 4.5005
R22805 VSS.n2650 VSS.n2390 4.5005
R22806 VSS.n2651 VSS.n2390 4.5005
R22807 VSS.n2653 VSS.n2390 4.5005
R22808 VSS.n2656 VSS.n2390 4.5005
R22809 VSS.n2658 VSS.n2390 4.5005
R22810 VSS.n2659 VSS.n2390 4.5005
R22811 VSS.n2661 VSS.n2390 4.5005
R22812 VSS.n2664 VSS.n2390 4.5005
R22813 VSS.n2666 VSS.n2390 4.5005
R22814 VSS.n2667 VSS.n2390 4.5005
R22815 VSS.n2669 VSS.n2390 4.5005
R22816 VSS.n2672 VSS.n2390 4.5005
R22817 VSS.n2674 VSS.n2390 4.5005
R22818 VSS.n2675 VSS.n2390 4.5005
R22819 VSS.n2677 VSS.n2390 4.5005
R22820 VSS.n2680 VSS.n2390 4.5005
R22821 VSS.n2682 VSS.n2390 4.5005
R22822 VSS.n2683 VSS.n2390 4.5005
R22823 VSS.n2685 VSS.n2390 4.5005
R22824 VSS.n2688 VSS.n2390 4.5005
R22825 VSS.n2690 VSS.n2390 4.5005
R22826 VSS.n2691 VSS.n2390 4.5005
R22827 VSS.n2693 VSS.n2390 4.5005
R22828 VSS.n2696 VSS.n2390 4.5005
R22829 VSS.n2698 VSS.n2390 4.5005
R22830 VSS.n2699 VSS.n2390 4.5005
R22831 VSS.n2701 VSS.n2390 4.5005
R22832 VSS.n2704 VSS.n2390 4.5005
R22833 VSS.n2706 VSS.n2390 4.5005
R22834 VSS.n2707 VSS.n2390 4.5005
R22835 VSS.n2709 VSS.n2390 4.5005
R22836 VSS.n2712 VSS.n2390 4.5005
R22837 VSS.n2714 VSS.n2390 4.5005
R22838 VSS.n2715 VSS.n2390 4.5005
R22839 VSS.n2717 VSS.n2390 4.5005
R22840 VSS.n2720 VSS.n2390 4.5005
R22841 VSS.n2722 VSS.n2390 4.5005
R22842 VSS.n2723 VSS.n2390 4.5005
R22843 VSS.n2725 VSS.n2390 4.5005
R22844 VSS.n2793 VSS.n2390 4.5005
R22845 VSS.n2859 VSS.n2390 4.5005
R22846 VSS.n3051 VSS.n2442 4.5005
R22847 VSS.n2442 VSS.n2351 4.5005
R22848 VSS.n2483 VSS.n2442 4.5005
R22849 VSS.n2484 VSS.n2442 4.5005
R22850 VSS.n2486 VSS.n2442 4.5005
R22851 VSS.n2489 VSS.n2442 4.5005
R22852 VSS.n2491 VSS.n2442 4.5005
R22853 VSS.n2492 VSS.n2442 4.5005
R22854 VSS.n2494 VSS.n2442 4.5005
R22855 VSS.n2497 VSS.n2442 4.5005
R22856 VSS.n2499 VSS.n2442 4.5005
R22857 VSS.n2500 VSS.n2442 4.5005
R22858 VSS.n2502 VSS.n2442 4.5005
R22859 VSS.n2505 VSS.n2442 4.5005
R22860 VSS.n2507 VSS.n2442 4.5005
R22861 VSS.n2508 VSS.n2442 4.5005
R22862 VSS.n2510 VSS.n2442 4.5005
R22863 VSS.n2513 VSS.n2442 4.5005
R22864 VSS.n2515 VSS.n2442 4.5005
R22865 VSS.n2516 VSS.n2442 4.5005
R22866 VSS.n2518 VSS.n2442 4.5005
R22867 VSS.n2521 VSS.n2442 4.5005
R22868 VSS.n2523 VSS.n2442 4.5005
R22869 VSS.n2524 VSS.n2442 4.5005
R22870 VSS.n2526 VSS.n2442 4.5005
R22871 VSS.n2529 VSS.n2442 4.5005
R22872 VSS.n2531 VSS.n2442 4.5005
R22873 VSS.n2532 VSS.n2442 4.5005
R22874 VSS.n2534 VSS.n2442 4.5005
R22875 VSS.n2537 VSS.n2442 4.5005
R22876 VSS.n2539 VSS.n2442 4.5005
R22877 VSS.n2540 VSS.n2442 4.5005
R22878 VSS.n2542 VSS.n2442 4.5005
R22879 VSS.n2545 VSS.n2442 4.5005
R22880 VSS.n2547 VSS.n2442 4.5005
R22881 VSS.n2548 VSS.n2442 4.5005
R22882 VSS.n2550 VSS.n2442 4.5005
R22883 VSS.n2553 VSS.n2442 4.5005
R22884 VSS.n2555 VSS.n2442 4.5005
R22885 VSS.n2556 VSS.n2442 4.5005
R22886 VSS.n2558 VSS.n2442 4.5005
R22887 VSS.n2561 VSS.n2442 4.5005
R22888 VSS.n2563 VSS.n2442 4.5005
R22889 VSS.n2564 VSS.n2442 4.5005
R22890 VSS.n2566 VSS.n2442 4.5005
R22891 VSS.n2569 VSS.n2442 4.5005
R22892 VSS.n2571 VSS.n2442 4.5005
R22893 VSS.n2572 VSS.n2442 4.5005
R22894 VSS.n2574 VSS.n2442 4.5005
R22895 VSS.n2577 VSS.n2442 4.5005
R22896 VSS.n2579 VSS.n2442 4.5005
R22897 VSS.n2580 VSS.n2442 4.5005
R22898 VSS.n2582 VSS.n2442 4.5005
R22899 VSS.n2585 VSS.n2442 4.5005
R22900 VSS.n2587 VSS.n2442 4.5005
R22901 VSS.n2588 VSS.n2442 4.5005
R22902 VSS.n2590 VSS.n2442 4.5005
R22903 VSS.n2593 VSS.n2442 4.5005
R22904 VSS.n2595 VSS.n2442 4.5005
R22905 VSS.n2596 VSS.n2442 4.5005
R22906 VSS.n2598 VSS.n2442 4.5005
R22907 VSS.n2601 VSS.n2442 4.5005
R22908 VSS.n2603 VSS.n2442 4.5005
R22909 VSS.n2604 VSS.n2442 4.5005
R22910 VSS.n2606 VSS.n2442 4.5005
R22911 VSS.n2609 VSS.n2442 4.5005
R22912 VSS.n2611 VSS.n2442 4.5005
R22913 VSS.n2612 VSS.n2442 4.5005
R22914 VSS.n2614 VSS.n2442 4.5005
R22915 VSS.n2617 VSS.n2442 4.5005
R22916 VSS.n2619 VSS.n2442 4.5005
R22917 VSS.n2620 VSS.n2442 4.5005
R22918 VSS.n2622 VSS.n2442 4.5005
R22919 VSS.n2625 VSS.n2442 4.5005
R22920 VSS.n2627 VSS.n2442 4.5005
R22921 VSS.n2628 VSS.n2442 4.5005
R22922 VSS.n2630 VSS.n2442 4.5005
R22923 VSS.n2633 VSS.n2442 4.5005
R22924 VSS.n2635 VSS.n2442 4.5005
R22925 VSS.n2636 VSS.n2442 4.5005
R22926 VSS.n2638 VSS.n2442 4.5005
R22927 VSS.n2640 VSS.n2442 4.5005
R22928 VSS.n2642 VSS.n2442 4.5005
R22929 VSS.n2643 VSS.n2442 4.5005
R22930 VSS.n2645 VSS.n2442 4.5005
R22931 VSS.n2648 VSS.n2442 4.5005
R22932 VSS.n2650 VSS.n2442 4.5005
R22933 VSS.n2651 VSS.n2442 4.5005
R22934 VSS.n2653 VSS.n2442 4.5005
R22935 VSS.n2656 VSS.n2442 4.5005
R22936 VSS.n2658 VSS.n2442 4.5005
R22937 VSS.n2659 VSS.n2442 4.5005
R22938 VSS.n2661 VSS.n2442 4.5005
R22939 VSS.n2664 VSS.n2442 4.5005
R22940 VSS.n2666 VSS.n2442 4.5005
R22941 VSS.n2667 VSS.n2442 4.5005
R22942 VSS.n2669 VSS.n2442 4.5005
R22943 VSS.n2672 VSS.n2442 4.5005
R22944 VSS.n2674 VSS.n2442 4.5005
R22945 VSS.n2675 VSS.n2442 4.5005
R22946 VSS.n2677 VSS.n2442 4.5005
R22947 VSS.n2680 VSS.n2442 4.5005
R22948 VSS.n2682 VSS.n2442 4.5005
R22949 VSS.n2683 VSS.n2442 4.5005
R22950 VSS.n2685 VSS.n2442 4.5005
R22951 VSS.n2688 VSS.n2442 4.5005
R22952 VSS.n2690 VSS.n2442 4.5005
R22953 VSS.n2691 VSS.n2442 4.5005
R22954 VSS.n2693 VSS.n2442 4.5005
R22955 VSS.n2696 VSS.n2442 4.5005
R22956 VSS.n2698 VSS.n2442 4.5005
R22957 VSS.n2699 VSS.n2442 4.5005
R22958 VSS.n2701 VSS.n2442 4.5005
R22959 VSS.n2704 VSS.n2442 4.5005
R22960 VSS.n2706 VSS.n2442 4.5005
R22961 VSS.n2707 VSS.n2442 4.5005
R22962 VSS.n2709 VSS.n2442 4.5005
R22963 VSS.n2712 VSS.n2442 4.5005
R22964 VSS.n2714 VSS.n2442 4.5005
R22965 VSS.n2715 VSS.n2442 4.5005
R22966 VSS.n2717 VSS.n2442 4.5005
R22967 VSS.n2720 VSS.n2442 4.5005
R22968 VSS.n2722 VSS.n2442 4.5005
R22969 VSS.n2723 VSS.n2442 4.5005
R22970 VSS.n2725 VSS.n2442 4.5005
R22971 VSS.n2793 VSS.n2442 4.5005
R22972 VSS.n2859 VSS.n2442 4.5005
R22973 VSS.n3051 VSS.n2389 4.5005
R22974 VSS.n2389 VSS.n2351 4.5005
R22975 VSS.n2483 VSS.n2389 4.5005
R22976 VSS.n2484 VSS.n2389 4.5005
R22977 VSS.n2486 VSS.n2389 4.5005
R22978 VSS.n2489 VSS.n2389 4.5005
R22979 VSS.n2491 VSS.n2389 4.5005
R22980 VSS.n2492 VSS.n2389 4.5005
R22981 VSS.n2494 VSS.n2389 4.5005
R22982 VSS.n2497 VSS.n2389 4.5005
R22983 VSS.n2499 VSS.n2389 4.5005
R22984 VSS.n2500 VSS.n2389 4.5005
R22985 VSS.n2502 VSS.n2389 4.5005
R22986 VSS.n2505 VSS.n2389 4.5005
R22987 VSS.n2507 VSS.n2389 4.5005
R22988 VSS.n2508 VSS.n2389 4.5005
R22989 VSS.n2510 VSS.n2389 4.5005
R22990 VSS.n2513 VSS.n2389 4.5005
R22991 VSS.n2515 VSS.n2389 4.5005
R22992 VSS.n2516 VSS.n2389 4.5005
R22993 VSS.n2518 VSS.n2389 4.5005
R22994 VSS.n2521 VSS.n2389 4.5005
R22995 VSS.n2523 VSS.n2389 4.5005
R22996 VSS.n2524 VSS.n2389 4.5005
R22997 VSS.n2526 VSS.n2389 4.5005
R22998 VSS.n2529 VSS.n2389 4.5005
R22999 VSS.n2531 VSS.n2389 4.5005
R23000 VSS.n2532 VSS.n2389 4.5005
R23001 VSS.n2534 VSS.n2389 4.5005
R23002 VSS.n2537 VSS.n2389 4.5005
R23003 VSS.n2539 VSS.n2389 4.5005
R23004 VSS.n2540 VSS.n2389 4.5005
R23005 VSS.n2542 VSS.n2389 4.5005
R23006 VSS.n2545 VSS.n2389 4.5005
R23007 VSS.n2547 VSS.n2389 4.5005
R23008 VSS.n2548 VSS.n2389 4.5005
R23009 VSS.n2550 VSS.n2389 4.5005
R23010 VSS.n2553 VSS.n2389 4.5005
R23011 VSS.n2555 VSS.n2389 4.5005
R23012 VSS.n2556 VSS.n2389 4.5005
R23013 VSS.n2558 VSS.n2389 4.5005
R23014 VSS.n2561 VSS.n2389 4.5005
R23015 VSS.n2563 VSS.n2389 4.5005
R23016 VSS.n2564 VSS.n2389 4.5005
R23017 VSS.n2566 VSS.n2389 4.5005
R23018 VSS.n2569 VSS.n2389 4.5005
R23019 VSS.n2571 VSS.n2389 4.5005
R23020 VSS.n2572 VSS.n2389 4.5005
R23021 VSS.n2574 VSS.n2389 4.5005
R23022 VSS.n2577 VSS.n2389 4.5005
R23023 VSS.n2579 VSS.n2389 4.5005
R23024 VSS.n2580 VSS.n2389 4.5005
R23025 VSS.n2582 VSS.n2389 4.5005
R23026 VSS.n2585 VSS.n2389 4.5005
R23027 VSS.n2587 VSS.n2389 4.5005
R23028 VSS.n2588 VSS.n2389 4.5005
R23029 VSS.n2590 VSS.n2389 4.5005
R23030 VSS.n2593 VSS.n2389 4.5005
R23031 VSS.n2595 VSS.n2389 4.5005
R23032 VSS.n2596 VSS.n2389 4.5005
R23033 VSS.n2598 VSS.n2389 4.5005
R23034 VSS.n2601 VSS.n2389 4.5005
R23035 VSS.n2603 VSS.n2389 4.5005
R23036 VSS.n2604 VSS.n2389 4.5005
R23037 VSS.n2606 VSS.n2389 4.5005
R23038 VSS.n2609 VSS.n2389 4.5005
R23039 VSS.n2611 VSS.n2389 4.5005
R23040 VSS.n2612 VSS.n2389 4.5005
R23041 VSS.n2614 VSS.n2389 4.5005
R23042 VSS.n2617 VSS.n2389 4.5005
R23043 VSS.n2619 VSS.n2389 4.5005
R23044 VSS.n2620 VSS.n2389 4.5005
R23045 VSS.n2622 VSS.n2389 4.5005
R23046 VSS.n2625 VSS.n2389 4.5005
R23047 VSS.n2627 VSS.n2389 4.5005
R23048 VSS.n2628 VSS.n2389 4.5005
R23049 VSS.n2630 VSS.n2389 4.5005
R23050 VSS.n2633 VSS.n2389 4.5005
R23051 VSS.n2635 VSS.n2389 4.5005
R23052 VSS.n2636 VSS.n2389 4.5005
R23053 VSS.n2638 VSS.n2389 4.5005
R23054 VSS.n2640 VSS.n2389 4.5005
R23055 VSS.n2642 VSS.n2389 4.5005
R23056 VSS.n2643 VSS.n2389 4.5005
R23057 VSS.n2645 VSS.n2389 4.5005
R23058 VSS.n2648 VSS.n2389 4.5005
R23059 VSS.n2650 VSS.n2389 4.5005
R23060 VSS.n2651 VSS.n2389 4.5005
R23061 VSS.n2653 VSS.n2389 4.5005
R23062 VSS.n2656 VSS.n2389 4.5005
R23063 VSS.n2658 VSS.n2389 4.5005
R23064 VSS.n2659 VSS.n2389 4.5005
R23065 VSS.n2661 VSS.n2389 4.5005
R23066 VSS.n2664 VSS.n2389 4.5005
R23067 VSS.n2666 VSS.n2389 4.5005
R23068 VSS.n2667 VSS.n2389 4.5005
R23069 VSS.n2669 VSS.n2389 4.5005
R23070 VSS.n2672 VSS.n2389 4.5005
R23071 VSS.n2674 VSS.n2389 4.5005
R23072 VSS.n2675 VSS.n2389 4.5005
R23073 VSS.n2677 VSS.n2389 4.5005
R23074 VSS.n2680 VSS.n2389 4.5005
R23075 VSS.n2682 VSS.n2389 4.5005
R23076 VSS.n2683 VSS.n2389 4.5005
R23077 VSS.n2685 VSS.n2389 4.5005
R23078 VSS.n2688 VSS.n2389 4.5005
R23079 VSS.n2690 VSS.n2389 4.5005
R23080 VSS.n2691 VSS.n2389 4.5005
R23081 VSS.n2693 VSS.n2389 4.5005
R23082 VSS.n2696 VSS.n2389 4.5005
R23083 VSS.n2698 VSS.n2389 4.5005
R23084 VSS.n2699 VSS.n2389 4.5005
R23085 VSS.n2701 VSS.n2389 4.5005
R23086 VSS.n2704 VSS.n2389 4.5005
R23087 VSS.n2706 VSS.n2389 4.5005
R23088 VSS.n2707 VSS.n2389 4.5005
R23089 VSS.n2709 VSS.n2389 4.5005
R23090 VSS.n2712 VSS.n2389 4.5005
R23091 VSS.n2714 VSS.n2389 4.5005
R23092 VSS.n2715 VSS.n2389 4.5005
R23093 VSS.n2717 VSS.n2389 4.5005
R23094 VSS.n2720 VSS.n2389 4.5005
R23095 VSS.n2722 VSS.n2389 4.5005
R23096 VSS.n2723 VSS.n2389 4.5005
R23097 VSS.n2725 VSS.n2389 4.5005
R23098 VSS.n2793 VSS.n2389 4.5005
R23099 VSS.n2859 VSS.n2389 4.5005
R23100 VSS.n3051 VSS.n2443 4.5005
R23101 VSS.n2443 VSS.n2351 4.5005
R23102 VSS.n2483 VSS.n2443 4.5005
R23103 VSS.n2484 VSS.n2443 4.5005
R23104 VSS.n2486 VSS.n2443 4.5005
R23105 VSS.n2489 VSS.n2443 4.5005
R23106 VSS.n2491 VSS.n2443 4.5005
R23107 VSS.n2492 VSS.n2443 4.5005
R23108 VSS.n2494 VSS.n2443 4.5005
R23109 VSS.n2497 VSS.n2443 4.5005
R23110 VSS.n2499 VSS.n2443 4.5005
R23111 VSS.n2500 VSS.n2443 4.5005
R23112 VSS.n2502 VSS.n2443 4.5005
R23113 VSS.n2505 VSS.n2443 4.5005
R23114 VSS.n2507 VSS.n2443 4.5005
R23115 VSS.n2508 VSS.n2443 4.5005
R23116 VSS.n2510 VSS.n2443 4.5005
R23117 VSS.n2513 VSS.n2443 4.5005
R23118 VSS.n2515 VSS.n2443 4.5005
R23119 VSS.n2516 VSS.n2443 4.5005
R23120 VSS.n2518 VSS.n2443 4.5005
R23121 VSS.n2521 VSS.n2443 4.5005
R23122 VSS.n2523 VSS.n2443 4.5005
R23123 VSS.n2524 VSS.n2443 4.5005
R23124 VSS.n2526 VSS.n2443 4.5005
R23125 VSS.n2529 VSS.n2443 4.5005
R23126 VSS.n2531 VSS.n2443 4.5005
R23127 VSS.n2532 VSS.n2443 4.5005
R23128 VSS.n2534 VSS.n2443 4.5005
R23129 VSS.n2537 VSS.n2443 4.5005
R23130 VSS.n2539 VSS.n2443 4.5005
R23131 VSS.n2540 VSS.n2443 4.5005
R23132 VSS.n2542 VSS.n2443 4.5005
R23133 VSS.n2545 VSS.n2443 4.5005
R23134 VSS.n2547 VSS.n2443 4.5005
R23135 VSS.n2548 VSS.n2443 4.5005
R23136 VSS.n2550 VSS.n2443 4.5005
R23137 VSS.n2553 VSS.n2443 4.5005
R23138 VSS.n2555 VSS.n2443 4.5005
R23139 VSS.n2556 VSS.n2443 4.5005
R23140 VSS.n2558 VSS.n2443 4.5005
R23141 VSS.n2561 VSS.n2443 4.5005
R23142 VSS.n2563 VSS.n2443 4.5005
R23143 VSS.n2564 VSS.n2443 4.5005
R23144 VSS.n2566 VSS.n2443 4.5005
R23145 VSS.n2569 VSS.n2443 4.5005
R23146 VSS.n2571 VSS.n2443 4.5005
R23147 VSS.n2572 VSS.n2443 4.5005
R23148 VSS.n2574 VSS.n2443 4.5005
R23149 VSS.n2577 VSS.n2443 4.5005
R23150 VSS.n2579 VSS.n2443 4.5005
R23151 VSS.n2580 VSS.n2443 4.5005
R23152 VSS.n2582 VSS.n2443 4.5005
R23153 VSS.n2585 VSS.n2443 4.5005
R23154 VSS.n2587 VSS.n2443 4.5005
R23155 VSS.n2588 VSS.n2443 4.5005
R23156 VSS.n2590 VSS.n2443 4.5005
R23157 VSS.n2593 VSS.n2443 4.5005
R23158 VSS.n2595 VSS.n2443 4.5005
R23159 VSS.n2596 VSS.n2443 4.5005
R23160 VSS.n2598 VSS.n2443 4.5005
R23161 VSS.n2601 VSS.n2443 4.5005
R23162 VSS.n2603 VSS.n2443 4.5005
R23163 VSS.n2604 VSS.n2443 4.5005
R23164 VSS.n2606 VSS.n2443 4.5005
R23165 VSS.n2609 VSS.n2443 4.5005
R23166 VSS.n2611 VSS.n2443 4.5005
R23167 VSS.n2612 VSS.n2443 4.5005
R23168 VSS.n2614 VSS.n2443 4.5005
R23169 VSS.n2617 VSS.n2443 4.5005
R23170 VSS.n2619 VSS.n2443 4.5005
R23171 VSS.n2620 VSS.n2443 4.5005
R23172 VSS.n2622 VSS.n2443 4.5005
R23173 VSS.n2625 VSS.n2443 4.5005
R23174 VSS.n2627 VSS.n2443 4.5005
R23175 VSS.n2628 VSS.n2443 4.5005
R23176 VSS.n2630 VSS.n2443 4.5005
R23177 VSS.n2633 VSS.n2443 4.5005
R23178 VSS.n2635 VSS.n2443 4.5005
R23179 VSS.n2636 VSS.n2443 4.5005
R23180 VSS.n2638 VSS.n2443 4.5005
R23181 VSS.n2640 VSS.n2443 4.5005
R23182 VSS.n2642 VSS.n2443 4.5005
R23183 VSS.n2643 VSS.n2443 4.5005
R23184 VSS.n2645 VSS.n2443 4.5005
R23185 VSS.n2648 VSS.n2443 4.5005
R23186 VSS.n2650 VSS.n2443 4.5005
R23187 VSS.n2651 VSS.n2443 4.5005
R23188 VSS.n2653 VSS.n2443 4.5005
R23189 VSS.n2656 VSS.n2443 4.5005
R23190 VSS.n2658 VSS.n2443 4.5005
R23191 VSS.n2659 VSS.n2443 4.5005
R23192 VSS.n2661 VSS.n2443 4.5005
R23193 VSS.n2664 VSS.n2443 4.5005
R23194 VSS.n2666 VSS.n2443 4.5005
R23195 VSS.n2667 VSS.n2443 4.5005
R23196 VSS.n2669 VSS.n2443 4.5005
R23197 VSS.n2672 VSS.n2443 4.5005
R23198 VSS.n2674 VSS.n2443 4.5005
R23199 VSS.n2675 VSS.n2443 4.5005
R23200 VSS.n2677 VSS.n2443 4.5005
R23201 VSS.n2680 VSS.n2443 4.5005
R23202 VSS.n2682 VSS.n2443 4.5005
R23203 VSS.n2683 VSS.n2443 4.5005
R23204 VSS.n2685 VSS.n2443 4.5005
R23205 VSS.n2688 VSS.n2443 4.5005
R23206 VSS.n2690 VSS.n2443 4.5005
R23207 VSS.n2691 VSS.n2443 4.5005
R23208 VSS.n2693 VSS.n2443 4.5005
R23209 VSS.n2696 VSS.n2443 4.5005
R23210 VSS.n2698 VSS.n2443 4.5005
R23211 VSS.n2699 VSS.n2443 4.5005
R23212 VSS.n2701 VSS.n2443 4.5005
R23213 VSS.n2704 VSS.n2443 4.5005
R23214 VSS.n2706 VSS.n2443 4.5005
R23215 VSS.n2707 VSS.n2443 4.5005
R23216 VSS.n2709 VSS.n2443 4.5005
R23217 VSS.n2712 VSS.n2443 4.5005
R23218 VSS.n2714 VSS.n2443 4.5005
R23219 VSS.n2715 VSS.n2443 4.5005
R23220 VSS.n2717 VSS.n2443 4.5005
R23221 VSS.n2720 VSS.n2443 4.5005
R23222 VSS.n2722 VSS.n2443 4.5005
R23223 VSS.n2723 VSS.n2443 4.5005
R23224 VSS.n2725 VSS.n2443 4.5005
R23225 VSS.n2793 VSS.n2443 4.5005
R23226 VSS.n2859 VSS.n2443 4.5005
R23227 VSS.n3051 VSS.n2388 4.5005
R23228 VSS.n2388 VSS.n2351 4.5005
R23229 VSS.n2483 VSS.n2388 4.5005
R23230 VSS.n2484 VSS.n2388 4.5005
R23231 VSS.n2486 VSS.n2388 4.5005
R23232 VSS.n2489 VSS.n2388 4.5005
R23233 VSS.n2491 VSS.n2388 4.5005
R23234 VSS.n2492 VSS.n2388 4.5005
R23235 VSS.n2494 VSS.n2388 4.5005
R23236 VSS.n2497 VSS.n2388 4.5005
R23237 VSS.n2499 VSS.n2388 4.5005
R23238 VSS.n2500 VSS.n2388 4.5005
R23239 VSS.n2502 VSS.n2388 4.5005
R23240 VSS.n2505 VSS.n2388 4.5005
R23241 VSS.n2507 VSS.n2388 4.5005
R23242 VSS.n2508 VSS.n2388 4.5005
R23243 VSS.n2510 VSS.n2388 4.5005
R23244 VSS.n2513 VSS.n2388 4.5005
R23245 VSS.n2515 VSS.n2388 4.5005
R23246 VSS.n2516 VSS.n2388 4.5005
R23247 VSS.n2518 VSS.n2388 4.5005
R23248 VSS.n2521 VSS.n2388 4.5005
R23249 VSS.n2523 VSS.n2388 4.5005
R23250 VSS.n2524 VSS.n2388 4.5005
R23251 VSS.n2526 VSS.n2388 4.5005
R23252 VSS.n2529 VSS.n2388 4.5005
R23253 VSS.n2531 VSS.n2388 4.5005
R23254 VSS.n2532 VSS.n2388 4.5005
R23255 VSS.n2534 VSS.n2388 4.5005
R23256 VSS.n2537 VSS.n2388 4.5005
R23257 VSS.n2539 VSS.n2388 4.5005
R23258 VSS.n2540 VSS.n2388 4.5005
R23259 VSS.n2542 VSS.n2388 4.5005
R23260 VSS.n2545 VSS.n2388 4.5005
R23261 VSS.n2547 VSS.n2388 4.5005
R23262 VSS.n2548 VSS.n2388 4.5005
R23263 VSS.n2550 VSS.n2388 4.5005
R23264 VSS.n2553 VSS.n2388 4.5005
R23265 VSS.n2555 VSS.n2388 4.5005
R23266 VSS.n2556 VSS.n2388 4.5005
R23267 VSS.n2558 VSS.n2388 4.5005
R23268 VSS.n2561 VSS.n2388 4.5005
R23269 VSS.n2563 VSS.n2388 4.5005
R23270 VSS.n2564 VSS.n2388 4.5005
R23271 VSS.n2566 VSS.n2388 4.5005
R23272 VSS.n2569 VSS.n2388 4.5005
R23273 VSS.n2571 VSS.n2388 4.5005
R23274 VSS.n2572 VSS.n2388 4.5005
R23275 VSS.n2574 VSS.n2388 4.5005
R23276 VSS.n2577 VSS.n2388 4.5005
R23277 VSS.n2579 VSS.n2388 4.5005
R23278 VSS.n2580 VSS.n2388 4.5005
R23279 VSS.n2582 VSS.n2388 4.5005
R23280 VSS.n2585 VSS.n2388 4.5005
R23281 VSS.n2587 VSS.n2388 4.5005
R23282 VSS.n2588 VSS.n2388 4.5005
R23283 VSS.n2590 VSS.n2388 4.5005
R23284 VSS.n2593 VSS.n2388 4.5005
R23285 VSS.n2595 VSS.n2388 4.5005
R23286 VSS.n2596 VSS.n2388 4.5005
R23287 VSS.n2598 VSS.n2388 4.5005
R23288 VSS.n2601 VSS.n2388 4.5005
R23289 VSS.n2603 VSS.n2388 4.5005
R23290 VSS.n2604 VSS.n2388 4.5005
R23291 VSS.n2606 VSS.n2388 4.5005
R23292 VSS.n2609 VSS.n2388 4.5005
R23293 VSS.n2611 VSS.n2388 4.5005
R23294 VSS.n2612 VSS.n2388 4.5005
R23295 VSS.n2614 VSS.n2388 4.5005
R23296 VSS.n2617 VSS.n2388 4.5005
R23297 VSS.n2619 VSS.n2388 4.5005
R23298 VSS.n2620 VSS.n2388 4.5005
R23299 VSS.n2622 VSS.n2388 4.5005
R23300 VSS.n2625 VSS.n2388 4.5005
R23301 VSS.n2627 VSS.n2388 4.5005
R23302 VSS.n2628 VSS.n2388 4.5005
R23303 VSS.n2630 VSS.n2388 4.5005
R23304 VSS.n2633 VSS.n2388 4.5005
R23305 VSS.n2635 VSS.n2388 4.5005
R23306 VSS.n2636 VSS.n2388 4.5005
R23307 VSS.n2638 VSS.n2388 4.5005
R23308 VSS.n2640 VSS.n2388 4.5005
R23309 VSS.n2642 VSS.n2388 4.5005
R23310 VSS.n2643 VSS.n2388 4.5005
R23311 VSS.n2645 VSS.n2388 4.5005
R23312 VSS.n2648 VSS.n2388 4.5005
R23313 VSS.n2650 VSS.n2388 4.5005
R23314 VSS.n2651 VSS.n2388 4.5005
R23315 VSS.n2653 VSS.n2388 4.5005
R23316 VSS.n2656 VSS.n2388 4.5005
R23317 VSS.n2658 VSS.n2388 4.5005
R23318 VSS.n2659 VSS.n2388 4.5005
R23319 VSS.n2661 VSS.n2388 4.5005
R23320 VSS.n2664 VSS.n2388 4.5005
R23321 VSS.n2666 VSS.n2388 4.5005
R23322 VSS.n2667 VSS.n2388 4.5005
R23323 VSS.n2669 VSS.n2388 4.5005
R23324 VSS.n2672 VSS.n2388 4.5005
R23325 VSS.n2674 VSS.n2388 4.5005
R23326 VSS.n2675 VSS.n2388 4.5005
R23327 VSS.n2677 VSS.n2388 4.5005
R23328 VSS.n2680 VSS.n2388 4.5005
R23329 VSS.n2682 VSS.n2388 4.5005
R23330 VSS.n2683 VSS.n2388 4.5005
R23331 VSS.n2685 VSS.n2388 4.5005
R23332 VSS.n2688 VSS.n2388 4.5005
R23333 VSS.n2690 VSS.n2388 4.5005
R23334 VSS.n2691 VSS.n2388 4.5005
R23335 VSS.n2693 VSS.n2388 4.5005
R23336 VSS.n2696 VSS.n2388 4.5005
R23337 VSS.n2698 VSS.n2388 4.5005
R23338 VSS.n2699 VSS.n2388 4.5005
R23339 VSS.n2701 VSS.n2388 4.5005
R23340 VSS.n2704 VSS.n2388 4.5005
R23341 VSS.n2706 VSS.n2388 4.5005
R23342 VSS.n2707 VSS.n2388 4.5005
R23343 VSS.n2709 VSS.n2388 4.5005
R23344 VSS.n2712 VSS.n2388 4.5005
R23345 VSS.n2714 VSS.n2388 4.5005
R23346 VSS.n2715 VSS.n2388 4.5005
R23347 VSS.n2717 VSS.n2388 4.5005
R23348 VSS.n2720 VSS.n2388 4.5005
R23349 VSS.n2722 VSS.n2388 4.5005
R23350 VSS.n2723 VSS.n2388 4.5005
R23351 VSS.n2725 VSS.n2388 4.5005
R23352 VSS.n2793 VSS.n2388 4.5005
R23353 VSS.n2859 VSS.n2388 4.5005
R23354 VSS.n3051 VSS.n2444 4.5005
R23355 VSS.n2444 VSS.n2351 4.5005
R23356 VSS.n2483 VSS.n2444 4.5005
R23357 VSS.n2484 VSS.n2444 4.5005
R23358 VSS.n2486 VSS.n2444 4.5005
R23359 VSS.n2489 VSS.n2444 4.5005
R23360 VSS.n2491 VSS.n2444 4.5005
R23361 VSS.n2492 VSS.n2444 4.5005
R23362 VSS.n2494 VSS.n2444 4.5005
R23363 VSS.n2497 VSS.n2444 4.5005
R23364 VSS.n2499 VSS.n2444 4.5005
R23365 VSS.n2500 VSS.n2444 4.5005
R23366 VSS.n2502 VSS.n2444 4.5005
R23367 VSS.n2505 VSS.n2444 4.5005
R23368 VSS.n2507 VSS.n2444 4.5005
R23369 VSS.n2508 VSS.n2444 4.5005
R23370 VSS.n2510 VSS.n2444 4.5005
R23371 VSS.n2513 VSS.n2444 4.5005
R23372 VSS.n2515 VSS.n2444 4.5005
R23373 VSS.n2516 VSS.n2444 4.5005
R23374 VSS.n2518 VSS.n2444 4.5005
R23375 VSS.n2521 VSS.n2444 4.5005
R23376 VSS.n2523 VSS.n2444 4.5005
R23377 VSS.n2524 VSS.n2444 4.5005
R23378 VSS.n2526 VSS.n2444 4.5005
R23379 VSS.n2529 VSS.n2444 4.5005
R23380 VSS.n2531 VSS.n2444 4.5005
R23381 VSS.n2532 VSS.n2444 4.5005
R23382 VSS.n2534 VSS.n2444 4.5005
R23383 VSS.n2537 VSS.n2444 4.5005
R23384 VSS.n2539 VSS.n2444 4.5005
R23385 VSS.n2540 VSS.n2444 4.5005
R23386 VSS.n2542 VSS.n2444 4.5005
R23387 VSS.n2545 VSS.n2444 4.5005
R23388 VSS.n2547 VSS.n2444 4.5005
R23389 VSS.n2548 VSS.n2444 4.5005
R23390 VSS.n2550 VSS.n2444 4.5005
R23391 VSS.n2553 VSS.n2444 4.5005
R23392 VSS.n2555 VSS.n2444 4.5005
R23393 VSS.n2556 VSS.n2444 4.5005
R23394 VSS.n2558 VSS.n2444 4.5005
R23395 VSS.n2561 VSS.n2444 4.5005
R23396 VSS.n2563 VSS.n2444 4.5005
R23397 VSS.n2564 VSS.n2444 4.5005
R23398 VSS.n2566 VSS.n2444 4.5005
R23399 VSS.n2569 VSS.n2444 4.5005
R23400 VSS.n2571 VSS.n2444 4.5005
R23401 VSS.n2572 VSS.n2444 4.5005
R23402 VSS.n2574 VSS.n2444 4.5005
R23403 VSS.n2577 VSS.n2444 4.5005
R23404 VSS.n2579 VSS.n2444 4.5005
R23405 VSS.n2580 VSS.n2444 4.5005
R23406 VSS.n2582 VSS.n2444 4.5005
R23407 VSS.n2585 VSS.n2444 4.5005
R23408 VSS.n2587 VSS.n2444 4.5005
R23409 VSS.n2588 VSS.n2444 4.5005
R23410 VSS.n2590 VSS.n2444 4.5005
R23411 VSS.n2593 VSS.n2444 4.5005
R23412 VSS.n2595 VSS.n2444 4.5005
R23413 VSS.n2596 VSS.n2444 4.5005
R23414 VSS.n2598 VSS.n2444 4.5005
R23415 VSS.n2601 VSS.n2444 4.5005
R23416 VSS.n2603 VSS.n2444 4.5005
R23417 VSS.n2604 VSS.n2444 4.5005
R23418 VSS.n2606 VSS.n2444 4.5005
R23419 VSS.n2609 VSS.n2444 4.5005
R23420 VSS.n2611 VSS.n2444 4.5005
R23421 VSS.n2612 VSS.n2444 4.5005
R23422 VSS.n2614 VSS.n2444 4.5005
R23423 VSS.n2617 VSS.n2444 4.5005
R23424 VSS.n2619 VSS.n2444 4.5005
R23425 VSS.n2620 VSS.n2444 4.5005
R23426 VSS.n2622 VSS.n2444 4.5005
R23427 VSS.n2625 VSS.n2444 4.5005
R23428 VSS.n2627 VSS.n2444 4.5005
R23429 VSS.n2628 VSS.n2444 4.5005
R23430 VSS.n2630 VSS.n2444 4.5005
R23431 VSS.n2633 VSS.n2444 4.5005
R23432 VSS.n2635 VSS.n2444 4.5005
R23433 VSS.n2636 VSS.n2444 4.5005
R23434 VSS.n2638 VSS.n2444 4.5005
R23435 VSS.n2640 VSS.n2444 4.5005
R23436 VSS.n2642 VSS.n2444 4.5005
R23437 VSS.n2643 VSS.n2444 4.5005
R23438 VSS.n2645 VSS.n2444 4.5005
R23439 VSS.n2648 VSS.n2444 4.5005
R23440 VSS.n2650 VSS.n2444 4.5005
R23441 VSS.n2651 VSS.n2444 4.5005
R23442 VSS.n2653 VSS.n2444 4.5005
R23443 VSS.n2656 VSS.n2444 4.5005
R23444 VSS.n2658 VSS.n2444 4.5005
R23445 VSS.n2659 VSS.n2444 4.5005
R23446 VSS.n2661 VSS.n2444 4.5005
R23447 VSS.n2664 VSS.n2444 4.5005
R23448 VSS.n2666 VSS.n2444 4.5005
R23449 VSS.n2667 VSS.n2444 4.5005
R23450 VSS.n2669 VSS.n2444 4.5005
R23451 VSS.n2672 VSS.n2444 4.5005
R23452 VSS.n2674 VSS.n2444 4.5005
R23453 VSS.n2675 VSS.n2444 4.5005
R23454 VSS.n2677 VSS.n2444 4.5005
R23455 VSS.n2680 VSS.n2444 4.5005
R23456 VSS.n2682 VSS.n2444 4.5005
R23457 VSS.n2683 VSS.n2444 4.5005
R23458 VSS.n2685 VSS.n2444 4.5005
R23459 VSS.n2688 VSS.n2444 4.5005
R23460 VSS.n2690 VSS.n2444 4.5005
R23461 VSS.n2691 VSS.n2444 4.5005
R23462 VSS.n2693 VSS.n2444 4.5005
R23463 VSS.n2696 VSS.n2444 4.5005
R23464 VSS.n2698 VSS.n2444 4.5005
R23465 VSS.n2699 VSS.n2444 4.5005
R23466 VSS.n2701 VSS.n2444 4.5005
R23467 VSS.n2704 VSS.n2444 4.5005
R23468 VSS.n2706 VSS.n2444 4.5005
R23469 VSS.n2707 VSS.n2444 4.5005
R23470 VSS.n2709 VSS.n2444 4.5005
R23471 VSS.n2712 VSS.n2444 4.5005
R23472 VSS.n2714 VSS.n2444 4.5005
R23473 VSS.n2715 VSS.n2444 4.5005
R23474 VSS.n2717 VSS.n2444 4.5005
R23475 VSS.n2720 VSS.n2444 4.5005
R23476 VSS.n2722 VSS.n2444 4.5005
R23477 VSS.n2723 VSS.n2444 4.5005
R23478 VSS.n2725 VSS.n2444 4.5005
R23479 VSS.n2793 VSS.n2444 4.5005
R23480 VSS.n2859 VSS.n2444 4.5005
R23481 VSS.n3051 VSS.n2387 4.5005
R23482 VSS.n2387 VSS.n2351 4.5005
R23483 VSS.n2483 VSS.n2387 4.5005
R23484 VSS.n2484 VSS.n2387 4.5005
R23485 VSS.n2486 VSS.n2387 4.5005
R23486 VSS.n2489 VSS.n2387 4.5005
R23487 VSS.n2491 VSS.n2387 4.5005
R23488 VSS.n2492 VSS.n2387 4.5005
R23489 VSS.n2494 VSS.n2387 4.5005
R23490 VSS.n2497 VSS.n2387 4.5005
R23491 VSS.n2499 VSS.n2387 4.5005
R23492 VSS.n2500 VSS.n2387 4.5005
R23493 VSS.n2502 VSS.n2387 4.5005
R23494 VSS.n2505 VSS.n2387 4.5005
R23495 VSS.n2507 VSS.n2387 4.5005
R23496 VSS.n2508 VSS.n2387 4.5005
R23497 VSS.n2510 VSS.n2387 4.5005
R23498 VSS.n2513 VSS.n2387 4.5005
R23499 VSS.n2515 VSS.n2387 4.5005
R23500 VSS.n2516 VSS.n2387 4.5005
R23501 VSS.n2518 VSS.n2387 4.5005
R23502 VSS.n2521 VSS.n2387 4.5005
R23503 VSS.n2523 VSS.n2387 4.5005
R23504 VSS.n2524 VSS.n2387 4.5005
R23505 VSS.n2526 VSS.n2387 4.5005
R23506 VSS.n2529 VSS.n2387 4.5005
R23507 VSS.n2531 VSS.n2387 4.5005
R23508 VSS.n2532 VSS.n2387 4.5005
R23509 VSS.n2534 VSS.n2387 4.5005
R23510 VSS.n2537 VSS.n2387 4.5005
R23511 VSS.n2539 VSS.n2387 4.5005
R23512 VSS.n2540 VSS.n2387 4.5005
R23513 VSS.n2542 VSS.n2387 4.5005
R23514 VSS.n2545 VSS.n2387 4.5005
R23515 VSS.n2547 VSS.n2387 4.5005
R23516 VSS.n2548 VSS.n2387 4.5005
R23517 VSS.n2550 VSS.n2387 4.5005
R23518 VSS.n2553 VSS.n2387 4.5005
R23519 VSS.n2555 VSS.n2387 4.5005
R23520 VSS.n2556 VSS.n2387 4.5005
R23521 VSS.n2558 VSS.n2387 4.5005
R23522 VSS.n2561 VSS.n2387 4.5005
R23523 VSS.n2563 VSS.n2387 4.5005
R23524 VSS.n2564 VSS.n2387 4.5005
R23525 VSS.n2566 VSS.n2387 4.5005
R23526 VSS.n2569 VSS.n2387 4.5005
R23527 VSS.n2571 VSS.n2387 4.5005
R23528 VSS.n2572 VSS.n2387 4.5005
R23529 VSS.n2574 VSS.n2387 4.5005
R23530 VSS.n2577 VSS.n2387 4.5005
R23531 VSS.n2579 VSS.n2387 4.5005
R23532 VSS.n2580 VSS.n2387 4.5005
R23533 VSS.n2582 VSS.n2387 4.5005
R23534 VSS.n2585 VSS.n2387 4.5005
R23535 VSS.n2587 VSS.n2387 4.5005
R23536 VSS.n2588 VSS.n2387 4.5005
R23537 VSS.n2590 VSS.n2387 4.5005
R23538 VSS.n2593 VSS.n2387 4.5005
R23539 VSS.n2595 VSS.n2387 4.5005
R23540 VSS.n2596 VSS.n2387 4.5005
R23541 VSS.n2598 VSS.n2387 4.5005
R23542 VSS.n2601 VSS.n2387 4.5005
R23543 VSS.n2603 VSS.n2387 4.5005
R23544 VSS.n2604 VSS.n2387 4.5005
R23545 VSS.n2606 VSS.n2387 4.5005
R23546 VSS.n2609 VSS.n2387 4.5005
R23547 VSS.n2611 VSS.n2387 4.5005
R23548 VSS.n2612 VSS.n2387 4.5005
R23549 VSS.n2614 VSS.n2387 4.5005
R23550 VSS.n2617 VSS.n2387 4.5005
R23551 VSS.n2619 VSS.n2387 4.5005
R23552 VSS.n2620 VSS.n2387 4.5005
R23553 VSS.n2622 VSS.n2387 4.5005
R23554 VSS.n2625 VSS.n2387 4.5005
R23555 VSS.n2627 VSS.n2387 4.5005
R23556 VSS.n2628 VSS.n2387 4.5005
R23557 VSS.n2630 VSS.n2387 4.5005
R23558 VSS.n2633 VSS.n2387 4.5005
R23559 VSS.n2635 VSS.n2387 4.5005
R23560 VSS.n2636 VSS.n2387 4.5005
R23561 VSS.n2638 VSS.n2387 4.5005
R23562 VSS.n2640 VSS.n2387 4.5005
R23563 VSS.n2642 VSS.n2387 4.5005
R23564 VSS.n2643 VSS.n2387 4.5005
R23565 VSS.n2645 VSS.n2387 4.5005
R23566 VSS.n2648 VSS.n2387 4.5005
R23567 VSS.n2650 VSS.n2387 4.5005
R23568 VSS.n2651 VSS.n2387 4.5005
R23569 VSS.n2653 VSS.n2387 4.5005
R23570 VSS.n2656 VSS.n2387 4.5005
R23571 VSS.n2658 VSS.n2387 4.5005
R23572 VSS.n2659 VSS.n2387 4.5005
R23573 VSS.n2661 VSS.n2387 4.5005
R23574 VSS.n2664 VSS.n2387 4.5005
R23575 VSS.n2666 VSS.n2387 4.5005
R23576 VSS.n2667 VSS.n2387 4.5005
R23577 VSS.n2669 VSS.n2387 4.5005
R23578 VSS.n2672 VSS.n2387 4.5005
R23579 VSS.n2674 VSS.n2387 4.5005
R23580 VSS.n2675 VSS.n2387 4.5005
R23581 VSS.n2677 VSS.n2387 4.5005
R23582 VSS.n2680 VSS.n2387 4.5005
R23583 VSS.n2682 VSS.n2387 4.5005
R23584 VSS.n2683 VSS.n2387 4.5005
R23585 VSS.n2685 VSS.n2387 4.5005
R23586 VSS.n2688 VSS.n2387 4.5005
R23587 VSS.n2690 VSS.n2387 4.5005
R23588 VSS.n2691 VSS.n2387 4.5005
R23589 VSS.n2693 VSS.n2387 4.5005
R23590 VSS.n2696 VSS.n2387 4.5005
R23591 VSS.n2698 VSS.n2387 4.5005
R23592 VSS.n2699 VSS.n2387 4.5005
R23593 VSS.n2701 VSS.n2387 4.5005
R23594 VSS.n2704 VSS.n2387 4.5005
R23595 VSS.n2706 VSS.n2387 4.5005
R23596 VSS.n2707 VSS.n2387 4.5005
R23597 VSS.n2709 VSS.n2387 4.5005
R23598 VSS.n2712 VSS.n2387 4.5005
R23599 VSS.n2714 VSS.n2387 4.5005
R23600 VSS.n2715 VSS.n2387 4.5005
R23601 VSS.n2717 VSS.n2387 4.5005
R23602 VSS.n2720 VSS.n2387 4.5005
R23603 VSS.n2722 VSS.n2387 4.5005
R23604 VSS.n2723 VSS.n2387 4.5005
R23605 VSS.n2725 VSS.n2387 4.5005
R23606 VSS.n2793 VSS.n2387 4.5005
R23607 VSS.n2859 VSS.n2387 4.5005
R23608 VSS.n3051 VSS.n2445 4.5005
R23609 VSS.n2445 VSS.n2351 4.5005
R23610 VSS.n2483 VSS.n2445 4.5005
R23611 VSS.n2484 VSS.n2445 4.5005
R23612 VSS.n2486 VSS.n2445 4.5005
R23613 VSS.n2489 VSS.n2445 4.5005
R23614 VSS.n2491 VSS.n2445 4.5005
R23615 VSS.n2492 VSS.n2445 4.5005
R23616 VSS.n2494 VSS.n2445 4.5005
R23617 VSS.n2497 VSS.n2445 4.5005
R23618 VSS.n2499 VSS.n2445 4.5005
R23619 VSS.n2500 VSS.n2445 4.5005
R23620 VSS.n2502 VSS.n2445 4.5005
R23621 VSS.n2505 VSS.n2445 4.5005
R23622 VSS.n2507 VSS.n2445 4.5005
R23623 VSS.n2508 VSS.n2445 4.5005
R23624 VSS.n2510 VSS.n2445 4.5005
R23625 VSS.n2513 VSS.n2445 4.5005
R23626 VSS.n2515 VSS.n2445 4.5005
R23627 VSS.n2516 VSS.n2445 4.5005
R23628 VSS.n2518 VSS.n2445 4.5005
R23629 VSS.n2521 VSS.n2445 4.5005
R23630 VSS.n2523 VSS.n2445 4.5005
R23631 VSS.n2524 VSS.n2445 4.5005
R23632 VSS.n2526 VSS.n2445 4.5005
R23633 VSS.n2529 VSS.n2445 4.5005
R23634 VSS.n2531 VSS.n2445 4.5005
R23635 VSS.n2532 VSS.n2445 4.5005
R23636 VSS.n2534 VSS.n2445 4.5005
R23637 VSS.n2537 VSS.n2445 4.5005
R23638 VSS.n2539 VSS.n2445 4.5005
R23639 VSS.n2540 VSS.n2445 4.5005
R23640 VSS.n2542 VSS.n2445 4.5005
R23641 VSS.n2545 VSS.n2445 4.5005
R23642 VSS.n2547 VSS.n2445 4.5005
R23643 VSS.n2548 VSS.n2445 4.5005
R23644 VSS.n2550 VSS.n2445 4.5005
R23645 VSS.n2553 VSS.n2445 4.5005
R23646 VSS.n2555 VSS.n2445 4.5005
R23647 VSS.n2556 VSS.n2445 4.5005
R23648 VSS.n2558 VSS.n2445 4.5005
R23649 VSS.n2561 VSS.n2445 4.5005
R23650 VSS.n2563 VSS.n2445 4.5005
R23651 VSS.n2564 VSS.n2445 4.5005
R23652 VSS.n2566 VSS.n2445 4.5005
R23653 VSS.n2569 VSS.n2445 4.5005
R23654 VSS.n2571 VSS.n2445 4.5005
R23655 VSS.n2572 VSS.n2445 4.5005
R23656 VSS.n2574 VSS.n2445 4.5005
R23657 VSS.n2577 VSS.n2445 4.5005
R23658 VSS.n2579 VSS.n2445 4.5005
R23659 VSS.n2580 VSS.n2445 4.5005
R23660 VSS.n2582 VSS.n2445 4.5005
R23661 VSS.n2585 VSS.n2445 4.5005
R23662 VSS.n2587 VSS.n2445 4.5005
R23663 VSS.n2588 VSS.n2445 4.5005
R23664 VSS.n2590 VSS.n2445 4.5005
R23665 VSS.n2593 VSS.n2445 4.5005
R23666 VSS.n2595 VSS.n2445 4.5005
R23667 VSS.n2596 VSS.n2445 4.5005
R23668 VSS.n2598 VSS.n2445 4.5005
R23669 VSS.n2601 VSS.n2445 4.5005
R23670 VSS.n2603 VSS.n2445 4.5005
R23671 VSS.n2604 VSS.n2445 4.5005
R23672 VSS.n2606 VSS.n2445 4.5005
R23673 VSS.n2609 VSS.n2445 4.5005
R23674 VSS.n2611 VSS.n2445 4.5005
R23675 VSS.n2612 VSS.n2445 4.5005
R23676 VSS.n2614 VSS.n2445 4.5005
R23677 VSS.n2617 VSS.n2445 4.5005
R23678 VSS.n2619 VSS.n2445 4.5005
R23679 VSS.n2620 VSS.n2445 4.5005
R23680 VSS.n2622 VSS.n2445 4.5005
R23681 VSS.n2625 VSS.n2445 4.5005
R23682 VSS.n2627 VSS.n2445 4.5005
R23683 VSS.n2628 VSS.n2445 4.5005
R23684 VSS.n2630 VSS.n2445 4.5005
R23685 VSS.n2633 VSS.n2445 4.5005
R23686 VSS.n2635 VSS.n2445 4.5005
R23687 VSS.n2636 VSS.n2445 4.5005
R23688 VSS.n2638 VSS.n2445 4.5005
R23689 VSS.n2640 VSS.n2445 4.5005
R23690 VSS.n2642 VSS.n2445 4.5005
R23691 VSS.n2643 VSS.n2445 4.5005
R23692 VSS.n2645 VSS.n2445 4.5005
R23693 VSS.n2648 VSS.n2445 4.5005
R23694 VSS.n2650 VSS.n2445 4.5005
R23695 VSS.n2651 VSS.n2445 4.5005
R23696 VSS.n2653 VSS.n2445 4.5005
R23697 VSS.n2656 VSS.n2445 4.5005
R23698 VSS.n2658 VSS.n2445 4.5005
R23699 VSS.n2659 VSS.n2445 4.5005
R23700 VSS.n2661 VSS.n2445 4.5005
R23701 VSS.n2664 VSS.n2445 4.5005
R23702 VSS.n2666 VSS.n2445 4.5005
R23703 VSS.n2667 VSS.n2445 4.5005
R23704 VSS.n2669 VSS.n2445 4.5005
R23705 VSS.n2672 VSS.n2445 4.5005
R23706 VSS.n2674 VSS.n2445 4.5005
R23707 VSS.n2675 VSS.n2445 4.5005
R23708 VSS.n2677 VSS.n2445 4.5005
R23709 VSS.n2680 VSS.n2445 4.5005
R23710 VSS.n2682 VSS.n2445 4.5005
R23711 VSS.n2683 VSS.n2445 4.5005
R23712 VSS.n2685 VSS.n2445 4.5005
R23713 VSS.n2688 VSS.n2445 4.5005
R23714 VSS.n2690 VSS.n2445 4.5005
R23715 VSS.n2691 VSS.n2445 4.5005
R23716 VSS.n2693 VSS.n2445 4.5005
R23717 VSS.n2696 VSS.n2445 4.5005
R23718 VSS.n2698 VSS.n2445 4.5005
R23719 VSS.n2699 VSS.n2445 4.5005
R23720 VSS.n2701 VSS.n2445 4.5005
R23721 VSS.n2704 VSS.n2445 4.5005
R23722 VSS.n2706 VSS.n2445 4.5005
R23723 VSS.n2707 VSS.n2445 4.5005
R23724 VSS.n2709 VSS.n2445 4.5005
R23725 VSS.n2712 VSS.n2445 4.5005
R23726 VSS.n2714 VSS.n2445 4.5005
R23727 VSS.n2715 VSS.n2445 4.5005
R23728 VSS.n2717 VSS.n2445 4.5005
R23729 VSS.n2720 VSS.n2445 4.5005
R23730 VSS.n2722 VSS.n2445 4.5005
R23731 VSS.n2723 VSS.n2445 4.5005
R23732 VSS.n2725 VSS.n2445 4.5005
R23733 VSS.n2793 VSS.n2445 4.5005
R23734 VSS.n2859 VSS.n2445 4.5005
R23735 VSS.n3051 VSS.n2386 4.5005
R23736 VSS.n2386 VSS.n2351 4.5005
R23737 VSS.n2483 VSS.n2386 4.5005
R23738 VSS.n2484 VSS.n2386 4.5005
R23739 VSS.n2486 VSS.n2386 4.5005
R23740 VSS.n2489 VSS.n2386 4.5005
R23741 VSS.n2491 VSS.n2386 4.5005
R23742 VSS.n2492 VSS.n2386 4.5005
R23743 VSS.n2494 VSS.n2386 4.5005
R23744 VSS.n2497 VSS.n2386 4.5005
R23745 VSS.n2499 VSS.n2386 4.5005
R23746 VSS.n2500 VSS.n2386 4.5005
R23747 VSS.n2502 VSS.n2386 4.5005
R23748 VSS.n2505 VSS.n2386 4.5005
R23749 VSS.n2507 VSS.n2386 4.5005
R23750 VSS.n2508 VSS.n2386 4.5005
R23751 VSS.n2510 VSS.n2386 4.5005
R23752 VSS.n2513 VSS.n2386 4.5005
R23753 VSS.n2515 VSS.n2386 4.5005
R23754 VSS.n2516 VSS.n2386 4.5005
R23755 VSS.n2518 VSS.n2386 4.5005
R23756 VSS.n2521 VSS.n2386 4.5005
R23757 VSS.n2523 VSS.n2386 4.5005
R23758 VSS.n2524 VSS.n2386 4.5005
R23759 VSS.n2526 VSS.n2386 4.5005
R23760 VSS.n2529 VSS.n2386 4.5005
R23761 VSS.n2531 VSS.n2386 4.5005
R23762 VSS.n2532 VSS.n2386 4.5005
R23763 VSS.n2534 VSS.n2386 4.5005
R23764 VSS.n2537 VSS.n2386 4.5005
R23765 VSS.n2539 VSS.n2386 4.5005
R23766 VSS.n2540 VSS.n2386 4.5005
R23767 VSS.n2542 VSS.n2386 4.5005
R23768 VSS.n2545 VSS.n2386 4.5005
R23769 VSS.n2547 VSS.n2386 4.5005
R23770 VSS.n2548 VSS.n2386 4.5005
R23771 VSS.n2550 VSS.n2386 4.5005
R23772 VSS.n2553 VSS.n2386 4.5005
R23773 VSS.n2555 VSS.n2386 4.5005
R23774 VSS.n2556 VSS.n2386 4.5005
R23775 VSS.n2558 VSS.n2386 4.5005
R23776 VSS.n2561 VSS.n2386 4.5005
R23777 VSS.n2563 VSS.n2386 4.5005
R23778 VSS.n2564 VSS.n2386 4.5005
R23779 VSS.n2566 VSS.n2386 4.5005
R23780 VSS.n2569 VSS.n2386 4.5005
R23781 VSS.n2571 VSS.n2386 4.5005
R23782 VSS.n2572 VSS.n2386 4.5005
R23783 VSS.n2574 VSS.n2386 4.5005
R23784 VSS.n2577 VSS.n2386 4.5005
R23785 VSS.n2579 VSS.n2386 4.5005
R23786 VSS.n2580 VSS.n2386 4.5005
R23787 VSS.n2582 VSS.n2386 4.5005
R23788 VSS.n2585 VSS.n2386 4.5005
R23789 VSS.n2587 VSS.n2386 4.5005
R23790 VSS.n2588 VSS.n2386 4.5005
R23791 VSS.n2590 VSS.n2386 4.5005
R23792 VSS.n2593 VSS.n2386 4.5005
R23793 VSS.n2595 VSS.n2386 4.5005
R23794 VSS.n2596 VSS.n2386 4.5005
R23795 VSS.n2598 VSS.n2386 4.5005
R23796 VSS.n2601 VSS.n2386 4.5005
R23797 VSS.n2603 VSS.n2386 4.5005
R23798 VSS.n2604 VSS.n2386 4.5005
R23799 VSS.n2606 VSS.n2386 4.5005
R23800 VSS.n2609 VSS.n2386 4.5005
R23801 VSS.n2611 VSS.n2386 4.5005
R23802 VSS.n2612 VSS.n2386 4.5005
R23803 VSS.n2614 VSS.n2386 4.5005
R23804 VSS.n2617 VSS.n2386 4.5005
R23805 VSS.n2619 VSS.n2386 4.5005
R23806 VSS.n2620 VSS.n2386 4.5005
R23807 VSS.n2622 VSS.n2386 4.5005
R23808 VSS.n2625 VSS.n2386 4.5005
R23809 VSS.n2627 VSS.n2386 4.5005
R23810 VSS.n2628 VSS.n2386 4.5005
R23811 VSS.n2630 VSS.n2386 4.5005
R23812 VSS.n2633 VSS.n2386 4.5005
R23813 VSS.n2635 VSS.n2386 4.5005
R23814 VSS.n2636 VSS.n2386 4.5005
R23815 VSS.n2638 VSS.n2386 4.5005
R23816 VSS.n2640 VSS.n2386 4.5005
R23817 VSS.n2642 VSS.n2386 4.5005
R23818 VSS.n2643 VSS.n2386 4.5005
R23819 VSS.n2645 VSS.n2386 4.5005
R23820 VSS.n2648 VSS.n2386 4.5005
R23821 VSS.n2650 VSS.n2386 4.5005
R23822 VSS.n2651 VSS.n2386 4.5005
R23823 VSS.n2653 VSS.n2386 4.5005
R23824 VSS.n2656 VSS.n2386 4.5005
R23825 VSS.n2658 VSS.n2386 4.5005
R23826 VSS.n2659 VSS.n2386 4.5005
R23827 VSS.n2661 VSS.n2386 4.5005
R23828 VSS.n2664 VSS.n2386 4.5005
R23829 VSS.n2666 VSS.n2386 4.5005
R23830 VSS.n2667 VSS.n2386 4.5005
R23831 VSS.n2669 VSS.n2386 4.5005
R23832 VSS.n2672 VSS.n2386 4.5005
R23833 VSS.n2674 VSS.n2386 4.5005
R23834 VSS.n2675 VSS.n2386 4.5005
R23835 VSS.n2677 VSS.n2386 4.5005
R23836 VSS.n2680 VSS.n2386 4.5005
R23837 VSS.n2682 VSS.n2386 4.5005
R23838 VSS.n2683 VSS.n2386 4.5005
R23839 VSS.n2685 VSS.n2386 4.5005
R23840 VSS.n2688 VSS.n2386 4.5005
R23841 VSS.n2690 VSS.n2386 4.5005
R23842 VSS.n2691 VSS.n2386 4.5005
R23843 VSS.n2693 VSS.n2386 4.5005
R23844 VSS.n2696 VSS.n2386 4.5005
R23845 VSS.n2698 VSS.n2386 4.5005
R23846 VSS.n2699 VSS.n2386 4.5005
R23847 VSS.n2701 VSS.n2386 4.5005
R23848 VSS.n2704 VSS.n2386 4.5005
R23849 VSS.n2706 VSS.n2386 4.5005
R23850 VSS.n2707 VSS.n2386 4.5005
R23851 VSS.n2709 VSS.n2386 4.5005
R23852 VSS.n2712 VSS.n2386 4.5005
R23853 VSS.n2714 VSS.n2386 4.5005
R23854 VSS.n2715 VSS.n2386 4.5005
R23855 VSS.n2717 VSS.n2386 4.5005
R23856 VSS.n2720 VSS.n2386 4.5005
R23857 VSS.n2722 VSS.n2386 4.5005
R23858 VSS.n2723 VSS.n2386 4.5005
R23859 VSS.n2725 VSS.n2386 4.5005
R23860 VSS.n2793 VSS.n2386 4.5005
R23861 VSS.n2859 VSS.n2386 4.5005
R23862 VSS.n3051 VSS.n2446 4.5005
R23863 VSS.n2446 VSS.n2351 4.5005
R23864 VSS.n2483 VSS.n2446 4.5005
R23865 VSS.n2484 VSS.n2446 4.5005
R23866 VSS.n2486 VSS.n2446 4.5005
R23867 VSS.n2489 VSS.n2446 4.5005
R23868 VSS.n2491 VSS.n2446 4.5005
R23869 VSS.n2492 VSS.n2446 4.5005
R23870 VSS.n2494 VSS.n2446 4.5005
R23871 VSS.n2497 VSS.n2446 4.5005
R23872 VSS.n2499 VSS.n2446 4.5005
R23873 VSS.n2500 VSS.n2446 4.5005
R23874 VSS.n2502 VSS.n2446 4.5005
R23875 VSS.n2505 VSS.n2446 4.5005
R23876 VSS.n2507 VSS.n2446 4.5005
R23877 VSS.n2508 VSS.n2446 4.5005
R23878 VSS.n2510 VSS.n2446 4.5005
R23879 VSS.n2513 VSS.n2446 4.5005
R23880 VSS.n2515 VSS.n2446 4.5005
R23881 VSS.n2516 VSS.n2446 4.5005
R23882 VSS.n2518 VSS.n2446 4.5005
R23883 VSS.n2521 VSS.n2446 4.5005
R23884 VSS.n2523 VSS.n2446 4.5005
R23885 VSS.n2524 VSS.n2446 4.5005
R23886 VSS.n2526 VSS.n2446 4.5005
R23887 VSS.n2529 VSS.n2446 4.5005
R23888 VSS.n2531 VSS.n2446 4.5005
R23889 VSS.n2532 VSS.n2446 4.5005
R23890 VSS.n2534 VSS.n2446 4.5005
R23891 VSS.n2537 VSS.n2446 4.5005
R23892 VSS.n2539 VSS.n2446 4.5005
R23893 VSS.n2540 VSS.n2446 4.5005
R23894 VSS.n2542 VSS.n2446 4.5005
R23895 VSS.n2545 VSS.n2446 4.5005
R23896 VSS.n2547 VSS.n2446 4.5005
R23897 VSS.n2548 VSS.n2446 4.5005
R23898 VSS.n2550 VSS.n2446 4.5005
R23899 VSS.n2553 VSS.n2446 4.5005
R23900 VSS.n2555 VSS.n2446 4.5005
R23901 VSS.n2556 VSS.n2446 4.5005
R23902 VSS.n2558 VSS.n2446 4.5005
R23903 VSS.n2561 VSS.n2446 4.5005
R23904 VSS.n2563 VSS.n2446 4.5005
R23905 VSS.n2564 VSS.n2446 4.5005
R23906 VSS.n2566 VSS.n2446 4.5005
R23907 VSS.n2569 VSS.n2446 4.5005
R23908 VSS.n2571 VSS.n2446 4.5005
R23909 VSS.n2572 VSS.n2446 4.5005
R23910 VSS.n2574 VSS.n2446 4.5005
R23911 VSS.n2577 VSS.n2446 4.5005
R23912 VSS.n2579 VSS.n2446 4.5005
R23913 VSS.n2580 VSS.n2446 4.5005
R23914 VSS.n2582 VSS.n2446 4.5005
R23915 VSS.n2585 VSS.n2446 4.5005
R23916 VSS.n2587 VSS.n2446 4.5005
R23917 VSS.n2588 VSS.n2446 4.5005
R23918 VSS.n2590 VSS.n2446 4.5005
R23919 VSS.n2593 VSS.n2446 4.5005
R23920 VSS.n2595 VSS.n2446 4.5005
R23921 VSS.n2596 VSS.n2446 4.5005
R23922 VSS.n2598 VSS.n2446 4.5005
R23923 VSS.n2601 VSS.n2446 4.5005
R23924 VSS.n2603 VSS.n2446 4.5005
R23925 VSS.n2604 VSS.n2446 4.5005
R23926 VSS.n2606 VSS.n2446 4.5005
R23927 VSS.n2609 VSS.n2446 4.5005
R23928 VSS.n2611 VSS.n2446 4.5005
R23929 VSS.n2612 VSS.n2446 4.5005
R23930 VSS.n2614 VSS.n2446 4.5005
R23931 VSS.n2617 VSS.n2446 4.5005
R23932 VSS.n2619 VSS.n2446 4.5005
R23933 VSS.n2620 VSS.n2446 4.5005
R23934 VSS.n2622 VSS.n2446 4.5005
R23935 VSS.n2625 VSS.n2446 4.5005
R23936 VSS.n2627 VSS.n2446 4.5005
R23937 VSS.n2628 VSS.n2446 4.5005
R23938 VSS.n2630 VSS.n2446 4.5005
R23939 VSS.n2633 VSS.n2446 4.5005
R23940 VSS.n2635 VSS.n2446 4.5005
R23941 VSS.n2636 VSS.n2446 4.5005
R23942 VSS.n2638 VSS.n2446 4.5005
R23943 VSS.n2640 VSS.n2446 4.5005
R23944 VSS.n2642 VSS.n2446 4.5005
R23945 VSS.n2643 VSS.n2446 4.5005
R23946 VSS.n2645 VSS.n2446 4.5005
R23947 VSS.n2648 VSS.n2446 4.5005
R23948 VSS.n2650 VSS.n2446 4.5005
R23949 VSS.n2651 VSS.n2446 4.5005
R23950 VSS.n2653 VSS.n2446 4.5005
R23951 VSS.n2656 VSS.n2446 4.5005
R23952 VSS.n2658 VSS.n2446 4.5005
R23953 VSS.n2659 VSS.n2446 4.5005
R23954 VSS.n2661 VSS.n2446 4.5005
R23955 VSS.n2664 VSS.n2446 4.5005
R23956 VSS.n2666 VSS.n2446 4.5005
R23957 VSS.n2667 VSS.n2446 4.5005
R23958 VSS.n2669 VSS.n2446 4.5005
R23959 VSS.n2672 VSS.n2446 4.5005
R23960 VSS.n2674 VSS.n2446 4.5005
R23961 VSS.n2675 VSS.n2446 4.5005
R23962 VSS.n2677 VSS.n2446 4.5005
R23963 VSS.n2680 VSS.n2446 4.5005
R23964 VSS.n2682 VSS.n2446 4.5005
R23965 VSS.n2683 VSS.n2446 4.5005
R23966 VSS.n2685 VSS.n2446 4.5005
R23967 VSS.n2688 VSS.n2446 4.5005
R23968 VSS.n2690 VSS.n2446 4.5005
R23969 VSS.n2691 VSS.n2446 4.5005
R23970 VSS.n2693 VSS.n2446 4.5005
R23971 VSS.n2696 VSS.n2446 4.5005
R23972 VSS.n2698 VSS.n2446 4.5005
R23973 VSS.n2699 VSS.n2446 4.5005
R23974 VSS.n2701 VSS.n2446 4.5005
R23975 VSS.n2704 VSS.n2446 4.5005
R23976 VSS.n2706 VSS.n2446 4.5005
R23977 VSS.n2707 VSS.n2446 4.5005
R23978 VSS.n2709 VSS.n2446 4.5005
R23979 VSS.n2712 VSS.n2446 4.5005
R23980 VSS.n2714 VSS.n2446 4.5005
R23981 VSS.n2715 VSS.n2446 4.5005
R23982 VSS.n2717 VSS.n2446 4.5005
R23983 VSS.n2720 VSS.n2446 4.5005
R23984 VSS.n2722 VSS.n2446 4.5005
R23985 VSS.n2723 VSS.n2446 4.5005
R23986 VSS.n2725 VSS.n2446 4.5005
R23987 VSS.n2793 VSS.n2446 4.5005
R23988 VSS.n2859 VSS.n2446 4.5005
R23989 VSS.n3051 VSS.n2385 4.5005
R23990 VSS.n2385 VSS.n2351 4.5005
R23991 VSS.n2483 VSS.n2385 4.5005
R23992 VSS.n2484 VSS.n2385 4.5005
R23993 VSS.n2486 VSS.n2385 4.5005
R23994 VSS.n2489 VSS.n2385 4.5005
R23995 VSS.n2491 VSS.n2385 4.5005
R23996 VSS.n2492 VSS.n2385 4.5005
R23997 VSS.n2494 VSS.n2385 4.5005
R23998 VSS.n2497 VSS.n2385 4.5005
R23999 VSS.n2499 VSS.n2385 4.5005
R24000 VSS.n2500 VSS.n2385 4.5005
R24001 VSS.n2502 VSS.n2385 4.5005
R24002 VSS.n2505 VSS.n2385 4.5005
R24003 VSS.n2507 VSS.n2385 4.5005
R24004 VSS.n2508 VSS.n2385 4.5005
R24005 VSS.n2510 VSS.n2385 4.5005
R24006 VSS.n2513 VSS.n2385 4.5005
R24007 VSS.n2515 VSS.n2385 4.5005
R24008 VSS.n2516 VSS.n2385 4.5005
R24009 VSS.n2518 VSS.n2385 4.5005
R24010 VSS.n2521 VSS.n2385 4.5005
R24011 VSS.n2523 VSS.n2385 4.5005
R24012 VSS.n2524 VSS.n2385 4.5005
R24013 VSS.n2526 VSS.n2385 4.5005
R24014 VSS.n2529 VSS.n2385 4.5005
R24015 VSS.n2531 VSS.n2385 4.5005
R24016 VSS.n2532 VSS.n2385 4.5005
R24017 VSS.n2534 VSS.n2385 4.5005
R24018 VSS.n2537 VSS.n2385 4.5005
R24019 VSS.n2539 VSS.n2385 4.5005
R24020 VSS.n2540 VSS.n2385 4.5005
R24021 VSS.n2542 VSS.n2385 4.5005
R24022 VSS.n2545 VSS.n2385 4.5005
R24023 VSS.n2547 VSS.n2385 4.5005
R24024 VSS.n2548 VSS.n2385 4.5005
R24025 VSS.n2550 VSS.n2385 4.5005
R24026 VSS.n2553 VSS.n2385 4.5005
R24027 VSS.n2555 VSS.n2385 4.5005
R24028 VSS.n2556 VSS.n2385 4.5005
R24029 VSS.n2558 VSS.n2385 4.5005
R24030 VSS.n2561 VSS.n2385 4.5005
R24031 VSS.n2563 VSS.n2385 4.5005
R24032 VSS.n2564 VSS.n2385 4.5005
R24033 VSS.n2566 VSS.n2385 4.5005
R24034 VSS.n2569 VSS.n2385 4.5005
R24035 VSS.n2571 VSS.n2385 4.5005
R24036 VSS.n2572 VSS.n2385 4.5005
R24037 VSS.n2574 VSS.n2385 4.5005
R24038 VSS.n2577 VSS.n2385 4.5005
R24039 VSS.n2579 VSS.n2385 4.5005
R24040 VSS.n2580 VSS.n2385 4.5005
R24041 VSS.n2582 VSS.n2385 4.5005
R24042 VSS.n2585 VSS.n2385 4.5005
R24043 VSS.n2587 VSS.n2385 4.5005
R24044 VSS.n2588 VSS.n2385 4.5005
R24045 VSS.n2590 VSS.n2385 4.5005
R24046 VSS.n2593 VSS.n2385 4.5005
R24047 VSS.n2595 VSS.n2385 4.5005
R24048 VSS.n2596 VSS.n2385 4.5005
R24049 VSS.n2598 VSS.n2385 4.5005
R24050 VSS.n2601 VSS.n2385 4.5005
R24051 VSS.n2603 VSS.n2385 4.5005
R24052 VSS.n2604 VSS.n2385 4.5005
R24053 VSS.n2606 VSS.n2385 4.5005
R24054 VSS.n2609 VSS.n2385 4.5005
R24055 VSS.n2611 VSS.n2385 4.5005
R24056 VSS.n2612 VSS.n2385 4.5005
R24057 VSS.n2614 VSS.n2385 4.5005
R24058 VSS.n2617 VSS.n2385 4.5005
R24059 VSS.n2619 VSS.n2385 4.5005
R24060 VSS.n2620 VSS.n2385 4.5005
R24061 VSS.n2622 VSS.n2385 4.5005
R24062 VSS.n2625 VSS.n2385 4.5005
R24063 VSS.n2627 VSS.n2385 4.5005
R24064 VSS.n2628 VSS.n2385 4.5005
R24065 VSS.n2630 VSS.n2385 4.5005
R24066 VSS.n2633 VSS.n2385 4.5005
R24067 VSS.n2635 VSS.n2385 4.5005
R24068 VSS.n2636 VSS.n2385 4.5005
R24069 VSS.n2638 VSS.n2385 4.5005
R24070 VSS.n2640 VSS.n2385 4.5005
R24071 VSS.n2642 VSS.n2385 4.5005
R24072 VSS.n2643 VSS.n2385 4.5005
R24073 VSS.n2645 VSS.n2385 4.5005
R24074 VSS.n2648 VSS.n2385 4.5005
R24075 VSS.n2650 VSS.n2385 4.5005
R24076 VSS.n2651 VSS.n2385 4.5005
R24077 VSS.n2653 VSS.n2385 4.5005
R24078 VSS.n2656 VSS.n2385 4.5005
R24079 VSS.n2658 VSS.n2385 4.5005
R24080 VSS.n2659 VSS.n2385 4.5005
R24081 VSS.n2661 VSS.n2385 4.5005
R24082 VSS.n2664 VSS.n2385 4.5005
R24083 VSS.n2666 VSS.n2385 4.5005
R24084 VSS.n2667 VSS.n2385 4.5005
R24085 VSS.n2669 VSS.n2385 4.5005
R24086 VSS.n2672 VSS.n2385 4.5005
R24087 VSS.n2674 VSS.n2385 4.5005
R24088 VSS.n2675 VSS.n2385 4.5005
R24089 VSS.n2677 VSS.n2385 4.5005
R24090 VSS.n2680 VSS.n2385 4.5005
R24091 VSS.n2682 VSS.n2385 4.5005
R24092 VSS.n2683 VSS.n2385 4.5005
R24093 VSS.n2685 VSS.n2385 4.5005
R24094 VSS.n2688 VSS.n2385 4.5005
R24095 VSS.n2690 VSS.n2385 4.5005
R24096 VSS.n2691 VSS.n2385 4.5005
R24097 VSS.n2693 VSS.n2385 4.5005
R24098 VSS.n2696 VSS.n2385 4.5005
R24099 VSS.n2698 VSS.n2385 4.5005
R24100 VSS.n2699 VSS.n2385 4.5005
R24101 VSS.n2701 VSS.n2385 4.5005
R24102 VSS.n2704 VSS.n2385 4.5005
R24103 VSS.n2706 VSS.n2385 4.5005
R24104 VSS.n2707 VSS.n2385 4.5005
R24105 VSS.n2709 VSS.n2385 4.5005
R24106 VSS.n2712 VSS.n2385 4.5005
R24107 VSS.n2714 VSS.n2385 4.5005
R24108 VSS.n2715 VSS.n2385 4.5005
R24109 VSS.n2717 VSS.n2385 4.5005
R24110 VSS.n2720 VSS.n2385 4.5005
R24111 VSS.n2722 VSS.n2385 4.5005
R24112 VSS.n2723 VSS.n2385 4.5005
R24113 VSS.n2725 VSS.n2385 4.5005
R24114 VSS.n2793 VSS.n2385 4.5005
R24115 VSS.n2859 VSS.n2385 4.5005
R24116 VSS.n3051 VSS.n2447 4.5005
R24117 VSS.n2447 VSS.n2351 4.5005
R24118 VSS.n2483 VSS.n2447 4.5005
R24119 VSS.n2484 VSS.n2447 4.5005
R24120 VSS.n2486 VSS.n2447 4.5005
R24121 VSS.n2489 VSS.n2447 4.5005
R24122 VSS.n2491 VSS.n2447 4.5005
R24123 VSS.n2492 VSS.n2447 4.5005
R24124 VSS.n2494 VSS.n2447 4.5005
R24125 VSS.n2497 VSS.n2447 4.5005
R24126 VSS.n2499 VSS.n2447 4.5005
R24127 VSS.n2500 VSS.n2447 4.5005
R24128 VSS.n2502 VSS.n2447 4.5005
R24129 VSS.n2505 VSS.n2447 4.5005
R24130 VSS.n2507 VSS.n2447 4.5005
R24131 VSS.n2508 VSS.n2447 4.5005
R24132 VSS.n2510 VSS.n2447 4.5005
R24133 VSS.n2513 VSS.n2447 4.5005
R24134 VSS.n2515 VSS.n2447 4.5005
R24135 VSS.n2516 VSS.n2447 4.5005
R24136 VSS.n2518 VSS.n2447 4.5005
R24137 VSS.n2521 VSS.n2447 4.5005
R24138 VSS.n2523 VSS.n2447 4.5005
R24139 VSS.n2524 VSS.n2447 4.5005
R24140 VSS.n2526 VSS.n2447 4.5005
R24141 VSS.n2529 VSS.n2447 4.5005
R24142 VSS.n2531 VSS.n2447 4.5005
R24143 VSS.n2532 VSS.n2447 4.5005
R24144 VSS.n2534 VSS.n2447 4.5005
R24145 VSS.n2537 VSS.n2447 4.5005
R24146 VSS.n2539 VSS.n2447 4.5005
R24147 VSS.n2540 VSS.n2447 4.5005
R24148 VSS.n2542 VSS.n2447 4.5005
R24149 VSS.n2545 VSS.n2447 4.5005
R24150 VSS.n2547 VSS.n2447 4.5005
R24151 VSS.n2548 VSS.n2447 4.5005
R24152 VSS.n2550 VSS.n2447 4.5005
R24153 VSS.n2553 VSS.n2447 4.5005
R24154 VSS.n2555 VSS.n2447 4.5005
R24155 VSS.n2556 VSS.n2447 4.5005
R24156 VSS.n2558 VSS.n2447 4.5005
R24157 VSS.n2561 VSS.n2447 4.5005
R24158 VSS.n2563 VSS.n2447 4.5005
R24159 VSS.n2564 VSS.n2447 4.5005
R24160 VSS.n2566 VSS.n2447 4.5005
R24161 VSS.n2569 VSS.n2447 4.5005
R24162 VSS.n2571 VSS.n2447 4.5005
R24163 VSS.n2572 VSS.n2447 4.5005
R24164 VSS.n2574 VSS.n2447 4.5005
R24165 VSS.n2577 VSS.n2447 4.5005
R24166 VSS.n2579 VSS.n2447 4.5005
R24167 VSS.n2580 VSS.n2447 4.5005
R24168 VSS.n2582 VSS.n2447 4.5005
R24169 VSS.n2585 VSS.n2447 4.5005
R24170 VSS.n2587 VSS.n2447 4.5005
R24171 VSS.n2588 VSS.n2447 4.5005
R24172 VSS.n2590 VSS.n2447 4.5005
R24173 VSS.n2593 VSS.n2447 4.5005
R24174 VSS.n2595 VSS.n2447 4.5005
R24175 VSS.n2596 VSS.n2447 4.5005
R24176 VSS.n2598 VSS.n2447 4.5005
R24177 VSS.n2601 VSS.n2447 4.5005
R24178 VSS.n2603 VSS.n2447 4.5005
R24179 VSS.n2604 VSS.n2447 4.5005
R24180 VSS.n2606 VSS.n2447 4.5005
R24181 VSS.n2609 VSS.n2447 4.5005
R24182 VSS.n2611 VSS.n2447 4.5005
R24183 VSS.n2612 VSS.n2447 4.5005
R24184 VSS.n2614 VSS.n2447 4.5005
R24185 VSS.n2617 VSS.n2447 4.5005
R24186 VSS.n2619 VSS.n2447 4.5005
R24187 VSS.n2620 VSS.n2447 4.5005
R24188 VSS.n2622 VSS.n2447 4.5005
R24189 VSS.n2625 VSS.n2447 4.5005
R24190 VSS.n2627 VSS.n2447 4.5005
R24191 VSS.n2628 VSS.n2447 4.5005
R24192 VSS.n2630 VSS.n2447 4.5005
R24193 VSS.n2633 VSS.n2447 4.5005
R24194 VSS.n2635 VSS.n2447 4.5005
R24195 VSS.n2636 VSS.n2447 4.5005
R24196 VSS.n2638 VSS.n2447 4.5005
R24197 VSS.n2640 VSS.n2447 4.5005
R24198 VSS.n2642 VSS.n2447 4.5005
R24199 VSS.n2643 VSS.n2447 4.5005
R24200 VSS.n2645 VSS.n2447 4.5005
R24201 VSS.n2648 VSS.n2447 4.5005
R24202 VSS.n2650 VSS.n2447 4.5005
R24203 VSS.n2651 VSS.n2447 4.5005
R24204 VSS.n2653 VSS.n2447 4.5005
R24205 VSS.n2656 VSS.n2447 4.5005
R24206 VSS.n2658 VSS.n2447 4.5005
R24207 VSS.n2659 VSS.n2447 4.5005
R24208 VSS.n2661 VSS.n2447 4.5005
R24209 VSS.n2664 VSS.n2447 4.5005
R24210 VSS.n2666 VSS.n2447 4.5005
R24211 VSS.n2667 VSS.n2447 4.5005
R24212 VSS.n2669 VSS.n2447 4.5005
R24213 VSS.n2672 VSS.n2447 4.5005
R24214 VSS.n2674 VSS.n2447 4.5005
R24215 VSS.n2675 VSS.n2447 4.5005
R24216 VSS.n2677 VSS.n2447 4.5005
R24217 VSS.n2680 VSS.n2447 4.5005
R24218 VSS.n2682 VSS.n2447 4.5005
R24219 VSS.n2683 VSS.n2447 4.5005
R24220 VSS.n2685 VSS.n2447 4.5005
R24221 VSS.n2688 VSS.n2447 4.5005
R24222 VSS.n2690 VSS.n2447 4.5005
R24223 VSS.n2691 VSS.n2447 4.5005
R24224 VSS.n2693 VSS.n2447 4.5005
R24225 VSS.n2696 VSS.n2447 4.5005
R24226 VSS.n2698 VSS.n2447 4.5005
R24227 VSS.n2699 VSS.n2447 4.5005
R24228 VSS.n2701 VSS.n2447 4.5005
R24229 VSS.n2704 VSS.n2447 4.5005
R24230 VSS.n2706 VSS.n2447 4.5005
R24231 VSS.n2707 VSS.n2447 4.5005
R24232 VSS.n2709 VSS.n2447 4.5005
R24233 VSS.n2712 VSS.n2447 4.5005
R24234 VSS.n2714 VSS.n2447 4.5005
R24235 VSS.n2715 VSS.n2447 4.5005
R24236 VSS.n2717 VSS.n2447 4.5005
R24237 VSS.n2720 VSS.n2447 4.5005
R24238 VSS.n2722 VSS.n2447 4.5005
R24239 VSS.n2723 VSS.n2447 4.5005
R24240 VSS.n2725 VSS.n2447 4.5005
R24241 VSS.n2793 VSS.n2447 4.5005
R24242 VSS.n2859 VSS.n2447 4.5005
R24243 VSS.n3051 VSS.n2384 4.5005
R24244 VSS.n2384 VSS.n2351 4.5005
R24245 VSS.n2483 VSS.n2384 4.5005
R24246 VSS.n2484 VSS.n2384 4.5005
R24247 VSS.n2486 VSS.n2384 4.5005
R24248 VSS.n2489 VSS.n2384 4.5005
R24249 VSS.n2491 VSS.n2384 4.5005
R24250 VSS.n2492 VSS.n2384 4.5005
R24251 VSS.n2494 VSS.n2384 4.5005
R24252 VSS.n2497 VSS.n2384 4.5005
R24253 VSS.n2499 VSS.n2384 4.5005
R24254 VSS.n2500 VSS.n2384 4.5005
R24255 VSS.n2502 VSS.n2384 4.5005
R24256 VSS.n2505 VSS.n2384 4.5005
R24257 VSS.n2507 VSS.n2384 4.5005
R24258 VSS.n2508 VSS.n2384 4.5005
R24259 VSS.n2510 VSS.n2384 4.5005
R24260 VSS.n2513 VSS.n2384 4.5005
R24261 VSS.n2515 VSS.n2384 4.5005
R24262 VSS.n2516 VSS.n2384 4.5005
R24263 VSS.n2518 VSS.n2384 4.5005
R24264 VSS.n2521 VSS.n2384 4.5005
R24265 VSS.n2523 VSS.n2384 4.5005
R24266 VSS.n2524 VSS.n2384 4.5005
R24267 VSS.n2526 VSS.n2384 4.5005
R24268 VSS.n2529 VSS.n2384 4.5005
R24269 VSS.n2531 VSS.n2384 4.5005
R24270 VSS.n2532 VSS.n2384 4.5005
R24271 VSS.n2534 VSS.n2384 4.5005
R24272 VSS.n2537 VSS.n2384 4.5005
R24273 VSS.n2539 VSS.n2384 4.5005
R24274 VSS.n2540 VSS.n2384 4.5005
R24275 VSS.n2542 VSS.n2384 4.5005
R24276 VSS.n2545 VSS.n2384 4.5005
R24277 VSS.n2547 VSS.n2384 4.5005
R24278 VSS.n2548 VSS.n2384 4.5005
R24279 VSS.n2550 VSS.n2384 4.5005
R24280 VSS.n2553 VSS.n2384 4.5005
R24281 VSS.n2555 VSS.n2384 4.5005
R24282 VSS.n2556 VSS.n2384 4.5005
R24283 VSS.n2558 VSS.n2384 4.5005
R24284 VSS.n2561 VSS.n2384 4.5005
R24285 VSS.n2563 VSS.n2384 4.5005
R24286 VSS.n2564 VSS.n2384 4.5005
R24287 VSS.n2566 VSS.n2384 4.5005
R24288 VSS.n2569 VSS.n2384 4.5005
R24289 VSS.n2571 VSS.n2384 4.5005
R24290 VSS.n2572 VSS.n2384 4.5005
R24291 VSS.n2574 VSS.n2384 4.5005
R24292 VSS.n2577 VSS.n2384 4.5005
R24293 VSS.n2579 VSS.n2384 4.5005
R24294 VSS.n2580 VSS.n2384 4.5005
R24295 VSS.n2582 VSS.n2384 4.5005
R24296 VSS.n2585 VSS.n2384 4.5005
R24297 VSS.n2587 VSS.n2384 4.5005
R24298 VSS.n2588 VSS.n2384 4.5005
R24299 VSS.n2590 VSS.n2384 4.5005
R24300 VSS.n2593 VSS.n2384 4.5005
R24301 VSS.n2595 VSS.n2384 4.5005
R24302 VSS.n2596 VSS.n2384 4.5005
R24303 VSS.n2598 VSS.n2384 4.5005
R24304 VSS.n2601 VSS.n2384 4.5005
R24305 VSS.n2603 VSS.n2384 4.5005
R24306 VSS.n2604 VSS.n2384 4.5005
R24307 VSS.n2606 VSS.n2384 4.5005
R24308 VSS.n2609 VSS.n2384 4.5005
R24309 VSS.n2611 VSS.n2384 4.5005
R24310 VSS.n2612 VSS.n2384 4.5005
R24311 VSS.n2614 VSS.n2384 4.5005
R24312 VSS.n2617 VSS.n2384 4.5005
R24313 VSS.n2619 VSS.n2384 4.5005
R24314 VSS.n2620 VSS.n2384 4.5005
R24315 VSS.n2622 VSS.n2384 4.5005
R24316 VSS.n2625 VSS.n2384 4.5005
R24317 VSS.n2627 VSS.n2384 4.5005
R24318 VSS.n2628 VSS.n2384 4.5005
R24319 VSS.n2630 VSS.n2384 4.5005
R24320 VSS.n2633 VSS.n2384 4.5005
R24321 VSS.n2635 VSS.n2384 4.5005
R24322 VSS.n2636 VSS.n2384 4.5005
R24323 VSS.n2638 VSS.n2384 4.5005
R24324 VSS.n2640 VSS.n2384 4.5005
R24325 VSS.n2642 VSS.n2384 4.5005
R24326 VSS.n2643 VSS.n2384 4.5005
R24327 VSS.n2645 VSS.n2384 4.5005
R24328 VSS.n2648 VSS.n2384 4.5005
R24329 VSS.n2650 VSS.n2384 4.5005
R24330 VSS.n2651 VSS.n2384 4.5005
R24331 VSS.n2653 VSS.n2384 4.5005
R24332 VSS.n2656 VSS.n2384 4.5005
R24333 VSS.n2658 VSS.n2384 4.5005
R24334 VSS.n2659 VSS.n2384 4.5005
R24335 VSS.n2661 VSS.n2384 4.5005
R24336 VSS.n2664 VSS.n2384 4.5005
R24337 VSS.n2666 VSS.n2384 4.5005
R24338 VSS.n2667 VSS.n2384 4.5005
R24339 VSS.n2669 VSS.n2384 4.5005
R24340 VSS.n2672 VSS.n2384 4.5005
R24341 VSS.n2674 VSS.n2384 4.5005
R24342 VSS.n2675 VSS.n2384 4.5005
R24343 VSS.n2677 VSS.n2384 4.5005
R24344 VSS.n2680 VSS.n2384 4.5005
R24345 VSS.n2682 VSS.n2384 4.5005
R24346 VSS.n2683 VSS.n2384 4.5005
R24347 VSS.n2685 VSS.n2384 4.5005
R24348 VSS.n2688 VSS.n2384 4.5005
R24349 VSS.n2690 VSS.n2384 4.5005
R24350 VSS.n2691 VSS.n2384 4.5005
R24351 VSS.n2693 VSS.n2384 4.5005
R24352 VSS.n2696 VSS.n2384 4.5005
R24353 VSS.n2698 VSS.n2384 4.5005
R24354 VSS.n2699 VSS.n2384 4.5005
R24355 VSS.n2701 VSS.n2384 4.5005
R24356 VSS.n2704 VSS.n2384 4.5005
R24357 VSS.n2706 VSS.n2384 4.5005
R24358 VSS.n2707 VSS.n2384 4.5005
R24359 VSS.n2709 VSS.n2384 4.5005
R24360 VSS.n2712 VSS.n2384 4.5005
R24361 VSS.n2714 VSS.n2384 4.5005
R24362 VSS.n2715 VSS.n2384 4.5005
R24363 VSS.n2717 VSS.n2384 4.5005
R24364 VSS.n2720 VSS.n2384 4.5005
R24365 VSS.n2722 VSS.n2384 4.5005
R24366 VSS.n2723 VSS.n2384 4.5005
R24367 VSS.n2725 VSS.n2384 4.5005
R24368 VSS.n2793 VSS.n2384 4.5005
R24369 VSS.n2859 VSS.n2384 4.5005
R24370 VSS.n3051 VSS.n2448 4.5005
R24371 VSS.n2448 VSS.n2351 4.5005
R24372 VSS.n2483 VSS.n2448 4.5005
R24373 VSS.n2484 VSS.n2448 4.5005
R24374 VSS.n2486 VSS.n2448 4.5005
R24375 VSS.n2489 VSS.n2448 4.5005
R24376 VSS.n2491 VSS.n2448 4.5005
R24377 VSS.n2492 VSS.n2448 4.5005
R24378 VSS.n2494 VSS.n2448 4.5005
R24379 VSS.n2497 VSS.n2448 4.5005
R24380 VSS.n2499 VSS.n2448 4.5005
R24381 VSS.n2500 VSS.n2448 4.5005
R24382 VSS.n2502 VSS.n2448 4.5005
R24383 VSS.n2505 VSS.n2448 4.5005
R24384 VSS.n2507 VSS.n2448 4.5005
R24385 VSS.n2508 VSS.n2448 4.5005
R24386 VSS.n2510 VSS.n2448 4.5005
R24387 VSS.n2513 VSS.n2448 4.5005
R24388 VSS.n2515 VSS.n2448 4.5005
R24389 VSS.n2516 VSS.n2448 4.5005
R24390 VSS.n2518 VSS.n2448 4.5005
R24391 VSS.n2521 VSS.n2448 4.5005
R24392 VSS.n2523 VSS.n2448 4.5005
R24393 VSS.n2524 VSS.n2448 4.5005
R24394 VSS.n2526 VSS.n2448 4.5005
R24395 VSS.n2529 VSS.n2448 4.5005
R24396 VSS.n2531 VSS.n2448 4.5005
R24397 VSS.n2532 VSS.n2448 4.5005
R24398 VSS.n2534 VSS.n2448 4.5005
R24399 VSS.n2537 VSS.n2448 4.5005
R24400 VSS.n2539 VSS.n2448 4.5005
R24401 VSS.n2540 VSS.n2448 4.5005
R24402 VSS.n2542 VSS.n2448 4.5005
R24403 VSS.n2545 VSS.n2448 4.5005
R24404 VSS.n2547 VSS.n2448 4.5005
R24405 VSS.n2548 VSS.n2448 4.5005
R24406 VSS.n2550 VSS.n2448 4.5005
R24407 VSS.n2553 VSS.n2448 4.5005
R24408 VSS.n2555 VSS.n2448 4.5005
R24409 VSS.n2556 VSS.n2448 4.5005
R24410 VSS.n2558 VSS.n2448 4.5005
R24411 VSS.n2561 VSS.n2448 4.5005
R24412 VSS.n2563 VSS.n2448 4.5005
R24413 VSS.n2564 VSS.n2448 4.5005
R24414 VSS.n2566 VSS.n2448 4.5005
R24415 VSS.n2569 VSS.n2448 4.5005
R24416 VSS.n2571 VSS.n2448 4.5005
R24417 VSS.n2572 VSS.n2448 4.5005
R24418 VSS.n2574 VSS.n2448 4.5005
R24419 VSS.n2577 VSS.n2448 4.5005
R24420 VSS.n2579 VSS.n2448 4.5005
R24421 VSS.n2580 VSS.n2448 4.5005
R24422 VSS.n2582 VSS.n2448 4.5005
R24423 VSS.n2585 VSS.n2448 4.5005
R24424 VSS.n2587 VSS.n2448 4.5005
R24425 VSS.n2588 VSS.n2448 4.5005
R24426 VSS.n2590 VSS.n2448 4.5005
R24427 VSS.n2593 VSS.n2448 4.5005
R24428 VSS.n2595 VSS.n2448 4.5005
R24429 VSS.n2596 VSS.n2448 4.5005
R24430 VSS.n2598 VSS.n2448 4.5005
R24431 VSS.n2601 VSS.n2448 4.5005
R24432 VSS.n2603 VSS.n2448 4.5005
R24433 VSS.n2604 VSS.n2448 4.5005
R24434 VSS.n2606 VSS.n2448 4.5005
R24435 VSS.n2609 VSS.n2448 4.5005
R24436 VSS.n2611 VSS.n2448 4.5005
R24437 VSS.n2612 VSS.n2448 4.5005
R24438 VSS.n2614 VSS.n2448 4.5005
R24439 VSS.n2617 VSS.n2448 4.5005
R24440 VSS.n2619 VSS.n2448 4.5005
R24441 VSS.n2620 VSS.n2448 4.5005
R24442 VSS.n2622 VSS.n2448 4.5005
R24443 VSS.n2625 VSS.n2448 4.5005
R24444 VSS.n2627 VSS.n2448 4.5005
R24445 VSS.n2628 VSS.n2448 4.5005
R24446 VSS.n2630 VSS.n2448 4.5005
R24447 VSS.n2633 VSS.n2448 4.5005
R24448 VSS.n2635 VSS.n2448 4.5005
R24449 VSS.n2636 VSS.n2448 4.5005
R24450 VSS.n2638 VSS.n2448 4.5005
R24451 VSS.n2640 VSS.n2448 4.5005
R24452 VSS.n2642 VSS.n2448 4.5005
R24453 VSS.n2643 VSS.n2448 4.5005
R24454 VSS.n2645 VSS.n2448 4.5005
R24455 VSS.n2648 VSS.n2448 4.5005
R24456 VSS.n2650 VSS.n2448 4.5005
R24457 VSS.n2651 VSS.n2448 4.5005
R24458 VSS.n2653 VSS.n2448 4.5005
R24459 VSS.n2656 VSS.n2448 4.5005
R24460 VSS.n2658 VSS.n2448 4.5005
R24461 VSS.n2659 VSS.n2448 4.5005
R24462 VSS.n2661 VSS.n2448 4.5005
R24463 VSS.n2664 VSS.n2448 4.5005
R24464 VSS.n2666 VSS.n2448 4.5005
R24465 VSS.n2667 VSS.n2448 4.5005
R24466 VSS.n2669 VSS.n2448 4.5005
R24467 VSS.n2672 VSS.n2448 4.5005
R24468 VSS.n2674 VSS.n2448 4.5005
R24469 VSS.n2675 VSS.n2448 4.5005
R24470 VSS.n2677 VSS.n2448 4.5005
R24471 VSS.n2680 VSS.n2448 4.5005
R24472 VSS.n2682 VSS.n2448 4.5005
R24473 VSS.n2683 VSS.n2448 4.5005
R24474 VSS.n2685 VSS.n2448 4.5005
R24475 VSS.n2688 VSS.n2448 4.5005
R24476 VSS.n2690 VSS.n2448 4.5005
R24477 VSS.n2691 VSS.n2448 4.5005
R24478 VSS.n2693 VSS.n2448 4.5005
R24479 VSS.n2696 VSS.n2448 4.5005
R24480 VSS.n2698 VSS.n2448 4.5005
R24481 VSS.n2699 VSS.n2448 4.5005
R24482 VSS.n2701 VSS.n2448 4.5005
R24483 VSS.n2704 VSS.n2448 4.5005
R24484 VSS.n2706 VSS.n2448 4.5005
R24485 VSS.n2707 VSS.n2448 4.5005
R24486 VSS.n2709 VSS.n2448 4.5005
R24487 VSS.n2712 VSS.n2448 4.5005
R24488 VSS.n2714 VSS.n2448 4.5005
R24489 VSS.n2715 VSS.n2448 4.5005
R24490 VSS.n2717 VSS.n2448 4.5005
R24491 VSS.n2720 VSS.n2448 4.5005
R24492 VSS.n2722 VSS.n2448 4.5005
R24493 VSS.n2723 VSS.n2448 4.5005
R24494 VSS.n2725 VSS.n2448 4.5005
R24495 VSS.n2793 VSS.n2448 4.5005
R24496 VSS.n2859 VSS.n2448 4.5005
R24497 VSS.n3051 VSS.n2383 4.5005
R24498 VSS.n2383 VSS.n2351 4.5005
R24499 VSS.n2483 VSS.n2383 4.5005
R24500 VSS.n2484 VSS.n2383 4.5005
R24501 VSS.n2486 VSS.n2383 4.5005
R24502 VSS.n2489 VSS.n2383 4.5005
R24503 VSS.n2491 VSS.n2383 4.5005
R24504 VSS.n2492 VSS.n2383 4.5005
R24505 VSS.n2494 VSS.n2383 4.5005
R24506 VSS.n2497 VSS.n2383 4.5005
R24507 VSS.n2499 VSS.n2383 4.5005
R24508 VSS.n2500 VSS.n2383 4.5005
R24509 VSS.n2502 VSS.n2383 4.5005
R24510 VSS.n2505 VSS.n2383 4.5005
R24511 VSS.n2507 VSS.n2383 4.5005
R24512 VSS.n2508 VSS.n2383 4.5005
R24513 VSS.n2510 VSS.n2383 4.5005
R24514 VSS.n2513 VSS.n2383 4.5005
R24515 VSS.n2515 VSS.n2383 4.5005
R24516 VSS.n2516 VSS.n2383 4.5005
R24517 VSS.n2518 VSS.n2383 4.5005
R24518 VSS.n2521 VSS.n2383 4.5005
R24519 VSS.n2523 VSS.n2383 4.5005
R24520 VSS.n2524 VSS.n2383 4.5005
R24521 VSS.n2526 VSS.n2383 4.5005
R24522 VSS.n2529 VSS.n2383 4.5005
R24523 VSS.n2531 VSS.n2383 4.5005
R24524 VSS.n2532 VSS.n2383 4.5005
R24525 VSS.n2534 VSS.n2383 4.5005
R24526 VSS.n2537 VSS.n2383 4.5005
R24527 VSS.n2539 VSS.n2383 4.5005
R24528 VSS.n2540 VSS.n2383 4.5005
R24529 VSS.n2542 VSS.n2383 4.5005
R24530 VSS.n2545 VSS.n2383 4.5005
R24531 VSS.n2547 VSS.n2383 4.5005
R24532 VSS.n2548 VSS.n2383 4.5005
R24533 VSS.n2550 VSS.n2383 4.5005
R24534 VSS.n2553 VSS.n2383 4.5005
R24535 VSS.n2555 VSS.n2383 4.5005
R24536 VSS.n2556 VSS.n2383 4.5005
R24537 VSS.n2558 VSS.n2383 4.5005
R24538 VSS.n2561 VSS.n2383 4.5005
R24539 VSS.n2563 VSS.n2383 4.5005
R24540 VSS.n2564 VSS.n2383 4.5005
R24541 VSS.n2566 VSS.n2383 4.5005
R24542 VSS.n2569 VSS.n2383 4.5005
R24543 VSS.n2571 VSS.n2383 4.5005
R24544 VSS.n2572 VSS.n2383 4.5005
R24545 VSS.n2574 VSS.n2383 4.5005
R24546 VSS.n2577 VSS.n2383 4.5005
R24547 VSS.n2579 VSS.n2383 4.5005
R24548 VSS.n2580 VSS.n2383 4.5005
R24549 VSS.n2582 VSS.n2383 4.5005
R24550 VSS.n2585 VSS.n2383 4.5005
R24551 VSS.n2587 VSS.n2383 4.5005
R24552 VSS.n2588 VSS.n2383 4.5005
R24553 VSS.n2590 VSS.n2383 4.5005
R24554 VSS.n2593 VSS.n2383 4.5005
R24555 VSS.n2595 VSS.n2383 4.5005
R24556 VSS.n2596 VSS.n2383 4.5005
R24557 VSS.n2598 VSS.n2383 4.5005
R24558 VSS.n2601 VSS.n2383 4.5005
R24559 VSS.n2603 VSS.n2383 4.5005
R24560 VSS.n2604 VSS.n2383 4.5005
R24561 VSS.n2606 VSS.n2383 4.5005
R24562 VSS.n2609 VSS.n2383 4.5005
R24563 VSS.n2611 VSS.n2383 4.5005
R24564 VSS.n2612 VSS.n2383 4.5005
R24565 VSS.n2614 VSS.n2383 4.5005
R24566 VSS.n2617 VSS.n2383 4.5005
R24567 VSS.n2619 VSS.n2383 4.5005
R24568 VSS.n2620 VSS.n2383 4.5005
R24569 VSS.n2622 VSS.n2383 4.5005
R24570 VSS.n2625 VSS.n2383 4.5005
R24571 VSS.n2627 VSS.n2383 4.5005
R24572 VSS.n2628 VSS.n2383 4.5005
R24573 VSS.n2630 VSS.n2383 4.5005
R24574 VSS.n2633 VSS.n2383 4.5005
R24575 VSS.n2635 VSS.n2383 4.5005
R24576 VSS.n2636 VSS.n2383 4.5005
R24577 VSS.n2638 VSS.n2383 4.5005
R24578 VSS.n2640 VSS.n2383 4.5005
R24579 VSS.n2642 VSS.n2383 4.5005
R24580 VSS.n2643 VSS.n2383 4.5005
R24581 VSS.n2645 VSS.n2383 4.5005
R24582 VSS.n2648 VSS.n2383 4.5005
R24583 VSS.n2650 VSS.n2383 4.5005
R24584 VSS.n2651 VSS.n2383 4.5005
R24585 VSS.n2653 VSS.n2383 4.5005
R24586 VSS.n2656 VSS.n2383 4.5005
R24587 VSS.n2658 VSS.n2383 4.5005
R24588 VSS.n2659 VSS.n2383 4.5005
R24589 VSS.n2661 VSS.n2383 4.5005
R24590 VSS.n2664 VSS.n2383 4.5005
R24591 VSS.n2666 VSS.n2383 4.5005
R24592 VSS.n2667 VSS.n2383 4.5005
R24593 VSS.n2669 VSS.n2383 4.5005
R24594 VSS.n2672 VSS.n2383 4.5005
R24595 VSS.n2674 VSS.n2383 4.5005
R24596 VSS.n2675 VSS.n2383 4.5005
R24597 VSS.n2677 VSS.n2383 4.5005
R24598 VSS.n2680 VSS.n2383 4.5005
R24599 VSS.n2682 VSS.n2383 4.5005
R24600 VSS.n2683 VSS.n2383 4.5005
R24601 VSS.n2685 VSS.n2383 4.5005
R24602 VSS.n2688 VSS.n2383 4.5005
R24603 VSS.n2690 VSS.n2383 4.5005
R24604 VSS.n2691 VSS.n2383 4.5005
R24605 VSS.n2693 VSS.n2383 4.5005
R24606 VSS.n2696 VSS.n2383 4.5005
R24607 VSS.n2698 VSS.n2383 4.5005
R24608 VSS.n2699 VSS.n2383 4.5005
R24609 VSS.n2701 VSS.n2383 4.5005
R24610 VSS.n2704 VSS.n2383 4.5005
R24611 VSS.n2706 VSS.n2383 4.5005
R24612 VSS.n2707 VSS.n2383 4.5005
R24613 VSS.n2709 VSS.n2383 4.5005
R24614 VSS.n2712 VSS.n2383 4.5005
R24615 VSS.n2714 VSS.n2383 4.5005
R24616 VSS.n2715 VSS.n2383 4.5005
R24617 VSS.n2717 VSS.n2383 4.5005
R24618 VSS.n2720 VSS.n2383 4.5005
R24619 VSS.n2722 VSS.n2383 4.5005
R24620 VSS.n2723 VSS.n2383 4.5005
R24621 VSS.n2725 VSS.n2383 4.5005
R24622 VSS.n2793 VSS.n2383 4.5005
R24623 VSS.n2859 VSS.n2383 4.5005
R24624 VSS.n3051 VSS.n2449 4.5005
R24625 VSS.n2449 VSS.n2351 4.5005
R24626 VSS.n2483 VSS.n2449 4.5005
R24627 VSS.n2484 VSS.n2449 4.5005
R24628 VSS.n2486 VSS.n2449 4.5005
R24629 VSS.n2489 VSS.n2449 4.5005
R24630 VSS.n2491 VSS.n2449 4.5005
R24631 VSS.n2492 VSS.n2449 4.5005
R24632 VSS.n2494 VSS.n2449 4.5005
R24633 VSS.n2497 VSS.n2449 4.5005
R24634 VSS.n2499 VSS.n2449 4.5005
R24635 VSS.n2500 VSS.n2449 4.5005
R24636 VSS.n2502 VSS.n2449 4.5005
R24637 VSS.n2505 VSS.n2449 4.5005
R24638 VSS.n2507 VSS.n2449 4.5005
R24639 VSS.n2508 VSS.n2449 4.5005
R24640 VSS.n2510 VSS.n2449 4.5005
R24641 VSS.n2513 VSS.n2449 4.5005
R24642 VSS.n2515 VSS.n2449 4.5005
R24643 VSS.n2516 VSS.n2449 4.5005
R24644 VSS.n2518 VSS.n2449 4.5005
R24645 VSS.n2521 VSS.n2449 4.5005
R24646 VSS.n2523 VSS.n2449 4.5005
R24647 VSS.n2524 VSS.n2449 4.5005
R24648 VSS.n2526 VSS.n2449 4.5005
R24649 VSS.n2529 VSS.n2449 4.5005
R24650 VSS.n2531 VSS.n2449 4.5005
R24651 VSS.n2532 VSS.n2449 4.5005
R24652 VSS.n2534 VSS.n2449 4.5005
R24653 VSS.n2537 VSS.n2449 4.5005
R24654 VSS.n2539 VSS.n2449 4.5005
R24655 VSS.n2540 VSS.n2449 4.5005
R24656 VSS.n2542 VSS.n2449 4.5005
R24657 VSS.n2545 VSS.n2449 4.5005
R24658 VSS.n2547 VSS.n2449 4.5005
R24659 VSS.n2548 VSS.n2449 4.5005
R24660 VSS.n2550 VSS.n2449 4.5005
R24661 VSS.n2553 VSS.n2449 4.5005
R24662 VSS.n2555 VSS.n2449 4.5005
R24663 VSS.n2556 VSS.n2449 4.5005
R24664 VSS.n2558 VSS.n2449 4.5005
R24665 VSS.n2561 VSS.n2449 4.5005
R24666 VSS.n2563 VSS.n2449 4.5005
R24667 VSS.n2564 VSS.n2449 4.5005
R24668 VSS.n2566 VSS.n2449 4.5005
R24669 VSS.n2569 VSS.n2449 4.5005
R24670 VSS.n2571 VSS.n2449 4.5005
R24671 VSS.n2572 VSS.n2449 4.5005
R24672 VSS.n2574 VSS.n2449 4.5005
R24673 VSS.n2577 VSS.n2449 4.5005
R24674 VSS.n2579 VSS.n2449 4.5005
R24675 VSS.n2580 VSS.n2449 4.5005
R24676 VSS.n2582 VSS.n2449 4.5005
R24677 VSS.n2585 VSS.n2449 4.5005
R24678 VSS.n2587 VSS.n2449 4.5005
R24679 VSS.n2588 VSS.n2449 4.5005
R24680 VSS.n2590 VSS.n2449 4.5005
R24681 VSS.n2593 VSS.n2449 4.5005
R24682 VSS.n2595 VSS.n2449 4.5005
R24683 VSS.n2596 VSS.n2449 4.5005
R24684 VSS.n2598 VSS.n2449 4.5005
R24685 VSS.n2601 VSS.n2449 4.5005
R24686 VSS.n2603 VSS.n2449 4.5005
R24687 VSS.n2604 VSS.n2449 4.5005
R24688 VSS.n2606 VSS.n2449 4.5005
R24689 VSS.n2609 VSS.n2449 4.5005
R24690 VSS.n2611 VSS.n2449 4.5005
R24691 VSS.n2612 VSS.n2449 4.5005
R24692 VSS.n2614 VSS.n2449 4.5005
R24693 VSS.n2617 VSS.n2449 4.5005
R24694 VSS.n2619 VSS.n2449 4.5005
R24695 VSS.n2620 VSS.n2449 4.5005
R24696 VSS.n2622 VSS.n2449 4.5005
R24697 VSS.n2625 VSS.n2449 4.5005
R24698 VSS.n2627 VSS.n2449 4.5005
R24699 VSS.n2628 VSS.n2449 4.5005
R24700 VSS.n2630 VSS.n2449 4.5005
R24701 VSS.n2633 VSS.n2449 4.5005
R24702 VSS.n2635 VSS.n2449 4.5005
R24703 VSS.n2636 VSS.n2449 4.5005
R24704 VSS.n2638 VSS.n2449 4.5005
R24705 VSS.n2640 VSS.n2449 4.5005
R24706 VSS.n2642 VSS.n2449 4.5005
R24707 VSS.n2643 VSS.n2449 4.5005
R24708 VSS.n2645 VSS.n2449 4.5005
R24709 VSS.n2648 VSS.n2449 4.5005
R24710 VSS.n2650 VSS.n2449 4.5005
R24711 VSS.n2651 VSS.n2449 4.5005
R24712 VSS.n2653 VSS.n2449 4.5005
R24713 VSS.n2656 VSS.n2449 4.5005
R24714 VSS.n2658 VSS.n2449 4.5005
R24715 VSS.n2659 VSS.n2449 4.5005
R24716 VSS.n2661 VSS.n2449 4.5005
R24717 VSS.n2664 VSS.n2449 4.5005
R24718 VSS.n2666 VSS.n2449 4.5005
R24719 VSS.n2667 VSS.n2449 4.5005
R24720 VSS.n2669 VSS.n2449 4.5005
R24721 VSS.n2672 VSS.n2449 4.5005
R24722 VSS.n2674 VSS.n2449 4.5005
R24723 VSS.n2675 VSS.n2449 4.5005
R24724 VSS.n2677 VSS.n2449 4.5005
R24725 VSS.n2680 VSS.n2449 4.5005
R24726 VSS.n2682 VSS.n2449 4.5005
R24727 VSS.n2683 VSS.n2449 4.5005
R24728 VSS.n2685 VSS.n2449 4.5005
R24729 VSS.n2688 VSS.n2449 4.5005
R24730 VSS.n2690 VSS.n2449 4.5005
R24731 VSS.n2691 VSS.n2449 4.5005
R24732 VSS.n2693 VSS.n2449 4.5005
R24733 VSS.n2696 VSS.n2449 4.5005
R24734 VSS.n2698 VSS.n2449 4.5005
R24735 VSS.n2699 VSS.n2449 4.5005
R24736 VSS.n2701 VSS.n2449 4.5005
R24737 VSS.n2704 VSS.n2449 4.5005
R24738 VSS.n2706 VSS.n2449 4.5005
R24739 VSS.n2707 VSS.n2449 4.5005
R24740 VSS.n2709 VSS.n2449 4.5005
R24741 VSS.n2712 VSS.n2449 4.5005
R24742 VSS.n2714 VSS.n2449 4.5005
R24743 VSS.n2715 VSS.n2449 4.5005
R24744 VSS.n2717 VSS.n2449 4.5005
R24745 VSS.n2720 VSS.n2449 4.5005
R24746 VSS.n2722 VSS.n2449 4.5005
R24747 VSS.n2723 VSS.n2449 4.5005
R24748 VSS.n2725 VSS.n2449 4.5005
R24749 VSS.n2793 VSS.n2449 4.5005
R24750 VSS.n2859 VSS.n2449 4.5005
R24751 VSS.n3051 VSS.n2382 4.5005
R24752 VSS.n2382 VSS.n2351 4.5005
R24753 VSS.n2483 VSS.n2382 4.5005
R24754 VSS.n2484 VSS.n2382 4.5005
R24755 VSS.n2486 VSS.n2382 4.5005
R24756 VSS.n2489 VSS.n2382 4.5005
R24757 VSS.n2491 VSS.n2382 4.5005
R24758 VSS.n2492 VSS.n2382 4.5005
R24759 VSS.n2494 VSS.n2382 4.5005
R24760 VSS.n2497 VSS.n2382 4.5005
R24761 VSS.n2499 VSS.n2382 4.5005
R24762 VSS.n2500 VSS.n2382 4.5005
R24763 VSS.n2502 VSS.n2382 4.5005
R24764 VSS.n2505 VSS.n2382 4.5005
R24765 VSS.n2507 VSS.n2382 4.5005
R24766 VSS.n2508 VSS.n2382 4.5005
R24767 VSS.n2510 VSS.n2382 4.5005
R24768 VSS.n2513 VSS.n2382 4.5005
R24769 VSS.n2515 VSS.n2382 4.5005
R24770 VSS.n2516 VSS.n2382 4.5005
R24771 VSS.n2518 VSS.n2382 4.5005
R24772 VSS.n2521 VSS.n2382 4.5005
R24773 VSS.n2523 VSS.n2382 4.5005
R24774 VSS.n2524 VSS.n2382 4.5005
R24775 VSS.n2526 VSS.n2382 4.5005
R24776 VSS.n2529 VSS.n2382 4.5005
R24777 VSS.n2531 VSS.n2382 4.5005
R24778 VSS.n2532 VSS.n2382 4.5005
R24779 VSS.n2534 VSS.n2382 4.5005
R24780 VSS.n2537 VSS.n2382 4.5005
R24781 VSS.n2539 VSS.n2382 4.5005
R24782 VSS.n2540 VSS.n2382 4.5005
R24783 VSS.n2542 VSS.n2382 4.5005
R24784 VSS.n2545 VSS.n2382 4.5005
R24785 VSS.n2547 VSS.n2382 4.5005
R24786 VSS.n2548 VSS.n2382 4.5005
R24787 VSS.n2550 VSS.n2382 4.5005
R24788 VSS.n2553 VSS.n2382 4.5005
R24789 VSS.n2555 VSS.n2382 4.5005
R24790 VSS.n2556 VSS.n2382 4.5005
R24791 VSS.n2558 VSS.n2382 4.5005
R24792 VSS.n2561 VSS.n2382 4.5005
R24793 VSS.n2563 VSS.n2382 4.5005
R24794 VSS.n2564 VSS.n2382 4.5005
R24795 VSS.n2566 VSS.n2382 4.5005
R24796 VSS.n2569 VSS.n2382 4.5005
R24797 VSS.n2571 VSS.n2382 4.5005
R24798 VSS.n2572 VSS.n2382 4.5005
R24799 VSS.n2574 VSS.n2382 4.5005
R24800 VSS.n2577 VSS.n2382 4.5005
R24801 VSS.n2579 VSS.n2382 4.5005
R24802 VSS.n2580 VSS.n2382 4.5005
R24803 VSS.n2582 VSS.n2382 4.5005
R24804 VSS.n2585 VSS.n2382 4.5005
R24805 VSS.n2587 VSS.n2382 4.5005
R24806 VSS.n2588 VSS.n2382 4.5005
R24807 VSS.n2590 VSS.n2382 4.5005
R24808 VSS.n2593 VSS.n2382 4.5005
R24809 VSS.n2595 VSS.n2382 4.5005
R24810 VSS.n2596 VSS.n2382 4.5005
R24811 VSS.n2598 VSS.n2382 4.5005
R24812 VSS.n2601 VSS.n2382 4.5005
R24813 VSS.n2603 VSS.n2382 4.5005
R24814 VSS.n2604 VSS.n2382 4.5005
R24815 VSS.n2606 VSS.n2382 4.5005
R24816 VSS.n2609 VSS.n2382 4.5005
R24817 VSS.n2611 VSS.n2382 4.5005
R24818 VSS.n2612 VSS.n2382 4.5005
R24819 VSS.n2614 VSS.n2382 4.5005
R24820 VSS.n2617 VSS.n2382 4.5005
R24821 VSS.n2619 VSS.n2382 4.5005
R24822 VSS.n2620 VSS.n2382 4.5005
R24823 VSS.n2622 VSS.n2382 4.5005
R24824 VSS.n2625 VSS.n2382 4.5005
R24825 VSS.n2627 VSS.n2382 4.5005
R24826 VSS.n2628 VSS.n2382 4.5005
R24827 VSS.n2630 VSS.n2382 4.5005
R24828 VSS.n2633 VSS.n2382 4.5005
R24829 VSS.n2635 VSS.n2382 4.5005
R24830 VSS.n2636 VSS.n2382 4.5005
R24831 VSS.n2638 VSS.n2382 4.5005
R24832 VSS.n2640 VSS.n2382 4.5005
R24833 VSS.n2642 VSS.n2382 4.5005
R24834 VSS.n2643 VSS.n2382 4.5005
R24835 VSS.n2645 VSS.n2382 4.5005
R24836 VSS.n2648 VSS.n2382 4.5005
R24837 VSS.n2650 VSS.n2382 4.5005
R24838 VSS.n2651 VSS.n2382 4.5005
R24839 VSS.n2653 VSS.n2382 4.5005
R24840 VSS.n2656 VSS.n2382 4.5005
R24841 VSS.n2658 VSS.n2382 4.5005
R24842 VSS.n2659 VSS.n2382 4.5005
R24843 VSS.n2661 VSS.n2382 4.5005
R24844 VSS.n2664 VSS.n2382 4.5005
R24845 VSS.n2666 VSS.n2382 4.5005
R24846 VSS.n2667 VSS.n2382 4.5005
R24847 VSS.n2669 VSS.n2382 4.5005
R24848 VSS.n2672 VSS.n2382 4.5005
R24849 VSS.n2674 VSS.n2382 4.5005
R24850 VSS.n2675 VSS.n2382 4.5005
R24851 VSS.n2677 VSS.n2382 4.5005
R24852 VSS.n2680 VSS.n2382 4.5005
R24853 VSS.n2682 VSS.n2382 4.5005
R24854 VSS.n2683 VSS.n2382 4.5005
R24855 VSS.n2685 VSS.n2382 4.5005
R24856 VSS.n2688 VSS.n2382 4.5005
R24857 VSS.n2690 VSS.n2382 4.5005
R24858 VSS.n2691 VSS.n2382 4.5005
R24859 VSS.n2693 VSS.n2382 4.5005
R24860 VSS.n2696 VSS.n2382 4.5005
R24861 VSS.n2698 VSS.n2382 4.5005
R24862 VSS.n2699 VSS.n2382 4.5005
R24863 VSS.n2701 VSS.n2382 4.5005
R24864 VSS.n2704 VSS.n2382 4.5005
R24865 VSS.n2706 VSS.n2382 4.5005
R24866 VSS.n2707 VSS.n2382 4.5005
R24867 VSS.n2709 VSS.n2382 4.5005
R24868 VSS.n2712 VSS.n2382 4.5005
R24869 VSS.n2714 VSS.n2382 4.5005
R24870 VSS.n2715 VSS.n2382 4.5005
R24871 VSS.n2717 VSS.n2382 4.5005
R24872 VSS.n2720 VSS.n2382 4.5005
R24873 VSS.n2722 VSS.n2382 4.5005
R24874 VSS.n2723 VSS.n2382 4.5005
R24875 VSS.n2725 VSS.n2382 4.5005
R24876 VSS.n2793 VSS.n2382 4.5005
R24877 VSS.n2859 VSS.n2382 4.5005
R24878 VSS.n3051 VSS.n2450 4.5005
R24879 VSS.n2450 VSS.n2351 4.5005
R24880 VSS.n2483 VSS.n2450 4.5005
R24881 VSS.n2484 VSS.n2450 4.5005
R24882 VSS.n2486 VSS.n2450 4.5005
R24883 VSS.n2489 VSS.n2450 4.5005
R24884 VSS.n2491 VSS.n2450 4.5005
R24885 VSS.n2492 VSS.n2450 4.5005
R24886 VSS.n2494 VSS.n2450 4.5005
R24887 VSS.n2497 VSS.n2450 4.5005
R24888 VSS.n2499 VSS.n2450 4.5005
R24889 VSS.n2500 VSS.n2450 4.5005
R24890 VSS.n2502 VSS.n2450 4.5005
R24891 VSS.n2505 VSS.n2450 4.5005
R24892 VSS.n2507 VSS.n2450 4.5005
R24893 VSS.n2508 VSS.n2450 4.5005
R24894 VSS.n2510 VSS.n2450 4.5005
R24895 VSS.n2513 VSS.n2450 4.5005
R24896 VSS.n2515 VSS.n2450 4.5005
R24897 VSS.n2516 VSS.n2450 4.5005
R24898 VSS.n2518 VSS.n2450 4.5005
R24899 VSS.n2521 VSS.n2450 4.5005
R24900 VSS.n2523 VSS.n2450 4.5005
R24901 VSS.n2524 VSS.n2450 4.5005
R24902 VSS.n2526 VSS.n2450 4.5005
R24903 VSS.n2529 VSS.n2450 4.5005
R24904 VSS.n2531 VSS.n2450 4.5005
R24905 VSS.n2532 VSS.n2450 4.5005
R24906 VSS.n2534 VSS.n2450 4.5005
R24907 VSS.n2537 VSS.n2450 4.5005
R24908 VSS.n2539 VSS.n2450 4.5005
R24909 VSS.n2540 VSS.n2450 4.5005
R24910 VSS.n2542 VSS.n2450 4.5005
R24911 VSS.n2545 VSS.n2450 4.5005
R24912 VSS.n2547 VSS.n2450 4.5005
R24913 VSS.n2548 VSS.n2450 4.5005
R24914 VSS.n2550 VSS.n2450 4.5005
R24915 VSS.n2553 VSS.n2450 4.5005
R24916 VSS.n2555 VSS.n2450 4.5005
R24917 VSS.n2556 VSS.n2450 4.5005
R24918 VSS.n2558 VSS.n2450 4.5005
R24919 VSS.n2561 VSS.n2450 4.5005
R24920 VSS.n2563 VSS.n2450 4.5005
R24921 VSS.n2564 VSS.n2450 4.5005
R24922 VSS.n2566 VSS.n2450 4.5005
R24923 VSS.n2569 VSS.n2450 4.5005
R24924 VSS.n2571 VSS.n2450 4.5005
R24925 VSS.n2572 VSS.n2450 4.5005
R24926 VSS.n2574 VSS.n2450 4.5005
R24927 VSS.n2577 VSS.n2450 4.5005
R24928 VSS.n2579 VSS.n2450 4.5005
R24929 VSS.n2580 VSS.n2450 4.5005
R24930 VSS.n2582 VSS.n2450 4.5005
R24931 VSS.n2585 VSS.n2450 4.5005
R24932 VSS.n2587 VSS.n2450 4.5005
R24933 VSS.n2588 VSS.n2450 4.5005
R24934 VSS.n2590 VSS.n2450 4.5005
R24935 VSS.n2593 VSS.n2450 4.5005
R24936 VSS.n2595 VSS.n2450 4.5005
R24937 VSS.n2596 VSS.n2450 4.5005
R24938 VSS.n2598 VSS.n2450 4.5005
R24939 VSS.n2601 VSS.n2450 4.5005
R24940 VSS.n2603 VSS.n2450 4.5005
R24941 VSS.n2604 VSS.n2450 4.5005
R24942 VSS.n2606 VSS.n2450 4.5005
R24943 VSS.n2609 VSS.n2450 4.5005
R24944 VSS.n2611 VSS.n2450 4.5005
R24945 VSS.n2612 VSS.n2450 4.5005
R24946 VSS.n2614 VSS.n2450 4.5005
R24947 VSS.n2617 VSS.n2450 4.5005
R24948 VSS.n2619 VSS.n2450 4.5005
R24949 VSS.n2620 VSS.n2450 4.5005
R24950 VSS.n2622 VSS.n2450 4.5005
R24951 VSS.n2625 VSS.n2450 4.5005
R24952 VSS.n2627 VSS.n2450 4.5005
R24953 VSS.n2628 VSS.n2450 4.5005
R24954 VSS.n2630 VSS.n2450 4.5005
R24955 VSS.n2633 VSS.n2450 4.5005
R24956 VSS.n2635 VSS.n2450 4.5005
R24957 VSS.n2636 VSS.n2450 4.5005
R24958 VSS.n2638 VSS.n2450 4.5005
R24959 VSS.n2640 VSS.n2450 4.5005
R24960 VSS.n2642 VSS.n2450 4.5005
R24961 VSS.n2643 VSS.n2450 4.5005
R24962 VSS.n2645 VSS.n2450 4.5005
R24963 VSS.n2648 VSS.n2450 4.5005
R24964 VSS.n2650 VSS.n2450 4.5005
R24965 VSS.n2651 VSS.n2450 4.5005
R24966 VSS.n2653 VSS.n2450 4.5005
R24967 VSS.n2656 VSS.n2450 4.5005
R24968 VSS.n2658 VSS.n2450 4.5005
R24969 VSS.n2659 VSS.n2450 4.5005
R24970 VSS.n2661 VSS.n2450 4.5005
R24971 VSS.n2664 VSS.n2450 4.5005
R24972 VSS.n2666 VSS.n2450 4.5005
R24973 VSS.n2667 VSS.n2450 4.5005
R24974 VSS.n2669 VSS.n2450 4.5005
R24975 VSS.n2672 VSS.n2450 4.5005
R24976 VSS.n2674 VSS.n2450 4.5005
R24977 VSS.n2675 VSS.n2450 4.5005
R24978 VSS.n2677 VSS.n2450 4.5005
R24979 VSS.n2680 VSS.n2450 4.5005
R24980 VSS.n2682 VSS.n2450 4.5005
R24981 VSS.n2683 VSS.n2450 4.5005
R24982 VSS.n2685 VSS.n2450 4.5005
R24983 VSS.n2688 VSS.n2450 4.5005
R24984 VSS.n2690 VSS.n2450 4.5005
R24985 VSS.n2691 VSS.n2450 4.5005
R24986 VSS.n2693 VSS.n2450 4.5005
R24987 VSS.n2696 VSS.n2450 4.5005
R24988 VSS.n2698 VSS.n2450 4.5005
R24989 VSS.n2699 VSS.n2450 4.5005
R24990 VSS.n2701 VSS.n2450 4.5005
R24991 VSS.n2704 VSS.n2450 4.5005
R24992 VSS.n2706 VSS.n2450 4.5005
R24993 VSS.n2707 VSS.n2450 4.5005
R24994 VSS.n2709 VSS.n2450 4.5005
R24995 VSS.n2712 VSS.n2450 4.5005
R24996 VSS.n2714 VSS.n2450 4.5005
R24997 VSS.n2715 VSS.n2450 4.5005
R24998 VSS.n2717 VSS.n2450 4.5005
R24999 VSS.n2720 VSS.n2450 4.5005
R25000 VSS.n2722 VSS.n2450 4.5005
R25001 VSS.n2723 VSS.n2450 4.5005
R25002 VSS.n2725 VSS.n2450 4.5005
R25003 VSS.n2793 VSS.n2450 4.5005
R25004 VSS.n2859 VSS.n2450 4.5005
R25005 VSS.n3051 VSS.n2381 4.5005
R25006 VSS.n2381 VSS.n2351 4.5005
R25007 VSS.n2483 VSS.n2381 4.5005
R25008 VSS.n2484 VSS.n2381 4.5005
R25009 VSS.n2486 VSS.n2381 4.5005
R25010 VSS.n2489 VSS.n2381 4.5005
R25011 VSS.n2491 VSS.n2381 4.5005
R25012 VSS.n2492 VSS.n2381 4.5005
R25013 VSS.n2494 VSS.n2381 4.5005
R25014 VSS.n2497 VSS.n2381 4.5005
R25015 VSS.n2499 VSS.n2381 4.5005
R25016 VSS.n2500 VSS.n2381 4.5005
R25017 VSS.n2502 VSS.n2381 4.5005
R25018 VSS.n2505 VSS.n2381 4.5005
R25019 VSS.n2507 VSS.n2381 4.5005
R25020 VSS.n2508 VSS.n2381 4.5005
R25021 VSS.n2510 VSS.n2381 4.5005
R25022 VSS.n2513 VSS.n2381 4.5005
R25023 VSS.n2515 VSS.n2381 4.5005
R25024 VSS.n2516 VSS.n2381 4.5005
R25025 VSS.n2518 VSS.n2381 4.5005
R25026 VSS.n2521 VSS.n2381 4.5005
R25027 VSS.n2523 VSS.n2381 4.5005
R25028 VSS.n2524 VSS.n2381 4.5005
R25029 VSS.n2526 VSS.n2381 4.5005
R25030 VSS.n2529 VSS.n2381 4.5005
R25031 VSS.n2531 VSS.n2381 4.5005
R25032 VSS.n2532 VSS.n2381 4.5005
R25033 VSS.n2534 VSS.n2381 4.5005
R25034 VSS.n2537 VSS.n2381 4.5005
R25035 VSS.n2539 VSS.n2381 4.5005
R25036 VSS.n2540 VSS.n2381 4.5005
R25037 VSS.n2542 VSS.n2381 4.5005
R25038 VSS.n2545 VSS.n2381 4.5005
R25039 VSS.n2547 VSS.n2381 4.5005
R25040 VSS.n2548 VSS.n2381 4.5005
R25041 VSS.n2550 VSS.n2381 4.5005
R25042 VSS.n2553 VSS.n2381 4.5005
R25043 VSS.n2555 VSS.n2381 4.5005
R25044 VSS.n2556 VSS.n2381 4.5005
R25045 VSS.n2558 VSS.n2381 4.5005
R25046 VSS.n2561 VSS.n2381 4.5005
R25047 VSS.n2563 VSS.n2381 4.5005
R25048 VSS.n2564 VSS.n2381 4.5005
R25049 VSS.n2566 VSS.n2381 4.5005
R25050 VSS.n2569 VSS.n2381 4.5005
R25051 VSS.n2571 VSS.n2381 4.5005
R25052 VSS.n2572 VSS.n2381 4.5005
R25053 VSS.n2574 VSS.n2381 4.5005
R25054 VSS.n2577 VSS.n2381 4.5005
R25055 VSS.n2579 VSS.n2381 4.5005
R25056 VSS.n2580 VSS.n2381 4.5005
R25057 VSS.n2582 VSS.n2381 4.5005
R25058 VSS.n2585 VSS.n2381 4.5005
R25059 VSS.n2587 VSS.n2381 4.5005
R25060 VSS.n2588 VSS.n2381 4.5005
R25061 VSS.n2590 VSS.n2381 4.5005
R25062 VSS.n2593 VSS.n2381 4.5005
R25063 VSS.n2595 VSS.n2381 4.5005
R25064 VSS.n2596 VSS.n2381 4.5005
R25065 VSS.n2598 VSS.n2381 4.5005
R25066 VSS.n2601 VSS.n2381 4.5005
R25067 VSS.n2603 VSS.n2381 4.5005
R25068 VSS.n2604 VSS.n2381 4.5005
R25069 VSS.n2606 VSS.n2381 4.5005
R25070 VSS.n2609 VSS.n2381 4.5005
R25071 VSS.n2611 VSS.n2381 4.5005
R25072 VSS.n2612 VSS.n2381 4.5005
R25073 VSS.n2614 VSS.n2381 4.5005
R25074 VSS.n2617 VSS.n2381 4.5005
R25075 VSS.n2619 VSS.n2381 4.5005
R25076 VSS.n2620 VSS.n2381 4.5005
R25077 VSS.n2622 VSS.n2381 4.5005
R25078 VSS.n2625 VSS.n2381 4.5005
R25079 VSS.n2627 VSS.n2381 4.5005
R25080 VSS.n2628 VSS.n2381 4.5005
R25081 VSS.n2630 VSS.n2381 4.5005
R25082 VSS.n2633 VSS.n2381 4.5005
R25083 VSS.n2635 VSS.n2381 4.5005
R25084 VSS.n2636 VSS.n2381 4.5005
R25085 VSS.n2638 VSS.n2381 4.5005
R25086 VSS.n2640 VSS.n2381 4.5005
R25087 VSS.n2642 VSS.n2381 4.5005
R25088 VSS.n2643 VSS.n2381 4.5005
R25089 VSS.n2645 VSS.n2381 4.5005
R25090 VSS.n2648 VSS.n2381 4.5005
R25091 VSS.n2650 VSS.n2381 4.5005
R25092 VSS.n2651 VSS.n2381 4.5005
R25093 VSS.n2653 VSS.n2381 4.5005
R25094 VSS.n2656 VSS.n2381 4.5005
R25095 VSS.n2658 VSS.n2381 4.5005
R25096 VSS.n2659 VSS.n2381 4.5005
R25097 VSS.n2661 VSS.n2381 4.5005
R25098 VSS.n2664 VSS.n2381 4.5005
R25099 VSS.n2666 VSS.n2381 4.5005
R25100 VSS.n2667 VSS.n2381 4.5005
R25101 VSS.n2669 VSS.n2381 4.5005
R25102 VSS.n2672 VSS.n2381 4.5005
R25103 VSS.n2674 VSS.n2381 4.5005
R25104 VSS.n2675 VSS.n2381 4.5005
R25105 VSS.n2677 VSS.n2381 4.5005
R25106 VSS.n2680 VSS.n2381 4.5005
R25107 VSS.n2682 VSS.n2381 4.5005
R25108 VSS.n2683 VSS.n2381 4.5005
R25109 VSS.n2685 VSS.n2381 4.5005
R25110 VSS.n2688 VSS.n2381 4.5005
R25111 VSS.n2690 VSS.n2381 4.5005
R25112 VSS.n2691 VSS.n2381 4.5005
R25113 VSS.n2693 VSS.n2381 4.5005
R25114 VSS.n2696 VSS.n2381 4.5005
R25115 VSS.n2698 VSS.n2381 4.5005
R25116 VSS.n2699 VSS.n2381 4.5005
R25117 VSS.n2701 VSS.n2381 4.5005
R25118 VSS.n2704 VSS.n2381 4.5005
R25119 VSS.n2706 VSS.n2381 4.5005
R25120 VSS.n2707 VSS.n2381 4.5005
R25121 VSS.n2709 VSS.n2381 4.5005
R25122 VSS.n2712 VSS.n2381 4.5005
R25123 VSS.n2714 VSS.n2381 4.5005
R25124 VSS.n2715 VSS.n2381 4.5005
R25125 VSS.n2717 VSS.n2381 4.5005
R25126 VSS.n2720 VSS.n2381 4.5005
R25127 VSS.n2722 VSS.n2381 4.5005
R25128 VSS.n2723 VSS.n2381 4.5005
R25129 VSS.n2725 VSS.n2381 4.5005
R25130 VSS.n2793 VSS.n2381 4.5005
R25131 VSS.n2859 VSS.n2381 4.5005
R25132 VSS.n3051 VSS.n2451 4.5005
R25133 VSS.n2451 VSS.n2351 4.5005
R25134 VSS.n2483 VSS.n2451 4.5005
R25135 VSS.n2484 VSS.n2451 4.5005
R25136 VSS.n2486 VSS.n2451 4.5005
R25137 VSS.n2489 VSS.n2451 4.5005
R25138 VSS.n2491 VSS.n2451 4.5005
R25139 VSS.n2492 VSS.n2451 4.5005
R25140 VSS.n2494 VSS.n2451 4.5005
R25141 VSS.n2497 VSS.n2451 4.5005
R25142 VSS.n2499 VSS.n2451 4.5005
R25143 VSS.n2500 VSS.n2451 4.5005
R25144 VSS.n2502 VSS.n2451 4.5005
R25145 VSS.n2505 VSS.n2451 4.5005
R25146 VSS.n2507 VSS.n2451 4.5005
R25147 VSS.n2508 VSS.n2451 4.5005
R25148 VSS.n2510 VSS.n2451 4.5005
R25149 VSS.n2513 VSS.n2451 4.5005
R25150 VSS.n2515 VSS.n2451 4.5005
R25151 VSS.n2516 VSS.n2451 4.5005
R25152 VSS.n2518 VSS.n2451 4.5005
R25153 VSS.n2521 VSS.n2451 4.5005
R25154 VSS.n2523 VSS.n2451 4.5005
R25155 VSS.n2524 VSS.n2451 4.5005
R25156 VSS.n2526 VSS.n2451 4.5005
R25157 VSS.n2529 VSS.n2451 4.5005
R25158 VSS.n2531 VSS.n2451 4.5005
R25159 VSS.n2532 VSS.n2451 4.5005
R25160 VSS.n2534 VSS.n2451 4.5005
R25161 VSS.n2537 VSS.n2451 4.5005
R25162 VSS.n2539 VSS.n2451 4.5005
R25163 VSS.n2540 VSS.n2451 4.5005
R25164 VSS.n2542 VSS.n2451 4.5005
R25165 VSS.n2545 VSS.n2451 4.5005
R25166 VSS.n2547 VSS.n2451 4.5005
R25167 VSS.n2548 VSS.n2451 4.5005
R25168 VSS.n2550 VSS.n2451 4.5005
R25169 VSS.n2553 VSS.n2451 4.5005
R25170 VSS.n2555 VSS.n2451 4.5005
R25171 VSS.n2556 VSS.n2451 4.5005
R25172 VSS.n2558 VSS.n2451 4.5005
R25173 VSS.n2561 VSS.n2451 4.5005
R25174 VSS.n2563 VSS.n2451 4.5005
R25175 VSS.n2564 VSS.n2451 4.5005
R25176 VSS.n2566 VSS.n2451 4.5005
R25177 VSS.n2569 VSS.n2451 4.5005
R25178 VSS.n2571 VSS.n2451 4.5005
R25179 VSS.n2572 VSS.n2451 4.5005
R25180 VSS.n2574 VSS.n2451 4.5005
R25181 VSS.n2577 VSS.n2451 4.5005
R25182 VSS.n2579 VSS.n2451 4.5005
R25183 VSS.n2580 VSS.n2451 4.5005
R25184 VSS.n2582 VSS.n2451 4.5005
R25185 VSS.n2585 VSS.n2451 4.5005
R25186 VSS.n2587 VSS.n2451 4.5005
R25187 VSS.n2588 VSS.n2451 4.5005
R25188 VSS.n2590 VSS.n2451 4.5005
R25189 VSS.n2593 VSS.n2451 4.5005
R25190 VSS.n2595 VSS.n2451 4.5005
R25191 VSS.n2596 VSS.n2451 4.5005
R25192 VSS.n2598 VSS.n2451 4.5005
R25193 VSS.n2601 VSS.n2451 4.5005
R25194 VSS.n2603 VSS.n2451 4.5005
R25195 VSS.n2604 VSS.n2451 4.5005
R25196 VSS.n2606 VSS.n2451 4.5005
R25197 VSS.n2609 VSS.n2451 4.5005
R25198 VSS.n2611 VSS.n2451 4.5005
R25199 VSS.n2612 VSS.n2451 4.5005
R25200 VSS.n2614 VSS.n2451 4.5005
R25201 VSS.n2617 VSS.n2451 4.5005
R25202 VSS.n2619 VSS.n2451 4.5005
R25203 VSS.n2620 VSS.n2451 4.5005
R25204 VSS.n2622 VSS.n2451 4.5005
R25205 VSS.n2625 VSS.n2451 4.5005
R25206 VSS.n2627 VSS.n2451 4.5005
R25207 VSS.n2628 VSS.n2451 4.5005
R25208 VSS.n2630 VSS.n2451 4.5005
R25209 VSS.n2633 VSS.n2451 4.5005
R25210 VSS.n2635 VSS.n2451 4.5005
R25211 VSS.n2636 VSS.n2451 4.5005
R25212 VSS.n2638 VSS.n2451 4.5005
R25213 VSS.n2640 VSS.n2451 4.5005
R25214 VSS.n2642 VSS.n2451 4.5005
R25215 VSS.n2643 VSS.n2451 4.5005
R25216 VSS.n2645 VSS.n2451 4.5005
R25217 VSS.n2648 VSS.n2451 4.5005
R25218 VSS.n2650 VSS.n2451 4.5005
R25219 VSS.n2651 VSS.n2451 4.5005
R25220 VSS.n2653 VSS.n2451 4.5005
R25221 VSS.n2656 VSS.n2451 4.5005
R25222 VSS.n2658 VSS.n2451 4.5005
R25223 VSS.n2659 VSS.n2451 4.5005
R25224 VSS.n2661 VSS.n2451 4.5005
R25225 VSS.n2664 VSS.n2451 4.5005
R25226 VSS.n2666 VSS.n2451 4.5005
R25227 VSS.n2667 VSS.n2451 4.5005
R25228 VSS.n2669 VSS.n2451 4.5005
R25229 VSS.n2672 VSS.n2451 4.5005
R25230 VSS.n2674 VSS.n2451 4.5005
R25231 VSS.n2675 VSS.n2451 4.5005
R25232 VSS.n2677 VSS.n2451 4.5005
R25233 VSS.n2680 VSS.n2451 4.5005
R25234 VSS.n2682 VSS.n2451 4.5005
R25235 VSS.n2683 VSS.n2451 4.5005
R25236 VSS.n2685 VSS.n2451 4.5005
R25237 VSS.n2688 VSS.n2451 4.5005
R25238 VSS.n2690 VSS.n2451 4.5005
R25239 VSS.n2691 VSS.n2451 4.5005
R25240 VSS.n2693 VSS.n2451 4.5005
R25241 VSS.n2696 VSS.n2451 4.5005
R25242 VSS.n2698 VSS.n2451 4.5005
R25243 VSS.n2699 VSS.n2451 4.5005
R25244 VSS.n2701 VSS.n2451 4.5005
R25245 VSS.n2704 VSS.n2451 4.5005
R25246 VSS.n2706 VSS.n2451 4.5005
R25247 VSS.n2707 VSS.n2451 4.5005
R25248 VSS.n2709 VSS.n2451 4.5005
R25249 VSS.n2712 VSS.n2451 4.5005
R25250 VSS.n2714 VSS.n2451 4.5005
R25251 VSS.n2715 VSS.n2451 4.5005
R25252 VSS.n2717 VSS.n2451 4.5005
R25253 VSS.n2720 VSS.n2451 4.5005
R25254 VSS.n2722 VSS.n2451 4.5005
R25255 VSS.n2723 VSS.n2451 4.5005
R25256 VSS.n2725 VSS.n2451 4.5005
R25257 VSS.n2793 VSS.n2451 4.5005
R25258 VSS.n2859 VSS.n2451 4.5005
R25259 VSS.n3051 VSS.n2380 4.5005
R25260 VSS.n2380 VSS.n2351 4.5005
R25261 VSS.n2483 VSS.n2380 4.5005
R25262 VSS.n2484 VSS.n2380 4.5005
R25263 VSS.n2486 VSS.n2380 4.5005
R25264 VSS.n2489 VSS.n2380 4.5005
R25265 VSS.n2491 VSS.n2380 4.5005
R25266 VSS.n2492 VSS.n2380 4.5005
R25267 VSS.n2494 VSS.n2380 4.5005
R25268 VSS.n2497 VSS.n2380 4.5005
R25269 VSS.n2499 VSS.n2380 4.5005
R25270 VSS.n2500 VSS.n2380 4.5005
R25271 VSS.n2502 VSS.n2380 4.5005
R25272 VSS.n2505 VSS.n2380 4.5005
R25273 VSS.n2507 VSS.n2380 4.5005
R25274 VSS.n2508 VSS.n2380 4.5005
R25275 VSS.n2510 VSS.n2380 4.5005
R25276 VSS.n2513 VSS.n2380 4.5005
R25277 VSS.n2515 VSS.n2380 4.5005
R25278 VSS.n2516 VSS.n2380 4.5005
R25279 VSS.n2518 VSS.n2380 4.5005
R25280 VSS.n2521 VSS.n2380 4.5005
R25281 VSS.n2523 VSS.n2380 4.5005
R25282 VSS.n2524 VSS.n2380 4.5005
R25283 VSS.n2526 VSS.n2380 4.5005
R25284 VSS.n2529 VSS.n2380 4.5005
R25285 VSS.n2531 VSS.n2380 4.5005
R25286 VSS.n2532 VSS.n2380 4.5005
R25287 VSS.n2534 VSS.n2380 4.5005
R25288 VSS.n2537 VSS.n2380 4.5005
R25289 VSS.n2539 VSS.n2380 4.5005
R25290 VSS.n2540 VSS.n2380 4.5005
R25291 VSS.n2542 VSS.n2380 4.5005
R25292 VSS.n2545 VSS.n2380 4.5005
R25293 VSS.n2547 VSS.n2380 4.5005
R25294 VSS.n2548 VSS.n2380 4.5005
R25295 VSS.n2550 VSS.n2380 4.5005
R25296 VSS.n2553 VSS.n2380 4.5005
R25297 VSS.n2555 VSS.n2380 4.5005
R25298 VSS.n2556 VSS.n2380 4.5005
R25299 VSS.n2558 VSS.n2380 4.5005
R25300 VSS.n2561 VSS.n2380 4.5005
R25301 VSS.n2563 VSS.n2380 4.5005
R25302 VSS.n2564 VSS.n2380 4.5005
R25303 VSS.n2566 VSS.n2380 4.5005
R25304 VSS.n2569 VSS.n2380 4.5005
R25305 VSS.n2571 VSS.n2380 4.5005
R25306 VSS.n2572 VSS.n2380 4.5005
R25307 VSS.n2574 VSS.n2380 4.5005
R25308 VSS.n2577 VSS.n2380 4.5005
R25309 VSS.n2579 VSS.n2380 4.5005
R25310 VSS.n2580 VSS.n2380 4.5005
R25311 VSS.n2582 VSS.n2380 4.5005
R25312 VSS.n2585 VSS.n2380 4.5005
R25313 VSS.n2587 VSS.n2380 4.5005
R25314 VSS.n2588 VSS.n2380 4.5005
R25315 VSS.n2590 VSS.n2380 4.5005
R25316 VSS.n2593 VSS.n2380 4.5005
R25317 VSS.n2595 VSS.n2380 4.5005
R25318 VSS.n2596 VSS.n2380 4.5005
R25319 VSS.n2598 VSS.n2380 4.5005
R25320 VSS.n2601 VSS.n2380 4.5005
R25321 VSS.n2603 VSS.n2380 4.5005
R25322 VSS.n2604 VSS.n2380 4.5005
R25323 VSS.n2606 VSS.n2380 4.5005
R25324 VSS.n2609 VSS.n2380 4.5005
R25325 VSS.n2611 VSS.n2380 4.5005
R25326 VSS.n2612 VSS.n2380 4.5005
R25327 VSS.n2614 VSS.n2380 4.5005
R25328 VSS.n2617 VSS.n2380 4.5005
R25329 VSS.n2619 VSS.n2380 4.5005
R25330 VSS.n2620 VSS.n2380 4.5005
R25331 VSS.n2622 VSS.n2380 4.5005
R25332 VSS.n2625 VSS.n2380 4.5005
R25333 VSS.n2627 VSS.n2380 4.5005
R25334 VSS.n2628 VSS.n2380 4.5005
R25335 VSS.n2630 VSS.n2380 4.5005
R25336 VSS.n2633 VSS.n2380 4.5005
R25337 VSS.n2635 VSS.n2380 4.5005
R25338 VSS.n2636 VSS.n2380 4.5005
R25339 VSS.n2638 VSS.n2380 4.5005
R25340 VSS.n2640 VSS.n2380 4.5005
R25341 VSS.n2642 VSS.n2380 4.5005
R25342 VSS.n2643 VSS.n2380 4.5005
R25343 VSS.n2645 VSS.n2380 4.5005
R25344 VSS.n2648 VSS.n2380 4.5005
R25345 VSS.n2650 VSS.n2380 4.5005
R25346 VSS.n2651 VSS.n2380 4.5005
R25347 VSS.n2653 VSS.n2380 4.5005
R25348 VSS.n2656 VSS.n2380 4.5005
R25349 VSS.n2658 VSS.n2380 4.5005
R25350 VSS.n2659 VSS.n2380 4.5005
R25351 VSS.n2661 VSS.n2380 4.5005
R25352 VSS.n2664 VSS.n2380 4.5005
R25353 VSS.n2666 VSS.n2380 4.5005
R25354 VSS.n2667 VSS.n2380 4.5005
R25355 VSS.n2669 VSS.n2380 4.5005
R25356 VSS.n2672 VSS.n2380 4.5005
R25357 VSS.n2674 VSS.n2380 4.5005
R25358 VSS.n2675 VSS.n2380 4.5005
R25359 VSS.n2677 VSS.n2380 4.5005
R25360 VSS.n2680 VSS.n2380 4.5005
R25361 VSS.n2682 VSS.n2380 4.5005
R25362 VSS.n2683 VSS.n2380 4.5005
R25363 VSS.n2685 VSS.n2380 4.5005
R25364 VSS.n2688 VSS.n2380 4.5005
R25365 VSS.n2690 VSS.n2380 4.5005
R25366 VSS.n2691 VSS.n2380 4.5005
R25367 VSS.n2693 VSS.n2380 4.5005
R25368 VSS.n2696 VSS.n2380 4.5005
R25369 VSS.n2698 VSS.n2380 4.5005
R25370 VSS.n2699 VSS.n2380 4.5005
R25371 VSS.n2701 VSS.n2380 4.5005
R25372 VSS.n2704 VSS.n2380 4.5005
R25373 VSS.n2706 VSS.n2380 4.5005
R25374 VSS.n2707 VSS.n2380 4.5005
R25375 VSS.n2709 VSS.n2380 4.5005
R25376 VSS.n2712 VSS.n2380 4.5005
R25377 VSS.n2714 VSS.n2380 4.5005
R25378 VSS.n2715 VSS.n2380 4.5005
R25379 VSS.n2717 VSS.n2380 4.5005
R25380 VSS.n2720 VSS.n2380 4.5005
R25381 VSS.n2722 VSS.n2380 4.5005
R25382 VSS.n2723 VSS.n2380 4.5005
R25383 VSS.n2725 VSS.n2380 4.5005
R25384 VSS.n2793 VSS.n2380 4.5005
R25385 VSS.n2859 VSS.n2380 4.5005
R25386 VSS.n3051 VSS.n2452 4.5005
R25387 VSS.n2452 VSS.n2351 4.5005
R25388 VSS.n2483 VSS.n2452 4.5005
R25389 VSS.n2484 VSS.n2452 4.5005
R25390 VSS.n2486 VSS.n2452 4.5005
R25391 VSS.n2489 VSS.n2452 4.5005
R25392 VSS.n2491 VSS.n2452 4.5005
R25393 VSS.n2492 VSS.n2452 4.5005
R25394 VSS.n2494 VSS.n2452 4.5005
R25395 VSS.n2497 VSS.n2452 4.5005
R25396 VSS.n2499 VSS.n2452 4.5005
R25397 VSS.n2500 VSS.n2452 4.5005
R25398 VSS.n2502 VSS.n2452 4.5005
R25399 VSS.n2505 VSS.n2452 4.5005
R25400 VSS.n2507 VSS.n2452 4.5005
R25401 VSS.n2508 VSS.n2452 4.5005
R25402 VSS.n2510 VSS.n2452 4.5005
R25403 VSS.n2513 VSS.n2452 4.5005
R25404 VSS.n2515 VSS.n2452 4.5005
R25405 VSS.n2516 VSS.n2452 4.5005
R25406 VSS.n2518 VSS.n2452 4.5005
R25407 VSS.n2521 VSS.n2452 4.5005
R25408 VSS.n2523 VSS.n2452 4.5005
R25409 VSS.n2524 VSS.n2452 4.5005
R25410 VSS.n2526 VSS.n2452 4.5005
R25411 VSS.n2529 VSS.n2452 4.5005
R25412 VSS.n2531 VSS.n2452 4.5005
R25413 VSS.n2532 VSS.n2452 4.5005
R25414 VSS.n2534 VSS.n2452 4.5005
R25415 VSS.n2537 VSS.n2452 4.5005
R25416 VSS.n2539 VSS.n2452 4.5005
R25417 VSS.n2540 VSS.n2452 4.5005
R25418 VSS.n2542 VSS.n2452 4.5005
R25419 VSS.n2545 VSS.n2452 4.5005
R25420 VSS.n2547 VSS.n2452 4.5005
R25421 VSS.n2548 VSS.n2452 4.5005
R25422 VSS.n2550 VSS.n2452 4.5005
R25423 VSS.n2553 VSS.n2452 4.5005
R25424 VSS.n2555 VSS.n2452 4.5005
R25425 VSS.n2556 VSS.n2452 4.5005
R25426 VSS.n2558 VSS.n2452 4.5005
R25427 VSS.n2561 VSS.n2452 4.5005
R25428 VSS.n2563 VSS.n2452 4.5005
R25429 VSS.n2564 VSS.n2452 4.5005
R25430 VSS.n2566 VSS.n2452 4.5005
R25431 VSS.n2569 VSS.n2452 4.5005
R25432 VSS.n2571 VSS.n2452 4.5005
R25433 VSS.n2572 VSS.n2452 4.5005
R25434 VSS.n2574 VSS.n2452 4.5005
R25435 VSS.n2577 VSS.n2452 4.5005
R25436 VSS.n2579 VSS.n2452 4.5005
R25437 VSS.n2580 VSS.n2452 4.5005
R25438 VSS.n2582 VSS.n2452 4.5005
R25439 VSS.n2585 VSS.n2452 4.5005
R25440 VSS.n2587 VSS.n2452 4.5005
R25441 VSS.n2588 VSS.n2452 4.5005
R25442 VSS.n2590 VSS.n2452 4.5005
R25443 VSS.n2593 VSS.n2452 4.5005
R25444 VSS.n2595 VSS.n2452 4.5005
R25445 VSS.n2596 VSS.n2452 4.5005
R25446 VSS.n2598 VSS.n2452 4.5005
R25447 VSS.n2601 VSS.n2452 4.5005
R25448 VSS.n2603 VSS.n2452 4.5005
R25449 VSS.n2604 VSS.n2452 4.5005
R25450 VSS.n2606 VSS.n2452 4.5005
R25451 VSS.n2609 VSS.n2452 4.5005
R25452 VSS.n2611 VSS.n2452 4.5005
R25453 VSS.n2612 VSS.n2452 4.5005
R25454 VSS.n2614 VSS.n2452 4.5005
R25455 VSS.n2617 VSS.n2452 4.5005
R25456 VSS.n2619 VSS.n2452 4.5005
R25457 VSS.n2620 VSS.n2452 4.5005
R25458 VSS.n2622 VSS.n2452 4.5005
R25459 VSS.n2625 VSS.n2452 4.5005
R25460 VSS.n2627 VSS.n2452 4.5005
R25461 VSS.n2628 VSS.n2452 4.5005
R25462 VSS.n2630 VSS.n2452 4.5005
R25463 VSS.n2633 VSS.n2452 4.5005
R25464 VSS.n2635 VSS.n2452 4.5005
R25465 VSS.n2636 VSS.n2452 4.5005
R25466 VSS.n2638 VSS.n2452 4.5005
R25467 VSS.n2640 VSS.n2452 4.5005
R25468 VSS.n2642 VSS.n2452 4.5005
R25469 VSS.n2643 VSS.n2452 4.5005
R25470 VSS.n2645 VSS.n2452 4.5005
R25471 VSS.n2648 VSS.n2452 4.5005
R25472 VSS.n2650 VSS.n2452 4.5005
R25473 VSS.n2651 VSS.n2452 4.5005
R25474 VSS.n2653 VSS.n2452 4.5005
R25475 VSS.n2656 VSS.n2452 4.5005
R25476 VSS.n2658 VSS.n2452 4.5005
R25477 VSS.n2659 VSS.n2452 4.5005
R25478 VSS.n2661 VSS.n2452 4.5005
R25479 VSS.n2664 VSS.n2452 4.5005
R25480 VSS.n2666 VSS.n2452 4.5005
R25481 VSS.n2667 VSS.n2452 4.5005
R25482 VSS.n2669 VSS.n2452 4.5005
R25483 VSS.n2672 VSS.n2452 4.5005
R25484 VSS.n2674 VSS.n2452 4.5005
R25485 VSS.n2675 VSS.n2452 4.5005
R25486 VSS.n2677 VSS.n2452 4.5005
R25487 VSS.n2680 VSS.n2452 4.5005
R25488 VSS.n2682 VSS.n2452 4.5005
R25489 VSS.n2683 VSS.n2452 4.5005
R25490 VSS.n2685 VSS.n2452 4.5005
R25491 VSS.n2688 VSS.n2452 4.5005
R25492 VSS.n2690 VSS.n2452 4.5005
R25493 VSS.n2691 VSS.n2452 4.5005
R25494 VSS.n2693 VSS.n2452 4.5005
R25495 VSS.n2696 VSS.n2452 4.5005
R25496 VSS.n2698 VSS.n2452 4.5005
R25497 VSS.n2699 VSS.n2452 4.5005
R25498 VSS.n2701 VSS.n2452 4.5005
R25499 VSS.n2704 VSS.n2452 4.5005
R25500 VSS.n2706 VSS.n2452 4.5005
R25501 VSS.n2707 VSS.n2452 4.5005
R25502 VSS.n2709 VSS.n2452 4.5005
R25503 VSS.n2712 VSS.n2452 4.5005
R25504 VSS.n2714 VSS.n2452 4.5005
R25505 VSS.n2715 VSS.n2452 4.5005
R25506 VSS.n2717 VSS.n2452 4.5005
R25507 VSS.n2720 VSS.n2452 4.5005
R25508 VSS.n2722 VSS.n2452 4.5005
R25509 VSS.n2723 VSS.n2452 4.5005
R25510 VSS.n2725 VSS.n2452 4.5005
R25511 VSS.n2793 VSS.n2452 4.5005
R25512 VSS.n2859 VSS.n2452 4.5005
R25513 VSS.n3051 VSS.n2379 4.5005
R25514 VSS.n2379 VSS.n2351 4.5005
R25515 VSS.n2483 VSS.n2379 4.5005
R25516 VSS.n2484 VSS.n2379 4.5005
R25517 VSS.n2486 VSS.n2379 4.5005
R25518 VSS.n2489 VSS.n2379 4.5005
R25519 VSS.n2491 VSS.n2379 4.5005
R25520 VSS.n2492 VSS.n2379 4.5005
R25521 VSS.n2494 VSS.n2379 4.5005
R25522 VSS.n2497 VSS.n2379 4.5005
R25523 VSS.n2499 VSS.n2379 4.5005
R25524 VSS.n2500 VSS.n2379 4.5005
R25525 VSS.n2502 VSS.n2379 4.5005
R25526 VSS.n2505 VSS.n2379 4.5005
R25527 VSS.n2507 VSS.n2379 4.5005
R25528 VSS.n2508 VSS.n2379 4.5005
R25529 VSS.n2510 VSS.n2379 4.5005
R25530 VSS.n2513 VSS.n2379 4.5005
R25531 VSS.n2515 VSS.n2379 4.5005
R25532 VSS.n2516 VSS.n2379 4.5005
R25533 VSS.n2518 VSS.n2379 4.5005
R25534 VSS.n2521 VSS.n2379 4.5005
R25535 VSS.n2523 VSS.n2379 4.5005
R25536 VSS.n2524 VSS.n2379 4.5005
R25537 VSS.n2526 VSS.n2379 4.5005
R25538 VSS.n2529 VSS.n2379 4.5005
R25539 VSS.n2531 VSS.n2379 4.5005
R25540 VSS.n2532 VSS.n2379 4.5005
R25541 VSS.n2534 VSS.n2379 4.5005
R25542 VSS.n2537 VSS.n2379 4.5005
R25543 VSS.n2539 VSS.n2379 4.5005
R25544 VSS.n2540 VSS.n2379 4.5005
R25545 VSS.n2542 VSS.n2379 4.5005
R25546 VSS.n2545 VSS.n2379 4.5005
R25547 VSS.n2547 VSS.n2379 4.5005
R25548 VSS.n2548 VSS.n2379 4.5005
R25549 VSS.n2550 VSS.n2379 4.5005
R25550 VSS.n2553 VSS.n2379 4.5005
R25551 VSS.n2555 VSS.n2379 4.5005
R25552 VSS.n2556 VSS.n2379 4.5005
R25553 VSS.n2558 VSS.n2379 4.5005
R25554 VSS.n2561 VSS.n2379 4.5005
R25555 VSS.n2563 VSS.n2379 4.5005
R25556 VSS.n2564 VSS.n2379 4.5005
R25557 VSS.n2566 VSS.n2379 4.5005
R25558 VSS.n2569 VSS.n2379 4.5005
R25559 VSS.n2571 VSS.n2379 4.5005
R25560 VSS.n2572 VSS.n2379 4.5005
R25561 VSS.n2574 VSS.n2379 4.5005
R25562 VSS.n2577 VSS.n2379 4.5005
R25563 VSS.n2579 VSS.n2379 4.5005
R25564 VSS.n2580 VSS.n2379 4.5005
R25565 VSS.n2582 VSS.n2379 4.5005
R25566 VSS.n2585 VSS.n2379 4.5005
R25567 VSS.n2587 VSS.n2379 4.5005
R25568 VSS.n2588 VSS.n2379 4.5005
R25569 VSS.n2590 VSS.n2379 4.5005
R25570 VSS.n2593 VSS.n2379 4.5005
R25571 VSS.n2595 VSS.n2379 4.5005
R25572 VSS.n2596 VSS.n2379 4.5005
R25573 VSS.n2598 VSS.n2379 4.5005
R25574 VSS.n2601 VSS.n2379 4.5005
R25575 VSS.n2603 VSS.n2379 4.5005
R25576 VSS.n2604 VSS.n2379 4.5005
R25577 VSS.n2606 VSS.n2379 4.5005
R25578 VSS.n2609 VSS.n2379 4.5005
R25579 VSS.n2611 VSS.n2379 4.5005
R25580 VSS.n2612 VSS.n2379 4.5005
R25581 VSS.n2614 VSS.n2379 4.5005
R25582 VSS.n2617 VSS.n2379 4.5005
R25583 VSS.n2619 VSS.n2379 4.5005
R25584 VSS.n2620 VSS.n2379 4.5005
R25585 VSS.n2622 VSS.n2379 4.5005
R25586 VSS.n2625 VSS.n2379 4.5005
R25587 VSS.n2627 VSS.n2379 4.5005
R25588 VSS.n2628 VSS.n2379 4.5005
R25589 VSS.n2630 VSS.n2379 4.5005
R25590 VSS.n2633 VSS.n2379 4.5005
R25591 VSS.n2635 VSS.n2379 4.5005
R25592 VSS.n2636 VSS.n2379 4.5005
R25593 VSS.n2638 VSS.n2379 4.5005
R25594 VSS.n2640 VSS.n2379 4.5005
R25595 VSS.n2642 VSS.n2379 4.5005
R25596 VSS.n2643 VSS.n2379 4.5005
R25597 VSS.n2645 VSS.n2379 4.5005
R25598 VSS.n2648 VSS.n2379 4.5005
R25599 VSS.n2650 VSS.n2379 4.5005
R25600 VSS.n2651 VSS.n2379 4.5005
R25601 VSS.n2653 VSS.n2379 4.5005
R25602 VSS.n2656 VSS.n2379 4.5005
R25603 VSS.n2658 VSS.n2379 4.5005
R25604 VSS.n2659 VSS.n2379 4.5005
R25605 VSS.n2661 VSS.n2379 4.5005
R25606 VSS.n2664 VSS.n2379 4.5005
R25607 VSS.n2666 VSS.n2379 4.5005
R25608 VSS.n2667 VSS.n2379 4.5005
R25609 VSS.n2669 VSS.n2379 4.5005
R25610 VSS.n2672 VSS.n2379 4.5005
R25611 VSS.n2674 VSS.n2379 4.5005
R25612 VSS.n2675 VSS.n2379 4.5005
R25613 VSS.n2677 VSS.n2379 4.5005
R25614 VSS.n2680 VSS.n2379 4.5005
R25615 VSS.n2682 VSS.n2379 4.5005
R25616 VSS.n2683 VSS.n2379 4.5005
R25617 VSS.n2685 VSS.n2379 4.5005
R25618 VSS.n2688 VSS.n2379 4.5005
R25619 VSS.n2690 VSS.n2379 4.5005
R25620 VSS.n2691 VSS.n2379 4.5005
R25621 VSS.n2693 VSS.n2379 4.5005
R25622 VSS.n2696 VSS.n2379 4.5005
R25623 VSS.n2698 VSS.n2379 4.5005
R25624 VSS.n2699 VSS.n2379 4.5005
R25625 VSS.n2701 VSS.n2379 4.5005
R25626 VSS.n2704 VSS.n2379 4.5005
R25627 VSS.n2706 VSS.n2379 4.5005
R25628 VSS.n2707 VSS.n2379 4.5005
R25629 VSS.n2709 VSS.n2379 4.5005
R25630 VSS.n2712 VSS.n2379 4.5005
R25631 VSS.n2714 VSS.n2379 4.5005
R25632 VSS.n2715 VSS.n2379 4.5005
R25633 VSS.n2717 VSS.n2379 4.5005
R25634 VSS.n2720 VSS.n2379 4.5005
R25635 VSS.n2722 VSS.n2379 4.5005
R25636 VSS.n2723 VSS.n2379 4.5005
R25637 VSS.n2725 VSS.n2379 4.5005
R25638 VSS.n2793 VSS.n2379 4.5005
R25639 VSS.n2859 VSS.n2379 4.5005
R25640 VSS.n3051 VSS.n2453 4.5005
R25641 VSS.n2453 VSS.n2351 4.5005
R25642 VSS.n2483 VSS.n2453 4.5005
R25643 VSS.n2484 VSS.n2453 4.5005
R25644 VSS.n2486 VSS.n2453 4.5005
R25645 VSS.n2489 VSS.n2453 4.5005
R25646 VSS.n2491 VSS.n2453 4.5005
R25647 VSS.n2492 VSS.n2453 4.5005
R25648 VSS.n2494 VSS.n2453 4.5005
R25649 VSS.n2497 VSS.n2453 4.5005
R25650 VSS.n2499 VSS.n2453 4.5005
R25651 VSS.n2500 VSS.n2453 4.5005
R25652 VSS.n2502 VSS.n2453 4.5005
R25653 VSS.n2505 VSS.n2453 4.5005
R25654 VSS.n2507 VSS.n2453 4.5005
R25655 VSS.n2508 VSS.n2453 4.5005
R25656 VSS.n2510 VSS.n2453 4.5005
R25657 VSS.n2513 VSS.n2453 4.5005
R25658 VSS.n2515 VSS.n2453 4.5005
R25659 VSS.n2516 VSS.n2453 4.5005
R25660 VSS.n2518 VSS.n2453 4.5005
R25661 VSS.n2521 VSS.n2453 4.5005
R25662 VSS.n2523 VSS.n2453 4.5005
R25663 VSS.n2524 VSS.n2453 4.5005
R25664 VSS.n2526 VSS.n2453 4.5005
R25665 VSS.n2529 VSS.n2453 4.5005
R25666 VSS.n2531 VSS.n2453 4.5005
R25667 VSS.n2532 VSS.n2453 4.5005
R25668 VSS.n2534 VSS.n2453 4.5005
R25669 VSS.n2537 VSS.n2453 4.5005
R25670 VSS.n2539 VSS.n2453 4.5005
R25671 VSS.n2540 VSS.n2453 4.5005
R25672 VSS.n2542 VSS.n2453 4.5005
R25673 VSS.n2545 VSS.n2453 4.5005
R25674 VSS.n2547 VSS.n2453 4.5005
R25675 VSS.n2548 VSS.n2453 4.5005
R25676 VSS.n2550 VSS.n2453 4.5005
R25677 VSS.n2553 VSS.n2453 4.5005
R25678 VSS.n2555 VSS.n2453 4.5005
R25679 VSS.n2556 VSS.n2453 4.5005
R25680 VSS.n2558 VSS.n2453 4.5005
R25681 VSS.n2561 VSS.n2453 4.5005
R25682 VSS.n2563 VSS.n2453 4.5005
R25683 VSS.n2564 VSS.n2453 4.5005
R25684 VSS.n2566 VSS.n2453 4.5005
R25685 VSS.n2569 VSS.n2453 4.5005
R25686 VSS.n2571 VSS.n2453 4.5005
R25687 VSS.n2572 VSS.n2453 4.5005
R25688 VSS.n2574 VSS.n2453 4.5005
R25689 VSS.n2577 VSS.n2453 4.5005
R25690 VSS.n2579 VSS.n2453 4.5005
R25691 VSS.n2580 VSS.n2453 4.5005
R25692 VSS.n2582 VSS.n2453 4.5005
R25693 VSS.n2585 VSS.n2453 4.5005
R25694 VSS.n2587 VSS.n2453 4.5005
R25695 VSS.n2588 VSS.n2453 4.5005
R25696 VSS.n2590 VSS.n2453 4.5005
R25697 VSS.n2593 VSS.n2453 4.5005
R25698 VSS.n2595 VSS.n2453 4.5005
R25699 VSS.n2596 VSS.n2453 4.5005
R25700 VSS.n2598 VSS.n2453 4.5005
R25701 VSS.n2601 VSS.n2453 4.5005
R25702 VSS.n2603 VSS.n2453 4.5005
R25703 VSS.n2604 VSS.n2453 4.5005
R25704 VSS.n2606 VSS.n2453 4.5005
R25705 VSS.n2609 VSS.n2453 4.5005
R25706 VSS.n2611 VSS.n2453 4.5005
R25707 VSS.n2612 VSS.n2453 4.5005
R25708 VSS.n2614 VSS.n2453 4.5005
R25709 VSS.n2617 VSS.n2453 4.5005
R25710 VSS.n2619 VSS.n2453 4.5005
R25711 VSS.n2620 VSS.n2453 4.5005
R25712 VSS.n2622 VSS.n2453 4.5005
R25713 VSS.n2625 VSS.n2453 4.5005
R25714 VSS.n2627 VSS.n2453 4.5005
R25715 VSS.n2628 VSS.n2453 4.5005
R25716 VSS.n2630 VSS.n2453 4.5005
R25717 VSS.n2633 VSS.n2453 4.5005
R25718 VSS.n2635 VSS.n2453 4.5005
R25719 VSS.n2636 VSS.n2453 4.5005
R25720 VSS.n2638 VSS.n2453 4.5005
R25721 VSS.n2640 VSS.n2453 4.5005
R25722 VSS.n2642 VSS.n2453 4.5005
R25723 VSS.n2643 VSS.n2453 4.5005
R25724 VSS.n2645 VSS.n2453 4.5005
R25725 VSS.n2648 VSS.n2453 4.5005
R25726 VSS.n2650 VSS.n2453 4.5005
R25727 VSS.n2651 VSS.n2453 4.5005
R25728 VSS.n2653 VSS.n2453 4.5005
R25729 VSS.n2656 VSS.n2453 4.5005
R25730 VSS.n2658 VSS.n2453 4.5005
R25731 VSS.n2659 VSS.n2453 4.5005
R25732 VSS.n2661 VSS.n2453 4.5005
R25733 VSS.n2664 VSS.n2453 4.5005
R25734 VSS.n2666 VSS.n2453 4.5005
R25735 VSS.n2667 VSS.n2453 4.5005
R25736 VSS.n2669 VSS.n2453 4.5005
R25737 VSS.n2672 VSS.n2453 4.5005
R25738 VSS.n2674 VSS.n2453 4.5005
R25739 VSS.n2675 VSS.n2453 4.5005
R25740 VSS.n2677 VSS.n2453 4.5005
R25741 VSS.n2680 VSS.n2453 4.5005
R25742 VSS.n2682 VSS.n2453 4.5005
R25743 VSS.n2683 VSS.n2453 4.5005
R25744 VSS.n2685 VSS.n2453 4.5005
R25745 VSS.n2688 VSS.n2453 4.5005
R25746 VSS.n2690 VSS.n2453 4.5005
R25747 VSS.n2691 VSS.n2453 4.5005
R25748 VSS.n2693 VSS.n2453 4.5005
R25749 VSS.n2696 VSS.n2453 4.5005
R25750 VSS.n2698 VSS.n2453 4.5005
R25751 VSS.n2699 VSS.n2453 4.5005
R25752 VSS.n2701 VSS.n2453 4.5005
R25753 VSS.n2704 VSS.n2453 4.5005
R25754 VSS.n2706 VSS.n2453 4.5005
R25755 VSS.n2707 VSS.n2453 4.5005
R25756 VSS.n2709 VSS.n2453 4.5005
R25757 VSS.n2712 VSS.n2453 4.5005
R25758 VSS.n2714 VSS.n2453 4.5005
R25759 VSS.n2715 VSS.n2453 4.5005
R25760 VSS.n2717 VSS.n2453 4.5005
R25761 VSS.n2720 VSS.n2453 4.5005
R25762 VSS.n2722 VSS.n2453 4.5005
R25763 VSS.n2723 VSS.n2453 4.5005
R25764 VSS.n2725 VSS.n2453 4.5005
R25765 VSS.n2793 VSS.n2453 4.5005
R25766 VSS.n2859 VSS.n2453 4.5005
R25767 VSS.n3051 VSS.n2378 4.5005
R25768 VSS.n2378 VSS.n2351 4.5005
R25769 VSS.n2483 VSS.n2378 4.5005
R25770 VSS.n2484 VSS.n2378 4.5005
R25771 VSS.n2486 VSS.n2378 4.5005
R25772 VSS.n2489 VSS.n2378 4.5005
R25773 VSS.n2491 VSS.n2378 4.5005
R25774 VSS.n2492 VSS.n2378 4.5005
R25775 VSS.n2494 VSS.n2378 4.5005
R25776 VSS.n2497 VSS.n2378 4.5005
R25777 VSS.n2499 VSS.n2378 4.5005
R25778 VSS.n2500 VSS.n2378 4.5005
R25779 VSS.n2502 VSS.n2378 4.5005
R25780 VSS.n2505 VSS.n2378 4.5005
R25781 VSS.n2507 VSS.n2378 4.5005
R25782 VSS.n2508 VSS.n2378 4.5005
R25783 VSS.n2510 VSS.n2378 4.5005
R25784 VSS.n2513 VSS.n2378 4.5005
R25785 VSS.n2515 VSS.n2378 4.5005
R25786 VSS.n2516 VSS.n2378 4.5005
R25787 VSS.n2518 VSS.n2378 4.5005
R25788 VSS.n2521 VSS.n2378 4.5005
R25789 VSS.n2523 VSS.n2378 4.5005
R25790 VSS.n2524 VSS.n2378 4.5005
R25791 VSS.n2526 VSS.n2378 4.5005
R25792 VSS.n2529 VSS.n2378 4.5005
R25793 VSS.n2531 VSS.n2378 4.5005
R25794 VSS.n2532 VSS.n2378 4.5005
R25795 VSS.n2534 VSS.n2378 4.5005
R25796 VSS.n2537 VSS.n2378 4.5005
R25797 VSS.n2539 VSS.n2378 4.5005
R25798 VSS.n2540 VSS.n2378 4.5005
R25799 VSS.n2542 VSS.n2378 4.5005
R25800 VSS.n2545 VSS.n2378 4.5005
R25801 VSS.n2547 VSS.n2378 4.5005
R25802 VSS.n2548 VSS.n2378 4.5005
R25803 VSS.n2550 VSS.n2378 4.5005
R25804 VSS.n2553 VSS.n2378 4.5005
R25805 VSS.n2555 VSS.n2378 4.5005
R25806 VSS.n2556 VSS.n2378 4.5005
R25807 VSS.n2558 VSS.n2378 4.5005
R25808 VSS.n2561 VSS.n2378 4.5005
R25809 VSS.n2563 VSS.n2378 4.5005
R25810 VSS.n2564 VSS.n2378 4.5005
R25811 VSS.n2566 VSS.n2378 4.5005
R25812 VSS.n2569 VSS.n2378 4.5005
R25813 VSS.n2571 VSS.n2378 4.5005
R25814 VSS.n2572 VSS.n2378 4.5005
R25815 VSS.n2574 VSS.n2378 4.5005
R25816 VSS.n2577 VSS.n2378 4.5005
R25817 VSS.n2579 VSS.n2378 4.5005
R25818 VSS.n2580 VSS.n2378 4.5005
R25819 VSS.n2582 VSS.n2378 4.5005
R25820 VSS.n2585 VSS.n2378 4.5005
R25821 VSS.n2587 VSS.n2378 4.5005
R25822 VSS.n2588 VSS.n2378 4.5005
R25823 VSS.n2590 VSS.n2378 4.5005
R25824 VSS.n2593 VSS.n2378 4.5005
R25825 VSS.n2595 VSS.n2378 4.5005
R25826 VSS.n2596 VSS.n2378 4.5005
R25827 VSS.n2598 VSS.n2378 4.5005
R25828 VSS.n2601 VSS.n2378 4.5005
R25829 VSS.n2603 VSS.n2378 4.5005
R25830 VSS.n2604 VSS.n2378 4.5005
R25831 VSS.n2606 VSS.n2378 4.5005
R25832 VSS.n2609 VSS.n2378 4.5005
R25833 VSS.n2611 VSS.n2378 4.5005
R25834 VSS.n2612 VSS.n2378 4.5005
R25835 VSS.n2614 VSS.n2378 4.5005
R25836 VSS.n2617 VSS.n2378 4.5005
R25837 VSS.n2619 VSS.n2378 4.5005
R25838 VSS.n2620 VSS.n2378 4.5005
R25839 VSS.n2622 VSS.n2378 4.5005
R25840 VSS.n2625 VSS.n2378 4.5005
R25841 VSS.n2627 VSS.n2378 4.5005
R25842 VSS.n2628 VSS.n2378 4.5005
R25843 VSS.n2630 VSS.n2378 4.5005
R25844 VSS.n2633 VSS.n2378 4.5005
R25845 VSS.n2635 VSS.n2378 4.5005
R25846 VSS.n2636 VSS.n2378 4.5005
R25847 VSS.n2638 VSS.n2378 4.5005
R25848 VSS.n2640 VSS.n2378 4.5005
R25849 VSS.n2642 VSS.n2378 4.5005
R25850 VSS.n2643 VSS.n2378 4.5005
R25851 VSS.n2645 VSS.n2378 4.5005
R25852 VSS.n2648 VSS.n2378 4.5005
R25853 VSS.n2650 VSS.n2378 4.5005
R25854 VSS.n2651 VSS.n2378 4.5005
R25855 VSS.n2653 VSS.n2378 4.5005
R25856 VSS.n2656 VSS.n2378 4.5005
R25857 VSS.n2658 VSS.n2378 4.5005
R25858 VSS.n2659 VSS.n2378 4.5005
R25859 VSS.n2661 VSS.n2378 4.5005
R25860 VSS.n2664 VSS.n2378 4.5005
R25861 VSS.n2666 VSS.n2378 4.5005
R25862 VSS.n2667 VSS.n2378 4.5005
R25863 VSS.n2669 VSS.n2378 4.5005
R25864 VSS.n2672 VSS.n2378 4.5005
R25865 VSS.n2674 VSS.n2378 4.5005
R25866 VSS.n2675 VSS.n2378 4.5005
R25867 VSS.n2677 VSS.n2378 4.5005
R25868 VSS.n2680 VSS.n2378 4.5005
R25869 VSS.n2682 VSS.n2378 4.5005
R25870 VSS.n2683 VSS.n2378 4.5005
R25871 VSS.n2685 VSS.n2378 4.5005
R25872 VSS.n2688 VSS.n2378 4.5005
R25873 VSS.n2690 VSS.n2378 4.5005
R25874 VSS.n2691 VSS.n2378 4.5005
R25875 VSS.n2693 VSS.n2378 4.5005
R25876 VSS.n2696 VSS.n2378 4.5005
R25877 VSS.n2698 VSS.n2378 4.5005
R25878 VSS.n2699 VSS.n2378 4.5005
R25879 VSS.n2701 VSS.n2378 4.5005
R25880 VSS.n2704 VSS.n2378 4.5005
R25881 VSS.n2706 VSS.n2378 4.5005
R25882 VSS.n2707 VSS.n2378 4.5005
R25883 VSS.n2709 VSS.n2378 4.5005
R25884 VSS.n2712 VSS.n2378 4.5005
R25885 VSS.n2714 VSS.n2378 4.5005
R25886 VSS.n2715 VSS.n2378 4.5005
R25887 VSS.n2717 VSS.n2378 4.5005
R25888 VSS.n2720 VSS.n2378 4.5005
R25889 VSS.n2722 VSS.n2378 4.5005
R25890 VSS.n2723 VSS.n2378 4.5005
R25891 VSS.n2725 VSS.n2378 4.5005
R25892 VSS.n2793 VSS.n2378 4.5005
R25893 VSS.n2859 VSS.n2378 4.5005
R25894 VSS.n3051 VSS.n2454 4.5005
R25895 VSS.n2454 VSS.n2351 4.5005
R25896 VSS.n2483 VSS.n2454 4.5005
R25897 VSS.n2484 VSS.n2454 4.5005
R25898 VSS.n2486 VSS.n2454 4.5005
R25899 VSS.n2489 VSS.n2454 4.5005
R25900 VSS.n2491 VSS.n2454 4.5005
R25901 VSS.n2492 VSS.n2454 4.5005
R25902 VSS.n2494 VSS.n2454 4.5005
R25903 VSS.n2497 VSS.n2454 4.5005
R25904 VSS.n2499 VSS.n2454 4.5005
R25905 VSS.n2500 VSS.n2454 4.5005
R25906 VSS.n2502 VSS.n2454 4.5005
R25907 VSS.n2505 VSS.n2454 4.5005
R25908 VSS.n2507 VSS.n2454 4.5005
R25909 VSS.n2508 VSS.n2454 4.5005
R25910 VSS.n2510 VSS.n2454 4.5005
R25911 VSS.n2513 VSS.n2454 4.5005
R25912 VSS.n2515 VSS.n2454 4.5005
R25913 VSS.n2516 VSS.n2454 4.5005
R25914 VSS.n2518 VSS.n2454 4.5005
R25915 VSS.n2521 VSS.n2454 4.5005
R25916 VSS.n2523 VSS.n2454 4.5005
R25917 VSS.n2524 VSS.n2454 4.5005
R25918 VSS.n2526 VSS.n2454 4.5005
R25919 VSS.n2529 VSS.n2454 4.5005
R25920 VSS.n2531 VSS.n2454 4.5005
R25921 VSS.n2532 VSS.n2454 4.5005
R25922 VSS.n2534 VSS.n2454 4.5005
R25923 VSS.n2537 VSS.n2454 4.5005
R25924 VSS.n2539 VSS.n2454 4.5005
R25925 VSS.n2540 VSS.n2454 4.5005
R25926 VSS.n2542 VSS.n2454 4.5005
R25927 VSS.n2545 VSS.n2454 4.5005
R25928 VSS.n2547 VSS.n2454 4.5005
R25929 VSS.n2548 VSS.n2454 4.5005
R25930 VSS.n2550 VSS.n2454 4.5005
R25931 VSS.n2553 VSS.n2454 4.5005
R25932 VSS.n2555 VSS.n2454 4.5005
R25933 VSS.n2556 VSS.n2454 4.5005
R25934 VSS.n2558 VSS.n2454 4.5005
R25935 VSS.n2561 VSS.n2454 4.5005
R25936 VSS.n2563 VSS.n2454 4.5005
R25937 VSS.n2564 VSS.n2454 4.5005
R25938 VSS.n2566 VSS.n2454 4.5005
R25939 VSS.n2569 VSS.n2454 4.5005
R25940 VSS.n2571 VSS.n2454 4.5005
R25941 VSS.n2572 VSS.n2454 4.5005
R25942 VSS.n2574 VSS.n2454 4.5005
R25943 VSS.n2577 VSS.n2454 4.5005
R25944 VSS.n2579 VSS.n2454 4.5005
R25945 VSS.n2580 VSS.n2454 4.5005
R25946 VSS.n2582 VSS.n2454 4.5005
R25947 VSS.n2585 VSS.n2454 4.5005
R25948 VSS.n2587 VSS.n2454 4.5005
R25949 VSS.n2588 VSS.n2454 4.5005
R25950 VSS.n2590 VSS.n2454 4.5005
R25951 VSS.n2593 VSS.n2454 4.5005
R25952 VSS.n2595 VSS.n2454 4.5005
R25953 VSS.n2596 VSS.n2454 4.5005
R25954 VSS.n2598 VSS.n2454 4.5005
R25955 VSS.n2601 VSS.n2454 4.5005
R25956 VSS.n2603 VSS.n2454 4.5005
R25957 VSS.n2604 VSS.n2454 4.5005
R25958 VSS.n2606 VSS.n2454 4.5005
R25959 VSS.n2609 VSS.n2454 4.5005
R25960 VSS.n2611 VSS.n2454 4.5005
R25961 VSS.n2612 VSS.n2454 4.5005
R25962 VSS.n2614 VSS.n2454 4.5005
R25963 VSS.n2617 VSS.n2454 4.5005
R25964 VSS.n2619 VSS.n2454 4.5005
R25965 VSS.n2620 VSS.n2454 4.5005
R25966 VSS.n2622 VSS.n2454 4.5005
R25967 VSS.n2625 VSS.n2454 4.5005
R25968 VSS.n2627 VSS.n2454 4.5005
R25969 VSS.n2628 VSS.n2454 4.5005
R25970 VSS.n2630 VSS.n2454 4.5005
R25971 VSS.n2633 VSS.n2454 4.5005
R25972 VSS.n2635 VSS.n2454 4.5005
R25973 VSS.n2636 VSS.n2454 4.5005
R25974 VSS.n2638 VSS.n2454 4.5005
R25975 VSS.n2640 VSS.n2454 4.5005
R25976 VSS.n2642 VSS.n2454 4.5005
R25977 VSS.n2643 VSS.n2454 4.5005
R25978 VSS.n2645 VSS.n2454 4.5005
R25979 VSS.n2648 VSS.n2454 4.5005
R25980 VSS.n2650 VSS.n2454 4.5005
R25981 VSS.n2651 VSS.n2454 4.5005
R25982 VSS.n2653 VSS.n2454 4.5005
R25983 VSS.n2656 VSS.n2454 4.5005
R25984 VSS.n2658 VSS.n2454 4.5005
R25985 VSS.n2659 VSS.n2454 4.5005
R25986 VSS.n2661 VSS.n2454 4.5005
R25987 VSS.n2664 VSS.n2454 4.5005
R25988 VSS.n2666 VSS.n2454 4.5005
R25989 VSS.n2667 VSS.n2454 4.5005
R25990 VSS.n2669 VSS.n2454 4.5005
R25991 VSS.n2672 VSS.n2454 4.5005
R25992 VSS.n2674 VSS.n2454 4.5005
R25993 VSS.n2675 VSS.n2454 4.5005
R25994 VSS.n2677 VSS.n2454 4.5005
R25995 VSS.n2680 VSS.n2454 4.5005
R25996 VSS.n2682 VSS.n2454 4.5005
R25997 VSS.n2683 VSS.n2454 4.5005
R25998 VSS.n2685 VSS.n2454 4.5005
R25999 VSS.n2688 VSS.n2454 4.5005
R26000 VSS.n2690 VSS.n2454 4.5005
R26001 VSS.n2691 VSS.n2454 4.5005
R26002 VSS.n2693 VSS.n2454 4.5005
R26003 VSS.n2696 VSS.n2454 4.5005
R26004 VSS.n2698 VSS.n2454 4.5005
R26005 VSS.n2699 VSS.n2454 4.5005
R26006 VSS.n2701 VSS.n2454 4.5005
R26007 VSS.n2704 VSS.n2454 4.5005
R26008 VSS.n2706 VSS.n2454 4.5005
R26009 VSS.n2707 VSS.n2454 4.5005
R26010 VSS.n2709 VSS.n2454 4.5005
R26011 VSS.n2712 VSS.n2454 4.5005
R26012 VSS.n2714 VSS.n2454 4.5005
R26013 VSS.n2715 VSS.n2454 4.5005
R26014 VSS.n2717 VSS.n2454 4.5005
R26015 VSS.n2720 VSS.n2454 4.5005
R26016 VSS.n2722 VSS.n2454 4.5005
R26017 VSS.n2723 VSS.n2454 4.5005
R26018 VSS.n2725 VSS.n2454 4.5005
R26019 VSS.n2793 VSS.n2454 4.5005
R26020 VSS.n2859 VSS.n2454 4.5005
R26021 VSS.n3051 VSS.n2377 4.5005
R26022 VSS.n2377 VSS.n2351 4.5005
R26023 VSS.n2483 VSS.n2377 4.5005
R26024 VSS.n2484 VSS.n2377 4.5005
R26025 VSS.n2486 VSS.n2377 4.5005
R26026 VSS.n2489 VSS.n2377 4.5005
R26027 VSS.n2491 VSS.n2377 4.5005
R26028 VSS.n2492 VSS.n2377 4.5005
R26029 VSS.n2494 VSS.n2377 4.5005
R26030 VSS.n2497 VSS.n2377 4.5005
R26031 VSS.n2499 VSS.n2377 4.5005
R26032 VSS.n2500 VSS.n2377 4.5005
R26033 VSS.n2502 VSS.n2377 4.5005
R26034 VSS.n2505 VSS.n2377 4.5005
R26035 VSS.n2507 VSS.n2377 4.5005
R26036 VSS.n2508 VSS.n2377 4.5005
R26037 VSS.n2510 VSS.n2377 4.5005
R26038 VSS.n2513 VSS.n2377 4.5005
R26039 VSS.n2515 VSS.n2377 4.5005
R26040 VSS.n2516 VSS.n2377 4.5005
R26041 VSS.n2518 VSS.n2377 4.5005
R26042 VSS.n2521 VSS.n2377 4.5005
R26043 VSS.n2523 VSS.n2377 4.5005
R26044 VSS.n2524 VSS.n2377 4.5005
R26045 VSS.n2526 VSS.n2377 4.5005
R26046 VSS.n2529 VSS.n2377 4.5005
R26047 VSS.n2531 VSS.n2377 4.5005
R26048 VSS.n2532 VSS.n2377 4.5005
R26049 VSS.n2534 VSS.n2377 4.5005
R26050 VSS.n2537 VSS.n2377 4.5005
R26051 VSS.n2539 VSS.n2377 4.5005
R26052 VSS.n2540 VSS.n2377 4.5005
R26053 VSS.n2542 VSS.n2377 4.5005
R26054 VSS.n2545 VSS.n2377 4.5005
R26055 VSS.n2547 VSS.n2377 4.5005
R26056 VSS.n2548 VSS.n2377 4.5005
R26057 VSS.n2550 VSS.n2377 4.5005
R26058 VSS.n2553 VSS.n2377 4.5005
R26059 VSS.n2555 VSS.n2377 4.5005
R26060 VSS.n2556 VSS.n2377 4.5005
R26061 VSS.n2558 VSS.n2377 4.5005
R26062 VSS.n2561 VSS.n2377 4.5005
R26063 VSS.n2563 VSS.n2377 4.5005
R26064 VSS.n2564 VSS.n2377 4.5005
R26065 VSS.n2566 VSS.n2377 4.5005
R26066 VSS.n2569 VSS.n2377 4.5005
R26067 VSS.n2571 VSS.n2377 4.5005
R26068 VSS.n2572 VSS.n2377 4.5005
R26069 VSS.n2574 VSS.n2377 4.5005
R26070 VSS.n2577 VSS.n2377 4.5005
R26071 VSS.n2579 VSS.n2377 4.5005
R26072 VSS.n2580 VSS.n2377 4.5005
R26073 VSS.n2582 VSS.n2377 4.5005
R26074 VSS.n2585 VSS.n2377 4.5005
R26075 VSS.n2587 VSS.n2377 4.5005
R26076 VSS.n2588 VSS.n2377 4.5005
R26077 VSS.n2590 VSS.n2377 4.5005
R26078 VSS.n2593 VSS.n2377 4.5005
R26079 VSS.n2595 VSS.n2377 4.5005
R26080 VSS.n2596 VSS.n2377 4.5005
R26081 VSS.n2598 VSS.n2377 4.5005
R26082 VSS.n2601 VSS.n2377 4.5005
R26083 VSS.n2603 VSS.n2377 4.5005
R26084 VSS.n2604 VSS.n2377 4.5005
R26085 VSS.n2606 VSS.n2377 4.5005
R26086 VSS.n2609 VSS.n2377 4.5005
R26087 VSS.n2611 VSS.n2377 4.5005
R26088 VSS.n2612 VSS.n2377 4.5005
R26089 VSS.n2614 VSS.n2377 4.5005
R26090 VSS.n2617 VSS.n2377 4.5005
R26091 VSS.n2619 VSS.n2377 4.5005
R26092 VSS.n2620 VSS.n2377 4.5005
R26093 VSS.n2622 VSS.n2377 4.5005
R26094 VSS.n2625 VSS.n2377 4.5005
R26095 VSS.n2627 VSS.n2377 4.5005
R26096 VSS.n2628 VSS.n2377 4.5005
R26097 VSS.n2630 VSS.n2377 4.5005
R26098 VSS.n2633 VSS.n2377 4.5005
R26099 VSS.n2635 VSS.n2377 4.5005
R26100 VSS.n2636 VSS.n2377 4.5005
R26101 VSS.n2638 VSS.n2377 4.5005
R26102 VSS.n2640 VSS.n2377 4.5005
R26103 VSS.n2642 VSS.n2377 4.5005
R26104 VSS.n2643 VSS.n2377 4.5005
R26105 VSS.n2645 VSS.n2377 4.5005
R26106 VSS.n2648 VSS.n2377 4.5005
R26107 VSS.n2650 VSS.n2377 4.5005
R26108 VSS.n2651 VSS.n2377 4.5005
R26109 VSS.n2653 VSS.n2377 4.5005
R26110 VSS.n2656 VSS.n2377 4.5005
R26111 VSS.n2658 VSS.n2377 4.5005
R26112 VSS.n2659 VSS.n2377 4.5005
R26113 VSS.n2661 VSS.n2377 4.5005
R26114 VSS.n2664 VSS.n2377 4.5005
R26115 VSS.n2666 VSS.n2377 4.5005
R26116 VSS.n2667 VSS.n2377 4.5005
R26117 VSS.n2669 VSS.n2377 4.5005
R26118 VSS.n2672 VSS.n2377 4.5005
R26119 VSS.n2674 VSS.n2377 4.5005
R26120 VSS.n2675 VSS.n2377 4.5005
R26121 VSS.n2677 VSS.n2377 4.5005
R26122 VSS.n2680 VSS.n2377 4.5005
R26123 VSS.n2682 VSS.n2377 4.5005
R26124 VSS.n2683 VSS.n2377 4.5005
R26125 VSS.n2685 VSS.n2377 4.5005
R26126 VSS.n2688 VSS.n2377 4.5005
R26127 VSS.n2690 VSS.n2377 4.5005
R26128 VSS.n2691 VSS.n2377 4.5005
R26129 VSS.n2693 VSS.n2377 4.5005
R26130 VSS.n2696 VSS.n2377 4.5005
R26131 VSS.n2698 VSS.n2377 4.5005
R26132 VSS.n2699 VSS.n2377 4.5005
R26133 VSS.n2701 VSS.n2377 4.5005
R26134 VSS.n2704 VSS.n2377 4.5005
R26135 VSS.n2706 VSS.n2377 4.5005
R26136 VSS.n2707 VSS.n2377 4.5005
R26137 VSS.n2709 VSS.n2377 4.5005
R26138 VSS.n2712 VSS.n2377 4.5005
R26139 VSS.n2714 VSS.n2377 4.5005
R26140 VSS.n2715 VSS.n2377 4.5005
R26141 VSS.n2717 VSS.n2377 4.5005
R26142 VSS.n2720 VSS.n2377 4.5005
R26143 VSS.n2722 VSS.n2377 4.5005
R26144 VSS.n2723 VSS.n2377 4.5005
R26145 VSS.n2725 VSS.n2377 4.5005
R26146 VSS.n2793 VSS.n2377 4.5005
R26147 VSS.n2859 VSS.n2377 4.5005
R26148 VSS.n3051 VSS.n2455 4.5005
R26149 VSS.n2455 VSS.n2351 4.5005
R26150 VSS.n2483 VSS.n2455 4.5005
R26151 VSS.n2484 VSS.n2455 4.5005
R26152 VSS.n2486 VSS.n2455 4.5005
R26153 VSS.n2489 VSS.n2455 4.5005
R26154 VSS.n2491 VSS.n2455 4.5005
R26155 VSS.n2492 VSS.n2455 4.5005
R26156 VSS.n2494 VSS.n2455 4.5005
R26157 VSS.n2497 VSS.n2455 4.5005
R26158 VSS.n2499 VSS.n2455 4.5005
R26159 VSS.n2500 VSS.n2455 4.5005
R26160 VSS.n2502 VSS.n2455 4.5005
R26161 VSS.n2505 VSS.n2455 4.5005
R26162 VSS.n2507 VSS.n2455 4.5005
R26163 VSS.n2508 VSS.n2455 4.5005
R26164 VSS.n2510 VSS.n2455 4.5005
R26165 VSS.n2513 VSS.n2455 4.5005
R26166 VSS.n2515 VSS.n2455 4.5005
R26167 VSS.n2516 VSS.n2455 4.5005
R26168 VSS.n2518 VSS.n2455 4.5005
R26169 VSS.n2521 VSS.n2455 4.5005
R26170 VSS.n2523 VSS.n2455 4.5005
R26171 VSS.n2524 VSS.n2455 4.5005
R26172 VSS.n2526 VSS.n2455 4.5005
R26173 VSS.n2529 VSS.n2455 4.5005
R26174 VSS.n2531 VSS.n2455 4.5005
R26175 VSS.n2532 VSS.n2455 4.5005
R26176 VSS.n2534 VSS.n2455 4.5005
R26177 VSS.n2537 VSS.n2455 4.5005
R26178 VSS.n2539 VSS.n2455 4.5005
R26179 VSS.n2540 VSS.n2455 4.5005
R26180 VSS.n2542 VSS.n2455 4.5005
R26181 VSS.n2545 VSS.n2455 4.5005
R26182 VSS.n2547 VSS.n2455 4.5005
R26183 VSS.n2548 VSS.n2455 4.5005
R26184 VSS.n2550 VSS.n2455 4.5005
R26185 VSS.n2553 VSS.n2455 4.5005
R26186 VSS.n2555 VSS.n2455 4.5005
R26187 VSS.n2556 VSS.n2455 4.5005
R26188 VSS.n2558 VSS.n2455 4.5005
R26189 VSS.n2561 VSS.n2455 4.5005
R26190 VSS.n2563 VSS.n2455 4.5005
R26191 VSS.n2564 VSS.n2455 4.5005
R26192 VSS.n2566 VSS.n2455 4.5005
R26193 VSS.n2569 VSS.n2455 4.5005
R26194 VSS.n2571 VSS.n2455 4.5005
R26195 VSS.n2572 VSS.n2455 4.5005
R26196 VSS.n2574 VSS.n2455 4.5005
R26197 VSS.n2577 VSS.n2455 4.5005
R26198 VSS.n2579 VSS.n2455 4.5005
R26199 VSS.n2580 VSS.n2455 4.5005
R26200 VSS.n2582 VSS.n2455 4.5005
R26201 VSS.n2585 VSS.n2455 4.5005
R26202 VSS.n2587 VSS.n2455 4.5005
R26203 VSS.n2588 VSS.n2455 4.5005
R26204 VSS.n2590 VSS.n2455 4.5005
R26205 VSS.n2593 VSS.n2455 4.5005
R26206 VSS.n2595 VSS.n2455 4.5005
R26207 VSS.n2596 VSS.n2455 4.5005
R26208 VSS.n2598 VSS.n2455 4.5005
R26209 VSS.n2601 VSS.n2455 4.5005
R26210 VSS.n2603 VSS.n2455 4.5005
R26211 VSS.n2604 VSS.n2455 4.5005
R26212 VSS.n2606 VSS.n2455 4.5005
R26213 VSS.n2609 VSS.n2455 4.5005
R26214 VSS.n2611 VSS.n2455 4.5005
R26215 VSS.n2612 VSS.n2455 4.5005
R26216 VSS.n2614 VSS.n2455 4.5005
R26217 VSS.n2617 VSS.n2455 4.5005
R26218 VSS.n2619 VSS.n2455 4.5005
R26219 VSS.n2620 VSS.n2455 4.5005
R26220 VSS.n2622 VSS.n2455 4.5005
R26221 VSS.n2625 VSS.n2455 4.5005
R26222 VSS.n2627 VSS.n2455 4.5005
R26223 VSS.n2628 VSS.n2455 4.5005
R26224 VSS.n2630 VSS.n2455 4.5005
R26225 VSS.n2633 VSS.n2455 4.5005
R26226 VSS.n2635 VSS.n2455 4.5005
R26227 VSS.n2636 VSS.n2455 4.5005
R26228 VSS.n2638 VSS.n2455 4.5005
R26229 VSS.n2640 VSS.n2455 4.5005
R26230 VSS.n2642 VSS.n2455 4.5005
R26231 VSS.n2643 VSS.n2455 4.5005
R26232 VSS.n2645 VSS.n2455 4.5005
R26233 VSS.n2648 VSS.n2455 4.5005
R26234 VSS.n2650 VSS.n2455 4.5005
R26235 VSS.n2651 VSS.n2455 4.5005
R26236 VSS.n2653 VSS.n2455 4.5005
R26237 VSS.n2656 VSS.n2455 4.5005
R26238 VSS.n2658 VSS.n2455 4.5005
R26239 VSS.n2659 VSS.n2455 4.5005
R26240 VSS.n2661 VSS.n2455 4.5005
R26241 VSS.n2664 VSS.n2455 4.5005
R26242 VSS.n2666 VSS.n2455 4.5005
R26243 VSS.n2667 VSS.n2455 4.5005
R26244 VSS.n2669 VSS.n2455 4.5005
R26245 VSS.n2672 VSS.n2455 4.5005
R26246 VSS.n2674 VSS.n2455 4.5005
R26247 VSS.n2675 VSS.n2455 4.5005
R26248 VSS.n2677 VSS.n2455 4.5005
R26249 VSS.n2680 VSS.n2455 4.5005
R26250 VSS.n2682 VSS.n2455 4.5005
R26251 VSS.n2683 VSS.n2455 4.5005
R26252 VSS.n2685 VSS.n2455 4.5005
R26253 VSS.n2688 VSS.n2455 4.5005
R26254 VSS.n2690 VSS.n2455 4.5005
R26255 VSS.n2691 VSS.n2455 4.5005
R26256 VSS.n2693 VSS.n2455 4.5005
R26257 VSS.n2696 VSS.n2455 4.5005
R26258 VSS.n2698 VSS.n2455 4.5005
R26259 VSS.n2699 VSS.n2455 4.5005
R26260 VSS.n2701 VSS.n2455 4.5005
R26261 VSS.n2704 VSS.n2455 4.5005
R26262 VSS.n2706 VSS.n2455 4.5005
R26263 VSS.n2707 VSS.n2455 4.5005
R26264 VSS.n2709 VSS.n2455 4.5005
R26265 VSS.n2712 VSS.n2455 4.5005
R26266 VSS.n2714 VSS.n2455 4.5005
R26267 VSS.n2715 VSS.n2455 4.5005
R26268 VSS.n2717 VSS.n2455 4.5005
R26269 VSS.n2720 VSS.n2455 4.5005
R26270 VSS.n2722 VSS.n2455 4.5005
R26271 VSS.n2723 VSS.n2455 4.5005
R26272 VSS.n2725 VSS.n2455 4.5005
R26273 VSS.n2793 VSS.n2455 4.5005
R26274 VSS.n2859 VSS.n2455 4.5005
R26275 VSS.n3051 VSS.n2376 4.5005
R26276 VSS.n2376 VSS.n2351 4.5005
R26277 VSS.n2483 VSS.n2376 4.5005
R26278 VSS.n2484 VSS.n2376 4.5005
R26279 VSS.n2486 VSS.n2376 4.5005
R26280 VSS.n2489 VSS.n2376 4.5005
R26281 VSS.n2491 VSS.n2376 4.5005
R26282 VSS.n2492 VSS.n2376 4.5005
R26283 VSS.n2494 VSS.n2376 4.5005
R26284 VSS.n2497 VSS.n2376 4.5005
R26285 VSS.n2499 VSS.n2376 4.5005
R26286 VSS.n2500 VSS.n2376 4.5005
R26287 VSS.n2502 VSS.n2376 4.5005
R26288 VSS.n2505 VSS.n2376 4.5005
R26289 VSS.n2507 VSS.n2376 4.5005
R26290 VSS.n2508 VSS.n2376 4.5005
R26291 VSS.n2510 VSS.n2376 4.5005
R26292 VSS.n2513 VSS.n2376 4.5005
R26293 VSS.n2515 VSS.n2376 4.5005
R26294 VSS.n2516 VSS.n2376 4.5005
R26295 VSS.n2518 VSS.n2376 4.5005
R26296 VSS.n2521 VSS.n2376 4.5005
R26297 VSS.n2523 VSS.n2376 4.5005
R26298 VSS.n2524 VSS.n2376 4.5005
R26299 VSS.n2526 VSS.n2376 4.5005
R26300 VSS.n2529 VSS.n2376 4.5005
R26301 VSS.n2531 VSS.n2376 4.5005
R26302 VSS.n2532 VSS.n2376 4.5005
R26303 VSS.n2534 VSS.n2376 4.5005
R26304 VSS.n2537 VSS.n2376 4.5005
R26305 VSS.n2539 VSS.n2376 4.5005
R26306 VSS.n2540 VSS.n2376 4.5005
R26307 VSS.n2542 VSS.n2376 4.5005
R26308 VSS.n2545 VSS.n2376 4.5005
R26309 VSS.n2547 VSS.n2376 4.5005
R26310 VSS.n2548 VSS.n2376 4.5005
R26311 VSS.n2550 VSS.n2376 4.5005
R26312 VSS.n2553 VSS.n2376 4.5005
R26313 VSS.n2555 VSS.n2376 4.5005
R26314 VSS.n2556 VSS.n2376 4.5005
R26315 VSS.n2558 VSS.n2376 4.5005
R26316 VSS.n2561 VSS.n2376 4.5005
R26317 VSS.n2563 VSS.n2376 4.5005
R26318 VSS.n2564 VSS.n2376 4.5005
R26319 VSS.n2566 VSS.n2376 4.5005
R26320 VSS.n2569 VSS.n2376 4.5005
R26321 VSS.n2571 VSS.n2376 4.5005
R26322 VSS.n2572 VSS.n2376 4.5005
R26323 VSS.n2574 VSS.n2376 4.5005
R26324 VSS.n2577 VSS.n2376 4.5005
R26325 VSS.n2579 VSS.n2376 4.5005
R26326 VSS.n2580 VSS.n2376 4.5005
R26327 VSS.n2582 VSS.n2376 4.5005
R26328 VSS.n2585 VSS.n2376 4.5005
R26329 VSS.n2587 VSS.n2376 4.5005
R26330 VSS.n2588 VSS.n2376 4.5005
R26331 VSS.n2590 VSS.n2376 4.5005
R26332 VSS.n2593 VSS.n2376 4.5005
R26333 VSS.n2595 VSS.n2376 4.5005
R26334 VSS.n2596 VSS.n2376 4.5005
R26335 VSS.n2598 VSS.n2376 4.5005
R26336 VSS.n2601 VSS.n2376 4.5005
R26337 VSS.n2603 VSS.n2376 4.5005
R26338 VSS.n2604 VSS.n2376 4.5005
R26339 VSS.n2606 VSS.n2376 4.5005
R26340 VSS.n2609 VSS.n2376 4.5005
R26341 VSS.n2611 VSS.n2376 4.5005
R26342 VSS.n2612 VSS.n2376 4.5005
R26343 VSS.n2614 VSS.n2376 4.5005
R26344 VSS.n2617 VSS.n2376 4.5005
R26345 VSS.n2619 VSS.n2376 4.5005
R26346 VSS.n2620 VSS.n2376 4.5005
R26347 VSS.n2622 VSS.n2376 4.5005
R26348 VSS.n2625 VSS.n2376 4.5005
R26349 VSS.n2627 VSS.n2376 4.5005
R26350 VSS.n2628 VSS.n2376 4.5005
R26351 VSS.n2630 VSS.n2376 4.5005
R26352 VSS.n2633 VSS.n2376 4.5005
R26353 VSS.n2635 VSS.n2376 4.5005
R26354 VSS.n2636 VSS.n2376 4.5005
R26355 VSS.n2638 VSS.n2376 4.5005
R26356 VSS.n2640 VSS.n2376 4.5005
R26357 VSS.n2642 VSS.n2376 4.5005
R26358 VSS.n2643 VSS.n2376 4.5005
R26359 VSS.n2645 VSS.n2376 4.5005
R26360 VSS.n2648 VSS.n2376 4.5005
R26361 VSS.n2650 VSS.n2376 4.5005
R26362 VSS.n2651 VSS.n2376 4.5005
R26363 VSS.n2653 VSS.n2376 4.5005
R26364 VSS.n2656 VSS.n2376 4.5005
R26365 VSS.n2658 VSS.n2376 4.5005
R26366 VSS.n2659 VSS.n2376 4.5005
R26367 VSS.n2661 VSS.n2376 4.5005
R26368 VSS.n2664 VSS.n2376 4.5005
R26369 VSS.n2666 VSS.n2376 4.5005
R26370 VSS.n2667 VSS.n2376 4.5005
R26371 VSS.n2669 VSS.n2376 4.5005
R26372 VSS.n2672 VSS.n2376 4.5005
R26373 VSS.n2674 VSS.n2376 4.5005
R26374 VSS.n2675 VSS.n2376 4.5005
R26375 VSS.n2677 VSS.n2376 4.5005
R26376 VSS.n2680 VSS.n2376 4.5005
R26377 VSS.n2682 VSS.n2376 4.5005
R26378 VSS.n2683 VSS.n2376 4.5005
R26379 VSS.n2685 VSS.n2376 4.5005
R26380 VSS.n2688 VSS.n2376 4.5005
R26381 VSS.n2690 VSS.n2376 4.5005
R26382 VSS.n2691 VSS.n2376 4.5005
R26383 VSS.n2693 VSS.n2376 4.5005
R26384 VSS.n2696 VSS.n2376 4.5005
R26385 VSS.n2698 VSS.n2376 4.5005
R26386 VSS.n2699 VSS.n2376 4.5005
R26387 VSS.n2701 VSS.n2376 4.5005
R26388 VSS.n2704 VSS.n2376 4.5005
R26389 VSS.n2706 VSS.n2376 4.5005
R26390 VSS.n2707 VSS.n2376 4.5005
R26391 VSS.n2709 VSS.n2376 4.5005
R26392 VSS.n2712 VSS.n2376 4.5005
R26393 VSS.n2714 VSS.n2376 4.5005
R26394 VSS.n2715 VSS.n2376 4.5005
R26395 VSS.n2717 VSS.n2376 4.5005
R26396 VSS.n2720 VSS.n2376 4.5005
R26397 VSS.n2722 VSS.n2376 4.5005
R26398 VSS.n2723 VSS.n2376 4.5005
R26399 VSS.n2725 VSS.n2376 4.5005
R26400 VSS.n2793 VSS.n2376 4.5005
R26401 VSS.n2859 VSS.n2376 4.5005
R26402 VSS.n3051 VSS.n2456 4.5005
R26403 VSS.n2456 VSS.n2351 4.5005
R26404 VSS.n2483 VSS.n2456 4.5005
R26405 VSS.n2484 VSS.n2456 4.5005
R26406 VSS.n2486 VSS.n2456 4.5005
R26407 VSS.n2489 VSS.n2456 4.5005
R26408 VSS.n2491 VSS.n2456 4.5005
R26409 VSS.n2492 VSS.n2456 4.5005
R26410 VSS.n2494 VSS.n2456 4.5005
R26411 VSS.n2497 VSS.n2456 4.5005
R26412 VSS.n2499 VSS.n2456 4.5005
R26413 VSS.n2500 VSS.n2456 4.5005
R26414 VSS.n2502 VSS.n2456 4.5005
R26415 VSS.n2505 VSS.n2456 4.5005
R26416 VSS.n2507 VSS.n2456 4.5005
R26417 VSS.n2508 VSS.n2456 4.5005
R26418 VSS.n2510 VSS.n2456 4.5005
R26419 VSS.n2513 VSS.n2456 4.5005
R26420 VSS.n2515 VSS.n2456 4.5005
R26421 VSS.n2516 VSS.n2456 4.5005
R26422 VSS.n2518 VSS.n2456 4.5005
R26423 VSS.n2521 VSS.n2456 4.5005
R26424 VSS.n2523 VSS.n2456 4.5005
R26425 VSS.n2524 VSS.n2456 4.5005
R26426 VSS.n2526 VSS.n2456 4.5005
R26427 VSS.n2529 VSS.n2456 4.5005
R26428 VSS.n2531 VSS.n2456 4.5005
R26429 VSS.n2532 VSS.n2456 4.5005
R26430 VSS.n2534 VSS.n2456 4.5005
R26431 VSS.n2537 VSS.n2456 4.5005
R26432 VSS.n2539 VSS.n2456 4.5005
R26433 VSS.n2540 VSS.n2456 4.5005
R26434 VSS.n2542 VSS.n2456 4.5005
R26435 VSS.n2545 VSS.n2456 4.5005
R26436 VSS.n2547 VSS.n2456 4.5005
R26437 VSS.n2548 VSS.n2456 4.5005
R26438 VSS.n2550 VSS.n2456 4.5005
R26439 VSS.n2553 VSS.n2456 4.5005
R26440 VSS.n2555 VSS.n2456 4.5005
R26441 VSS.n2556 VSS.n2456 4.5005
R26442 VSS.n2558 VSS.n2456 4.5005
R26443 VSS.n2561 VSS.n2456 4.5005
R26444 VSS.n2563 VSS.n2456 4.5005
R26445 VSS.n2564 VSS.n2456 4.5005
R26446 VSS.n2566 VSS.n2456 4.5005
R26447 VSS.n2569 VSS.n2456 4.5005
R26448 VSS.n2571 VSS.n2456 4.5005
R26449 VSS.n2572 VSS.n2456 4.5005
R26450 VSS.n2574 VSS.n2456 4.5005
R26451 VSS.n2577 VSS.n2456 4.5005
R26452 VSS.n2579 VSS.n2456 4.5005
R26453 VSS.n2580 VSS.n2456 4.5005
R26454 VSS.n2582 VSS.n2456 4.5005
R26455 VSS.n2585 VSS.n2456 4.5005
R26456 VSS.n2587 VSS.n2456 4.5005
R26457 VSS.n2588 VSS.n2456 4.5005
R26458 VSS.n2590 VSS.n2456 4.5005
R26459 VSS.n2593 VSS.n2456 4.5005
R26460 VSS.n2595 VSS.n2456 4.5005
R26461 VSS.n2596 VSS.n2456 4.5005
R26462 VSS.n2598 VSS.n2456 4.5005
R26463 VSS.n2601 VSS.n2456 4.5005
R26464 VSS.n2603 VSS.n2456 4.5005
R26465 VSS.n2604 VSS.n2456 4.5005
R26466 VSS.n2606 VSS.n2456 4.5005
R26467 VSS.n2609 VSS.n2456 4.5005
R26468 VSS.n2611 VSS.n2456 4.5005
R26469 VSS.n2612 VSS.n2456 4.5005
R26470 VSS.n2614 VSS.n2456 4.5005
R26471 VSS.n2617 VSS.n2456 4.5005
R26472 VSS.n2619 VSS.n2456 4.5005
R26473 VSS.n2620 VSS.n2456 4.5005
R26474 VSS.n2622 VSS.n2456 4.5005
R26475 VSS.n2625 VSS.n2456 4.5005
R26476 VSS.n2627 VSS.n2456 4.5005
R26477 VSS.n2628 VSS.n2456 4.5005
R26478 VSS.n2630 VSS.n2456 4.5005
R26479 VSS.n2633 VSS.n2456 4.5005
R26480 VSS.n2635 VSS.n2456 4.5005
R26481 VSS.n2636 VSS.n2456 4.5005
R26482 VSS.n2638 VSS.n2456 4.5005
R26483 VSS.n2640 VSS.n2456 4.5005
R26484 VSS.n2642 VSS.n2456 4.5005
R26485 VSS.n2643 VSS.n2456 4.5005
R26486 VSS.n2645 VSS.n2456 4.5005
R26487 VSS.n2648 VSS.n2456 4.5005
R26488 VSS.n2650 VSS.n2456 4.5005
R26489 VSS.n2651 VSS.n2456 4.5005
R26490 VSS.n2653 VSS.n2456 4.5005
R26491 VSS.n2656 VSS.n2456 4.5005
R26492 VSS.n2658 VSS.n2456 4.5005
R26493 VSS.n2659 VSS.n2456 4.5005
R26494 VSS.n2661 VSS.n2456 4.5005
R26495 VSS.n2664 VSS.n2456 4.5005
R26496 VSS.n2666 VSS.n2456 4.5005
R26497 VSS.n2667 VSS.n2456 4.5005
R26498 VSS.n2669 VSS.n2456 4.5005
R26499 VSS.n2672 VSS.n2456 4.5005
R26500 VSS.n2674 VSS.n2456 4.5005
R26501 VSS.n2675 VSS.n2456 4.5005
R26502 VSS.n2677 VSS.n2456 4.5005
R26503 VSS.n2680 VSS.n2456 4.5005
R26504 VSS.n2682 VSS.n2456 4.5005
R26505 VSS.n2683 VSS.n2456 4.5005
R26506 VSS.n2685 VSS.n2456 4.5005
R26507 VSS.n2688 VSS.n2456 4.5005
R26508 VSS.n2690 VSS.n2456 4.5005
R26509 VSS.n2691 VSS.n2456 4.5005
R26510 VSS.n2693 VSS.n2456 4.5005
R26511 VSS.n2696 VSS.n2456 4.5005
R26512 VSS.n2698 VSS.n2456 4.5005
R26513 VSS.n2699 VSS.n2456 4.5005
R26514 VSS.n2701 VSS.n2456 4.5005
R26515 VSS.n2704 VSS.n2456 4.5005
R26516 VSS.n2706 VSS.n2456 4.5005
R26517 VSS.n2707 VSS.n2456 4.5005
R26518 VSS.n2709 VSS.n2456 4.5005
R26519 VSS.n2712 VSS.n2456 4.5005
R26520 VSS.n2714 VSS.n2456 4.5005
R26521 VSS.n2715 VSS.n2456 4.5005
R26522 VSS.n2717 VSS.n2456 4.5005
R26523 VSS.n2720 VSS.n2456 4.5005
R26524 VSS.n2722 VSS.n2456 4.5005
R26525 VSS.n2723 VSS.n2456 4.5005
R26526 VSS.n2725 VSS.n2456 4.5005
R26527 VSS.n2793 VSS.n2456 4.5005
R26528 VSS.n2859 VSS.n2456 4.5005
R26529 VSS.n3051 VSS.n2375 4.5005
R26530 VSS.n2375 VSS.n2351 4.5005
R26531 VSS.n2483 VSS.n2375 4.5005
R26532 VSS.n2484 VSS.n2375 4.5005
R26533 VSS.n2486 VSS.n2375 4.5005
R26534 VSS.n2489 VSS.n2375 4.5005
R26535 VSS.n2491 VSS.n2375 4.5005
R26536 VSS.n2492 VSS.n2375 4.5005
R26537 VSS.n2494 VSS.n2375 4.5005
R26538 VSS.n2497 VSS.n2375 4.5005
R26539 VSS.n2499 VSS.n2375 4.5005
R26540 VSS.n2500 VSS.n2375 4.5005
R26541 VSS.n2502 VSS.n2375 4.5005
R26542 VSS.n2505 VSS.n2375 4.5005
R26543 VSS.n2507 VSS.n2375 4.5005
R26544 VSS.n2508 VSS.n2375 4.5005
R26545 VSS.n2510 VSS.n2375 4.5005
R26546 VSS.n2513 VSS.n2375 4.5005
R26547 VSS.n2515 VSS.n2375 4.5005
R26548 VSS.n2516 VSS.n2375 4.5005
R26549 VSS.n2518 VSS.n2375 4.5005
R26550 VSS.n2521 VSS.n2375 4.5005
R26551 VSS.n2523 VSS.n2375 4.5005
R26552 VSS.n2524 VSS.n2375 4.5005
R26553 VSS.n2526 VSS.n2375 4.5005
R26554 VSS.n2529 VSS.n2375 4.5005
R26555 VSS.n2531 VSS.n2375 4.5005
R26556 VSS.n2532 VSS.n2375 4.5005
R26557 VSS.n2534 VSS.n2375 4.5005
R26558 VSS.n2537 VSS.n2375 4.5005
R26559 VSS.n2539 VSS.n2375 4.5005
R26560 VSS.n2540 VSS.n2375 4.5005
R26561 VSS.n2542 VSS.n2375 4.5005
R26562 VSS.n2545 VSS.n2375 4.5005
R26563 VSS.n2547 VSS.n2375 4.5005
R26564 VSS.n2548 VSS.n2375 4.5005
R26565 VSS.n2550 VSS.n2375 4.5005
R26566 VSS.n2553 VSS.n2375 4.5005
R26567 VSS.n2555 VSS.n2375 4.5005
R26568 VSS.n2556 VSS.n2375 4.5005
R26569 VSS.n2558 VSS.n2375 4.5005
R26570 VSS.n2561 VSS.n2375 4.5005
R26571 VSS.n2563 VSS.n2375 4.5005
R26572 VSS.n2564 VSS.n2375 4.5005
R26573 VSS.n2566 VSS.n2375 4.5005
R26574 VSS.n2569 VSS.n2375 4.5005
R26575 VSS.n2571 VSS.n2375 4.5005
R26576 VSS.n2572 VSS.n2375 4.5005
R26577 VSS.n2574 VSS.n2375 4.5005
R26578 VSS.n2577 VSS.n2375 4.5005
R26579 VSS.n2579 VSS.n2375 4.5005
R26580 VSS.n2580 VSS.n2375 4.5005
R26581 VSS.n2582 VSS.n2375 4.5005
R26582 VSS.n2585 VSS.n2375 4.5005
R26583 VSS.n2587 VSS.n2375 4.5005
R26584 VSS.n2588 VSS.n2375 4.5005
R26585 VSS.n2590 VSS.n2375 4.5005
R26586 VSS.n2593 VSS.n2375 4.5005
R26587 VSS.n2595 VSS.n2375 4.5005
R26588 VSS.n2596 VSS.n2375 4.5005
R26589 VSS.n2598 VSS.n2375 4.5005
R26590 VSS.n2601 VSS.n2375 4.5005
R26591 VSS.n2603 VSS.n2375 4.5005
R26592 VSS.n2604 VSS.n2375 4.5005
R26593 VSS.n2606 VSS.n2375 4.5005
R26594 VSS.n2609 VSS.n2375 4.5005
R26595 VSS.n2611 VSS.n2375 4.5005
R26596 VSS.n2612 VSS.n2375 4.5005
R26597 VSS.n2614 VSS.n2375 4.5005
R26598 VSS.n2617 VSS.n2375 4.5005
R26599 VSS.n2619 VSS.n2375 4.5005
R26600 VSS.n2620 VSS.n2375 4.5005
R26601 VSS.n2622 VSS.n2375 4.5005
R26602 VSS.n2625 VSS.n2375 4.5005
R26603 VSS.n2627 VSS.n2375 4.5005
R26604 VSS.n2628 VSS.n2375 4.5005
R26605 VSS.n2630 VSS.n2375 4.5005
R26606 VSS.n2633 VSS.n2375 4.5005
R26607 VSS.n2635 VSS.n2375 4.5005
R26608 VSS.n2636 VSS.n2375 4.5005
R26609 VSS.n2638 VSS.n2375 4.5005
R26610 VSS.n2640 VSS.n2375 4.5005
R26611 VSS.n2642 VSS.n2375 4.5005
R26612 VSS.n2643 VSS.n2375 4.5005
R26613 VSS.n2645 VSS.n2375 4.5005
R26614 VSS.n2648 VSS.n2375 4.5005
R26615 VSS.n2650 VSS.n2375 4.5005
R26616 VSS.n2651 VSS.n2375 4.5005
R26617 VSS.n2653 VSS.n2375 4.5005
R26618 VSS.n2656 VSS.n2375 4.5005
R26619 VSS.n2658 VSS.n2375 4.5005
R26620 VSS.n2659 VSS.n2375 4.5005
R26621 VSS.n2661 VSS.n2375 4.5005
R26622 VSS.n2664 VSS.n2375 4.5005
R26623 VSS.n2666 VSS.n2375 4.5005
R26624 VSS.n2667 VSS.n2375 4.5005
R26625 VSS.n2669 VSS.n2375 4.5005
R26626 VSS.n2672 VSS.n2375 4.5005
R26627 VSS.n2674 VSS.n2375 4.5005
R26628 VSS.n2675 VSS.n2375 4.5005
R26629 VSS.n2677 VSS.n2375 4.5005
R26630 VSS.n2680 VSS.n2375 4.5005
R26631 VSS.n2682 VSS.n2375 4.5005
R26632 VSS.n2683 VSS.n2375 4.5005
R26633 VSS.n2685 VSS.n2375 4.5005
R26634 VSS.n2688 VSS.n2375 4.5005
R26635 VSS.n2690 VSS.n2375 4.5005
R26636 VSS.n2691 VSS.n2375 4.5005
R26637 VSS.n2693 VSS.n2375 4.5005
R26638 VSS.n2696 VSS.n2375 4.5005
R26639 VSS.n2698 VSS.n2375 4.5005
R26640 VSS.n2699 VSS.n2375 4.5005
R26641 VSS.n2701 VSS.n2375 4.5005
R26642 VSS.n2704 VSS.n2375 4.5005
R26643 VSS.n2706 VSS.n2375 4.5005
R26644 VSS.n2707 VSS.n2375 4.5005
R26645 VSS.n2709 VSS.n2375 4.5005
R26646 VSS.n2712 VSS.n2375 4.5005
R26647 VSS.n2714 VSS.n2375 4.5005
R26648 VSS.n2715 VSS.n2375 4.5005
R26649 VSS.n2717 VSS.n2375 4.5005
R26650 VSS.n2720 VSS.n2375 4.5005
R26651 VSS.n2722 VSS.n2375 4.5005
R26652 VSS.n2723 VSS.n2375 4.5005
R26653 VSS.n2725 VSS.n2375 4.5005
R26654 VSS.n2793 VSS.n2375 4.5005
R26655 VSS.n2859 VSS.n2375 4.5005
R26656 VSS.n3051 VSS.n2457 4.5005
R26657 VSS.n2457 VSS.n2351 4.5005
R26658 VSS.n2483 VSS.n2457 4.5005
R26659 VSS.n2484 VSS.n2457 4.5005
R26660 VSS.n2486 VSS.n2457 4.5005
R26661 VSS.n2489 VSS.n2457 4.5005
R26662 VSS.n2491 VSS.n2457 4.5005
R26663 VSS.n2492 VSS.n2457 4.5005
R26664 VSS.n2494 VSS.n2457 4.5005
R26665 VSS.n2497 VSS.n2457 4.5005
R26666 VSS.n2499 VSS.n2457 4.5005
R26667 VSS.n2500 VSS.n2457 4.5005
R26668 VSS.n2502 VSS.n2457 4.5005
R26669 VSS.n2505 VSS.n2457 4.5005
R26670 VSS.n2507 VSS.n2457 4.5005
R26671 VSS.n2508 VSS.n2457 4.5005
R26672 VSS.n2510 VSS.n2457 4.5005
R26673 VSS.n2513 VSS.n2457 4.5005
R26674 VSS.n2515 VSS.n2457 4.5005
R26675 VSS.n2516 VSS.n2457 4.5005
R26676 VSS.n2518 VSS.n2457 4.5005
R26677 VSS.n2521 VSS.n2457 4.5005
R26678 VSS.n2523 VSS.n2457 4.5005
R26679 VSS.n2524 VSS.n2457 4.5005
R26680 VSS.n2526 VSS.n2457 4.5005
R26681 VSS.n2529 VSS.n2457 4.5005
R26682 VSS.n2531 VSS.n2457 4.5005
R26683 VSS.n2532 VSS.n2457 4.5005
R26684 VSS.n2534 VSS.n2457 4.5005
R26685 VSS.n2537 VSS.n2457 4.5005
R26686 VSS.n2539 VSS.n2457 4.5005
R26687 VSS.n2540 VSS.n2457 4.5005
R26688 VSS.n2542 VSS.n2457 4.5005
R26689 VSS.n2545 VSS.n2457 4.5005
R26690 VSS.n2547 VSS.n2457 4.5005
R26691 VSS.n2548 VSS.n2457 4.5005
R26692 VSS.n2550 VSS.n2457 4.5005
R26693 VSS.n2553 VSS.n2457 4.5005
R26694 VSS.n2555 VSS.n2457 4.5005
R26695 VSS.n2556 VSS.n2457 4.5005
R26696 VSS.n2558 VSS.n2457 4.5005
R26697 VSS.n2561 VSS.n2457 4.5005
R26698 VSS.n2563 VSS.n2457 4.5005
R26699 VSS.n2564 VSS.n2457 4.5005
R26700 VSS.n2566 VSS.n2457 4.5005
R26701 VSS.n2569 VSS.n2457 4.5005
R26702 VSS.n2571 VSS.n2457 4.5005
R26703 VSS.n2572 VSS.n2457 4.5005
R26704 VSS.n2574 VSS.n2457 4.5005
R26705 VSS.n2577 VSS.n2457 4.5005
R26706 VSS.n2579 VSS.n2457 4.5005
R26707 VSS.n2580 VSS.n2457 4.5005
R26708 VSS.n2582 VSS.n2457 4.5005
R26709 VSS.n2585 VSS.n2457 4.5005
R26710 VSS.n2587 VSS.n2457 4.5005
R26711 VSS.n2588 VSS.n2457 4.5005
R26712 VSS.n2590 VSS.n2457 4.5005
R26713 VSS.n2593 VSS.n2457 4.5005
R26714 VSS.n2595 VSS.n2457 4.5005
R26715 VSS.n2596 VSS.n2457 4.5005
R26716 VSS.n2598 VSS.n2457 4.5005
R26717 VSS.n2601 VSS.n2457 4.5005
R26718 VSS.n2603 VSS.n2457 4.5005
R26719 VSS.n2604 VSS.n2457 4.5005
R26720 VSS.n2606 VSS.n2457 4.5005
R26721 VSS.n2609 VSS.n2457 4.5005
R26722 VSS.n2611 VSS.n2457 4.5005
R26723 VSS.n2612 VSS.n2457 4.5005
R26724 VSS.n2614 VSS.n2457 4.5005
R26725 VSS.n2617 VSS.n2457 4.5005
R26726 VSS.n2619 VSS.n2457 4.5005
R26727 VSS.n2620 VSS.n2457 4.5005
R26728 VSS.n2622 VSS.n2457 4.5005
R26729 VSS.n2625 VSS.n2457 4.5005
R26730 VSS.n2627 VSS.n2457 4.5005
R26731 VSS.n2628 VSS.n2457 4.5005
R26732 VSS.n2630 VSS.n2457 4.5005
R26733 VSS.n2633 VSS.n2457 4.5005
R26734 VSS.n2635 VSS.n2457 4.5005
R26735 VSS.n2636 VSS.n2457 4.5005
R26736 VSS.n2638 VSS.n2457 4.5005
R26737 VSS.n2640 VSS.n2457 4.5005
R26738 VSS.n2642 VSS.n2457 4.5005
R26739 VSS.n2643 VSS.n2457 4.5005
R26740 VSS.n2645 VSS.n2457 4.5005
R26741 VSS.n2648 VSS.n2457 4.5005
R26742 VSS.n2650 VSS.n2457 4.5005
R26743 VSS.n2651 VSS.n2457 4.5005
R26744 VSS.n2653 VSS.n2457 4.5005
R26745 VSS.n2656 VSS.n2457 4.5005
R26746 VSS.n2658 VSS.n2457 4.5005
R26747 VSS.n2659 VSS.n2457 4.5005
R26748 VSS.n2661 VSS.n2457 4.5005
R26749 VSS.n2664 VSS.n2457 4.5005
R26750 VSS.n2666 VSS.n2457 4.5005
R26751 VSS.n2667 VSS.n2457 4.5005
R26752 VSS.n2669 VSS.n2457 4.5005
R26753 VSS.n2672 VSS.n2457 4.5005
R26754 VSS.n2674 VSS.n2457 4.5005
R26755 VSS.n2675 VSS.n2457 4.5005
R26756 VSS.n2677 VSS.n2457 4.5005
R26757 VSS.n2680 VSS.n2457 4.5005
R26758 VSS.n2682 VSS.n2457 4.5005
R26759 VSS.n2683 VSS.n2457 4.5005
R26760 VSS.n2685 VSS.n2457 4.5005
R26761 VSS.n2688 VSS.n2457 4.5005
R26762 VSS.n2690 VSS.n2457 4.5005
R26763 VSS.n2691 VSS.n2457 4.5005
R26764 VSS.n2693 VSS.n2457 4.5005
R26765 VSS.n2696 VSS.n2457 4.5005
R26766 VSS.n2698 VSS.n2457 4.5005
R26767 VSS.n2699 VSS.n2457 4.5005
R26768 VSS.n2701 VSS.n2457 4.5005
R26769 VSS.n2704 VSS.n2457 4.5005
R26770 VSS.n2706 VSS.n2457 4.5005
R26771 VSS.n2707 VSS.n2457 4.5005
R26772 VSS.n2709 VSS.n2457 4.5005
R26773 VSS.n2712 VSS.n2457 4.5005
R26774 VSS.n2714 VSS.n2457 4.5005
R26775 VSS.n2715 VSS.n2457 4.5005
R26776 VSS.n2717 VSS.n2457 4.5005
R26777 VSS.n2720 VSS.n2457 4.5005
R26778 VSS.n2722 VSS.n2457 4.5005
R26779 VSS.n2723 VSS.n2457 4.5005
R26780 VSS.n2725 VSS.n2457 4.5005
R26781 VSS.n2793 VSS.n2457 4.5005
R26782 VSS.n2859 VSS.n2457 4.5005
R26783 VSS.n3051 VSS.n2374 4.5005
R26784 VSS.n2374 VSS.n2351 4.5005
R26785 VSS.n2483 VSS.n2374 4.5005
R26786 VSS.n2484 VSS.n2374 4.5005
R26787 VSS.n2486 VSS.n2374 4.5005
R26788 VSS.n2489 VSS.n2374 4.5005
R26789 VSS.n2491 VSS.n2374 4.5005
R26790 VSS.n2492 VSS.n2374 4.5005
R26791 VSS.n2494 VSS.n2374 4.5005
R26792 VSS.n2497 VSS.n2374 4.5005
R26793 VSS.n2499 VSS.n2374 4.5005
R26794 VSS.n2500 VSS.n2374 4.5005
R26795 VSS.n2502 VSS.n2374 4.5005
R26796 VSS.n2505 VSS.n2374 4.5005
R26797 VSS.n2507 VSS.n2374 4.5005
R26798 VSS.n2508 VSS.n2374 4.5005
R26799 VSS.n2510 VSS.n2374 4.5005
R26800 VSS.n2513 VSS.n2374 4.5005
R26801 VSS.n2515 VSS.n2374 4.5005
R26802 VSS.n2516 VSS.n2374 4.5005
R26803 VSS.n2518 VSS.n2374 4.5005
R26804 VSS.n2521 VSS.n2374 4.5005
R26805 VSS.n2523 VSS.n2374 4.5005
R26806 VSS.n2524 VSS.n2374 4.5005
R26807 VSS.n2526 VSS.n2374 4.5005
R26808 VSS.n2529 VSS.n2374 4.5005
R26809 VSS.n2531 VSS.n2374 4.5005
R26810 VSS.n2532 VSS.n2374 4.5005
R26811 VSS.n2534 VSS.n2374 4.5005
R26812 VSS.n2537 VSS.n2374 4.5005
R26813 VSS.n2539 VSS.n2374 4.5005
R26814 VSS.n2540 VSS.n2374 4.5005
R26815 VSS.n2542 VSS.n2374 4.5005
R26816 VSS.n2545 VSS.n2374 4.5005
R26817 VSS.n2547 VSS.n2374 4.5005
R26818 VSS.n2548 VSS.n2374 4.5005
R26819 VSS.n2550 VSS.n2374 4.5005
R26820 VSS.n2553 VSS.n2374 4.5005
R26821 VSS.n2555 VSS.n2374 4.5005
R26822 VSS.n2556 VSS.n2374 4.5005
R26823 VSS.n2558 VSS.n2374 4.5005
R26824 VSS.n2561 VSS.n2374 4.5005
R26825 VSS.n2563 VSS.n2374 4.5005
R26826 VSS.n2564 VSS.n2374 4.5005
R26827 VSS.n2566 VSS.n2374 4.5005
R26828 VSS.n2569 VSS.n2374 4.5005
R26829 VSS.n2571 VSS.n2374 4.5005
R26830 VSS.n2572 VSS.n2374 4.5005
R26831 VSS.n2574 VSS.n2374 4.5005
R26832 VSS.n2577 VSS.n2374 4.5005
R26833 VSS.n2579 VSS.n2374 4.5005
R26834 VSS.n2580 VSS.n2374 4.5005
R26835 VSS.n2582 VSS.n2374 4.5005
R26836 VSS.n2585 VSS.n2374 4.5005
R26837 VSS.n2587 VSS.n2374 4.5005
R26838 VSS.n2588 VSS.n2374 4.5005
R26839 VSS.n2590 VSS.n2374 4.5005
R26840 VSS.n2593 VSS.n2374 4.5005
R26841 VSS.n2595 VSS.n2374 4.5005
R26842 VSS.n2596 VSS.n2374 4.5005
R26843 VSS.n2598 VSS.n2374 4.5005
R26844 VSS.n2601 VSS.n2374 4.5005
R26845 VSS.n2603 VSS.n2374 4.5005
R26846 VSS.n2604 VSS.n2374 4.5005
R26847 VSS.n2606 VSS.n2374 4.5005
R26848 VSS.n2609 VSS.n2374 4.5005
R26849 VSS.n2611 VSS.n2374 4.5005
R26850 VSS.n2612 VSS.n2374 4.5005
R26851 VSS.n2614 VSS.n2374 4.5005
R26852 VSS.n2617 VSS.n2374 4.5005
R26853 VSS.n2619 VSS.n2374 4.5005
R26854 VSS.n2620 VSS.n2374 4.5005
R26855 VSS.n2622 VSS.n2374 4.5005
R26856 VSS.n2625 VSS.n2374 4.5005
R26857 VSS.n2627 VSS.n2374 4.5005
R26858 VSS.n2628 VSS.n2374 4.5005
R26859 VSS.n2630 VSS.n2374 4.5005
R26860 VSS.n2633 VSS.n2374 4.5005
R26861 VSS.n2635 VSS.n2374 4.5005
R26862 VSS.n2636 VSS.n2374 4.5005
R26863 VSS.n2638 VSS.n2374 4.5005
R26864 VSS.n2640 VSS.n2374 4.5005
R26865 VSS.n2642 VSS.n2374 4.5005
R26866 VSS.n2643 VSS.n2374 4.5005
R26867 VSS.n2645 VSS.n2374 4.5005
R26868 VSS.n2648 VSS.n2374 4.5005
R26869 VSS.n2650 VSS.n2374 4.5005
R26870 VSS.n2651 VSS.n2374 4.5005
R26871 VSS.n2653 VSS.n2374 4.5005
R26872 VSS.n2656 VSS.n2374 4.5005
R26873 VSS.n2658 VSS.n2374 4.5005
R26874 VSS.n2659 VSS.n2374 4.5005
R26875 VSS.n2661 VSS.n2374 4.5005
R26876 VSS.n2664 VSS.n2374 4.5005
R26877 VSS.n2666 VSS.n2374 4.5005
R26878 VSS.n2667 VSS.n2374 4.5005
R26879 VSS.n2669 VSS.n2374 4.5005
R26880 VSS.n2672 VSS.n2374 4.5005
R26881 VSS.n2674 VSS.n2374 4.5005
R26882 VSS.n2675 VSS.n2374 4.5005
R26883 VSS.n2677 VSS.n2374 4.5005
R26884 VSS.n2680 VSS.n2374 4.5005
R26885 VSS.n2682 VSS.n2374 4.5005
R26886 VSS.n2683 VSS.n2374 4.5005
R26887 VSS.n2685 VSS.n2374 4.5005
R26888 VSS.n2688 VSS.n2374 4.5005
R26889 VSS.n2690 VSS.n2374 4.5005
R26890 VSS.n2691 VSS.n2374 4.5005
R26891 VSS.n2693 VSS.n2374 4.5005
R26892 VSS.n2696 VSS.n2374 4.5005
R26893 VSS.n2698 VSS.n2374 4.5005
R26894 VSS.n2699 VSS.n2374 4.5005
R26895 VSS.n2701 VSS.n2374 4.5005
R26896 VSS.n2704 VSS.n2374 4.5005
R26897 VSS.n2706 VSS.n2374 4.5005
R26898 VSS.n2707 VSS.n2374 4.5005
R26899 VSS.n2709 VSS.n2374 4.5005
R26900 VSS.n2712 VSS.n2374 4.5005
R26901 VSS.n2714 VSS.n2374 4.5005
R26902 VSS.n2715 VSS.n2374 4.5005
R26903 VSS.n2717 VSS.n2374 4.5005
R26904 VSS.n2720 VSS.n2374 4.5005
R26905 VSS.n2722 VSS.n2374 4.5005
R26906 VSS.n2723 VSS.n2374 4.5005
R26907 VSS.n2725 VSS.n2374 4.5005
R26908 VSS.n2793 VSS.n2374 4.5005
R26909 VSS.n2859 VSS.n2374 4.5005
R26910 VSS.n3051 VSS.n2458 4.5005
R26911 VSS.n2458 VSS.n2351 4.5005
R26912 VSS.n2483 VSS.n2458 4.5005
R26913 VSS.n2484 VSS.n2458 4.5005
R26914 VSS.n2486 VSS.n2458 4.5005
R26915 VSS.n2489 VSS.n2458 4.5005
R26916 VSS.n2491 VSS.n2458 4.5005
R26917 VSS.n2492 VSS.n2458 4.5005
R26918 VSS.n2494 VSS.n2458 4.5005
R26919 VSS.n2497 VSS.n2458 4.5005
R26920 VSS.n2499 VSS.n2458 4.5005
R26921 VSS.n2500 VSS.n2458 4.5005
R26922 VSS.n2502 VSS.n2458 4.5005
R26923 VSS.n2505 VSS.n2458 4.5005
R26924 VSS.n2507 VSS.n2458 4.5005
R26925 VSS.n2508 VSS.n2458 4.5005
R26926 VSS.n2510 VSS.n2458 4.5005
R26927 VSS.n2513 VSS.n2458 4.5005
R26928 VSS.n2515 VSS.n2458 4.5005
R26929 VSS.n2516 VSS.n2458 4.5005
R26930 VSS.n2518 VSS.n2458 4.5005
R26931 VSS.n2521 VSS.n2458 4.5005
R26932 VSS.n2523 VSS.n2458 4.5005
R26933 VSS.n2524 VSS.n2458 4.5005
R26934 VSS.n2526 VSS.n2458 4.5005
R26935 VSS.n2529 VSS.n2458 4.5005
R26936 VSS.n2531 VSS.n2458 4.5005
R26937 VSS.n2532 VSS.n2458 4.5005
R26938 VSS.n2534 VSS.n2458 4.5005
R26939 VSS.n2537 VSS.n2458 4.5005
R26940 VSS.n2539 VSS.n2458 4.5005
R26941 VSS.n2540 VSS.n2458 4.5005
R26942 VSS.n2542 VSS.n2458 4.5005
R26943 VSS.n2545 VSS.n2458 4.5005
R26944 VSS.n2547 VSS.n2458 4.5005
R26945 VSS.n2548 VSS.n2458 4.5005
R26946 VSS.n2550 VSS.n2458 4.5005
R26947 VSS.n2553 VSS.n2458 4.5005
R26948 VSS.n2555 VSS.n2458 4.5005
R26949 VSS.n2556 VSS.n2458 4.5005
R26950 VSS.n2558 VSS.n2458 4.5005
R26951 VSS.n2561 VSS.n2458 4.5005
R26952 VSS.n2563 VSS.n2458 4.5005
R26953 VSS.n2564 VSS.n2458 4.5005
R26954 VSS.n2566 VSS.n2458 4.5005
R26955 VSS.n2569 VSS.n2458 4.5005
R26956 VSS.n2571 VSS.n2458 4.5005
R26957 VSS.n2572 VSS.n2458 4.5005
R26958 VSS.n2574 VSS.n2458 4.5005
R26959 VSS.n2577 VSS.n2458 4.5005
R26960 VSS.n2579 VSS.n2458 4.5005
R26961 VSS.n2580 VSS.n2458 4.5005
R26962 VSS.n2582 VSS.n2458 4.5005
R26963 VSS.n2585 VSS.n2458 4.5005
R26964 VSS.n2587 VSS.n2458 4.5005
R26965 VSS.n2588 VSS.n2458 4.5005
R26966 VSS.n2590 VSS.n2458 4.5005
R26967 VSS.n2593 VSS.n2458 4.5005
R26968 VSS.n2595 VSS.n2458 4.5005
R26969 VSS.n2596 VSS.n2458 4.5005
R26970 VSS.n2598 VSS.n2458 4.5005
R26971 VSS.n2601 VSS.n2458 4.5005
R26972 VSS.n2603 VSS.n2458 4.5005
R26973 VSS.n2604 VSS.n2458 4.5005
R26974 VSS.n2606 VSS.n2458 4.5005
R26975 VSS.n2609 VSS.n2458 4.5005
R26976 VSS.n2611 VSS.n2458 4.5005
R26977 VSS.n2612 VSS.n2458 4.5005
R26978 VSS.n2614 VSS.n2458 4.5005
R26979 VSS.n2617 VSS.n2458 4.5005
R26980 VSS.n2619 VSS.n2458 4.5005
R26981 VSS.n2620 VSS.n2458 4.5005
R26982 VSS.n2622 VSS.n2458 4.5005
R26983 VSS.n2625 VSS.n2458 4.5005
R26984 VSS.n2627 VSS.n2458 4.5005
R26985 VSS.n2628 VSS.n2458 4.5005
R26986 VSS.n2630 VSS.n2458 4.5005
R26987 VSS.n2633 VSS.n2458 4.5005
R26988 VSS.n2635 VSS.n2458 4.5005
R26989 VSS.n2636 VSS.n2458 4.5005
R26990 VSS.n2638 VSS.n2458 4.5005
R26991 VSS.n2640 VSS.n2458 4.5005
R26992 VSS.n2642 VSS.n2458 4.5005
R26993 VSS.n2643 VSS.n2458 4.5005
R26994 VSS.n2645 VSS.n2458 4.5005
R26995 VSS.n2648 VSS.n2458 4.5005
R26996 VSS.n2650 VSS.n2458 4.5005
R26997 VSS.n2651 VSS.n2458 4.5005
R26998 VSS.n2653 VSS.n2458 4.5005
R26999 VSS.n2656 VSS.n2458 4.5005
R27000 VSS.n2658 VSS.n2458 4.5005
R27001 VSS.n2659 VSS.n2458 4.5005
R27002 VSS.n2661 VSS.n2458 4.5005
R27003 VSS.n2664 VSS.n2458 4.5005
R27004 VSS.n2666 VSS.n2458 4.5005
R27005 VSS.n2667 VSS.n2458 4.5005
R27006 VSS.n2669 VSS.n2458 4.5005
R27007 VSS.n2672 VSS.n2458 4.5005
R27008 VSS.n2674 VSS.n2458 4.5005
R27009 VSS.n2675 VSS.n2458 4.5005
R27010 VSS.n2677 VSS.n2458 4.5005
R27011 VSS.n2680 VSS.n2458 4.5005
R27012 VSS.n2682 VSS.n2458 4.5005
R27013 VSS.n2683 VSS.n2458 4.5005
R27014 VSS.n2685 VSS.n2458 4.5005
R27015 VSS.n2688 VSS.n2458 4.5005
R27016 VSS.n2690 VSS.n2458 4.5005
R27017 VSS.n2691 VSS.n2458 4.5005
R27018 VSS.n2693 VSS.n2458 4.5005
R27019 VSS.n2696 VSS.n2458 4.5005
R27020 VSS.n2698 VSS.n2458 4.5005
R27021 VSS.n2699 VSS.n2458 4.5005
R27022 VSS.n2701 VSS.n2458 4.5005
R27023 VSS.n2704 VSS.n2458 4.5005
R27024 VSS.n2706 VSS.n2458 4.5005
R27025 VSS.n2707 VSS.n2458 4.5005
R27026 VSS.n2709 VSS.n2458 4.5005
R27027 VSS.n2712 VSS.n2458 4.5005
R27028 VSS.n2714 VSS.n2458 4.5005
R27029 VSS.n2715 VSS.n2458 4.5005
R27030 VSS.n2717 VSS.n2458 4.5005
R27031 VSS.n2720 VSS.n2458 4.5005
R27032 VSS.n2722 VSS.n2458 4.5005
R27033 VSS.n2723 VSS.n2458 4.5005
R27034 VSS.n2725 VSS.n2458 4.5005
R27035 VSS.n2793 VSS.n2458 4.5005
R27036 VSS.n2859 VSS.n2458 4.5005
R27037 VSS.n3051 VSS.n2373 4.5005
R27038 VSS.n2373 VSS.n2351 4.5005
R27039 VSS.n2483 VSS.n2373 4.5005
R27040 VSS.n2484 VSS.n2373 4.5005
R27041 VSS.n2486 VSS.n2373 4.5005
R27042 VSS.n2489 VSS.n2373 4.5005
R27043 VSS.n2491 VSS.n2373 4.5005
R27044 VSS.n2492 VSS.n2373 4.5005
R27045 VSS.n2494 VSS.n2373 4.5005
R27046 VSS.n2497 VSS.n2373 4.5005
R27047 VSS.n2499 VSS.n2373 4.5005
R27048 VSS.n2500 VSS.n2373 4.5005
R27049 VSS.n2502 VSS.n2373 4.5005
R27050 VSS.n2505 VSS.n2373 4.5005
R27051 VSS.n2507 VSS.n2373 4.5005
R27052 VSS.n2508 VSS.n2373 4.5005
R27053 VSS.n2510 VSS.n2373 4.5005
R27054 VSS.n2513 VSS.n2373 4.5005
R27055 VSS.n2515 VSS.n2373 4.5005
R27056 VSS.n2516 VSS.n2373 4.5005
R27057 VSS.n2518 VSS.n2373 4.5005
R27058 VSS.n2521 VSS.n2373 4.5005
R27059 VSS.n2523 VSS.n2373 4.5005
R27060 VSS.n2524 VSS.n2373 4.5005
R27061 VSS.n2526 VSS.n2373 4.5005
R27062 VSS.n2529 VSS.n2373 4.5005
R27063 VSS.n2531 VSS.n2373 4.5005
R27064 VSS.n2532 VSS.n2373 4.5005
R27065 VSS.n2534 VSS.n2373 4.5005
R27066 VSS.n2537 VSS.n2373 4.5005
R27067 VSS.n2539 VSS.n2373 4.5005
R27068 VSS.n2540 VSS.n2373 4.5005
R27069 VSS.n2542 VSS.n2373 4.5005
R27070 VSS.n2545 VSS.n2373 4.5005
R27071 VSS.n2547 VSS.n2373 4.5005
R27072 VSS.n2548 VSS.n2373 4.5005
R27073 VSS.n2550 VSS.n2373 4.5005
R27074 VSS.n2553 VSS.n2373 4.5005
R27075 VSS.n2555 VSS.n2373 4.5005
R27076 VSS.n2556 VSS.n2373 4.5005
R27077 VSS.n2558 VSS.n2373 4.5005
R27078 VSS.n2561 VSS.n2373 4.5005
R27079 VSS.n2563 VSS.n2373 4.5005
R27080 VSS.n2564 VSS.n2373 4.5005
R27081 VSS.n2566 VSS.n2373 4.5005
R27082 VSS.n2569 VSS.n2373 4.5005
R27083 VSS.n2571 VSS.n2373 4.5005
R27084 VSS.n2572 VSS.n2373 4.5005
R27085 VSS.n2574 VSS.n2373 4.5005
R27086 VSS.n2577 VSS.n2373 4.5005
R27087 VSS.n2579 VSS.n2373 4.5005
R27088 VSS.n2580 VSS.n2373 4.5005
R27089 VSS.n2582 VSS.n2373 4.5005
R27090 VSS.n2585 VSS.n2373 4.5005
R27091 VSS.n2587 VSS.n2373 4.5005
R27092 VSS.n2588 VSS.n2373 4.5005
R27093 VSS.n2590 VSS.n2373 4.5005
R27094 VSS.n2593 VSS.n2373 4.5005
R27095 VSS.n2595 VSS.n2373 4.5005
R27096 VSS.n2596 VSS.n2373 4.5005
R27097 VSS.n2598 VSS.n2373 4.5005
R27098 VSS.n2601 VSS.n2373 4.5005
R27099 VSS.n2603 VSS.n2373 4.5005
R27100 VSS.n2604 VSS.n2373 4.5005
R27101 VSS.n2606 VSS.n2373 4.5005
R27102 VSS.n2609 VSS.n2373 4.5005
R27103 VSS.n2611 VSS.n2373 4.5005
R27104 VSS.n2612 VSS.n2373 4.5005
R27105 VSS.n2614 VSS.n2373 4.5005
R27106 VSS.n2617 VSS.n2373 4.5005
R27107 VSS.n2619 VSS.n2373 4.5005
R27108 VSS.n2620 VSS.n2373 4.5005
R27109 VSS.n2622 VSS.n2373 4.5005
R27110 VSS.n2625 VSS.n2373 4.5005
R27111 VSS.n2627 VSS.n2373 4.5005
R27112 VSS.n2628 VSS.n2373 4.5005
R27113 VSS.n2630 VSS.n2373 4.5005
R27114 VSS.n2633 VSS.n2373 4.5005
R27115 VSS.n2635 VSS.n2373 4.5005
R27116 VSS.n2636 VSS.n2373 4.5005
R27117 VSS.n2638 VSS.n2373 4.5005
R27118 VSS.n2640 VSS.n2373 4.5005
R27119 VSS.n2642 VSS.n2373 4.5005
R27120 VSS.n2643 VSS.n2373 4.5005
R27121 VSS.n2645 VSS.n2373 4.5005
R27122 VSS.n2648 VSS.n2373 4.5005
R27123 VSS.n2650 VSS.n2373 4.5005
R27124 VSS.n2651 VSS.n2373 4.5005
R27125 VSS.n2653 VSS.n2373 4.5005
R27126 VSS.n2656 VSS.n2373 4.5005
R27127 VSS.n2658 VSS.n2373 4.5005
R27128 VSS.n2659 VSS.n2373 4.5005
R27129 VSS.n2661 VSS.n2373 4.5005
R27130 VSS.n2664 VSS.n2373 4.5005
R27131 VSS.n2666 VSS.n2373 4.5005
R27132 VSS.n2667 VSS.n2373 4.5005
R27133 VSS.n2669 VSS.n2373 4.5005
R27134 VSS.n2672 VSS.n2373 4.5005
R27135 VSS.n2674 VSS.n2373 4.5005
R27136 VSS.n2675 VSS.n2373 4.5005
R27137 VSS.n2677 VSS.n2373 4.5005
R27138 VSS.n2680 VSS.n2373 4.5005
R27139 VSS.n2682 VSS.n2373 4.5005
R27140 VSS.n2683 VSS.n2373 4.5005
R27141 VSS.n2685 VSS.n2373 4.5005
R27142 VSS.n2688 VSS.n2373 4.5005
R27143 VSS.n2690 VSS.n2373 4.5005
R27144 VSS.n2691 VSS.n2373 4.5005
R27145 VSS.n2693 VSS.n2373 4.5005
R27146 VSS.n2696 VSS.n2373 4.5005
R27147 VSS.n2698 VSS.n2373 4.5005
R27148 VSS.n2699 VSS.n2373 4.5005
R27149 VSS.n2701 VSS.n2373 4.5005
R27150 VSS.n2704 VSS.n2373 4.5005
R27151 VSS.n2706 VSS.n2373 4.5005
R27152 VSS.n2707 VSS.n2373 4.5005
R27153 VSS.n2709 VSS.n2373 4.5005
R27154 VSS.n2712 VSS.n2373 4.5005
R27155 VSS.n2714 VSS.n2373 4.5005
R27156 VSS.n2715 VSS.n2373 4.5005
R27157 VSS.n2717 VSS.n2373 4.5005
R27158 VSS.n2720 VSS.n2373 4.5005
R27159 VSS.n2722 VSS.n2373 4.5005
R27160 VSS.n2723 VSS.n2373 4.5005
R27161 VSS.n2725 VSS.n2373 4.5005
R27162 VSS.n2793 VSS.n2373 4.5005
R27163 VSS.n2859 VSS.n2373 4.5005
R27164 VSS.n3051 VSS.n2459 4.5005
R27165 VSS.n2459 VSS.n2351 4.5005
R27166 VSS.n2483 VSS.n2459 4.5005
R27167 VSS.n2484 VSS.n2459 4.5005
R27168 VSS.n2486 VSS.n2459 4.5005
R27169 VSS.n2489 VSS.n2459 4.5005
R27170 VSS.n2491 VSS.n2459 4.5005
R27171 VSS.n2492 VSS.n2459 4.5005
R27172 VSS.n2494 VSS.n2459 4.5005
R27173 VSS.n2497 VSS.n2459 4.5005
R27174 VSS.n2499 VSS.n2459 4.5005
R27175 VSS.n2500 VSS.n2459 4.5005
R27176 VSS.n2502 VSS.n2459 4.5005
R27177 VSS.n2505 VSS.n2459 4.5005
R27178 VSS.n2507 VSS.n2459 4.5005
R27179 VSS.n2508 VSS.n2459 4.5005
R27180 VSS.n2510 VSS.n2459 4.5005
R27181 VSS.n2513 VSS.n2459 4.5005
R27182 VSS.n2515 VSS.n2459 4.5005
R27183 VSS.n2516 VSS.n2459 4.5005
R27184 VSS.n2518 VSS.n2459 4.5005
R27185 VSS.n2521 VSS.n2459 4.5005
R27186 VSS.n2523 VSS.n2459 4.5005
R27187 VSS.n2524 VSS.n2459 4.5005
R27188 VSS.n2526 VSS.n2459 4.5005
R27189 VSS.n2529 VSS.n2459 4.5005
R27190 VSS.n2531 VSS.n2459 4.5005
R27191 VSS.n2532 VSS.n2459 4.5005
R27192 VSS.n2534 VSS.n2459 4.5005
R27193 VSS.n2537 VSS.n2459 4.5005
R27194 VSS.n2539 VSS.n2459 4.5005
R27195 VSS.n2540 VSS.n2459 4.5005
R27196 VSS.n2542 VSS.n2459 4.5005
R27197 VSS.n2545 VSS.n2459 4.5005
R27198 VSS.n2547 VSS.n2459 4.5005
R27199 VSS.n2548 VSS.n2459 4.5005
R27200 VSS.n2550 VSS.n2459 4.5005
R27201 VSS.n2553 VSS.n2459 4.5005
R27202 VSS.n2555 VSS.n2459 4.5005
R27203 VSS.n2556 VSS.n2459 4.5005
R27204 VSS.n2558 VSS.n2459 4.5005
R27205 VSS.n2561 VSS.n2459 4.5005
R27206 VSS.n2563 VSS.n2459 4.5005
R27207 VSS.n2564 VSS.n2459 4.5005
R27208 VSS.n2566 VSS.n2459 4.5005
R27209 VSS.n2569 VSS.n2459 4.5005
R27210 VSS.n2571 VSS.n2459 4.5005
R27211 VSS.n2572 VSS.n2459 4.5005
R27212 VSS.n2574 VSS.n2459 4.5005
R27213 VSS.n2577 VSS.n2459 4.5005
R27214 VSS.n2579 VSS.n2459 4.5005
R27215 VSS.n2580 VSS.n2459 4.5005
R27216 VSS.n2582 VSS.n2459 4.5005
R27217 VSS.n2585 VSS.n2459 4.5005
R27218 VSS.n2587 VSS.n2459 4.5005
R27219 VSS.n2588 VSS.n2459 4.5005
R27220 VSS.n2590 VSS.n2459 4.5005
R27221 VSS.n2593 VSS.n2459 4.5005
R27222 VSS.n2595 VSS.n2459 4.5005
R27223 VSS.n2596 VSS.n2459 4.5005
R27224 VSS.n2598 VSS.n2459 4.5005
R27225 VSS.n2601 VSS.n2459 4.5005
R27226 VSS.n2603 VSS.n2459 4.5005
R27227 VSS.n2604 VSS.n2459 4.5005
R27228 VSS.n2606 VSS.n2459 4.5005
R27229 VSS.n2609 VSS.n2459 4.5005
R27230 VSS.n2611 VSS.n2459 4.5005
R27231 VSS.n2612 VSS.n2459 4.5005
R27232 VSS.n2614 VSS.n2459 4.5005
R27233 VSS.n2617 VSS.n2459 4.5005
R27234 VSS.n2619 VSS.n2459 4.5005
R27235 VSS.n2620 VSS.n2459 4.5005
R27236 VSS.n2622 VSS.n2459 4.5005
R27237 VSS.n2625 VSS.n2459 4.5005
R27238 VSS.n2627 VSS.n2459 4.5005
R27239 VSS.n2628 VSS.n2459 4.5005
R27240 VSS.n2630 VSS.n2459 4.5005
R27241 VSS.n2633 VSS.n2459 4.5005
R27242 VSS.n2635 VSS.n2459 4.5005
R27243 VSS.n2636 VSS.n2459 4.5005
R27244 VSS.n2638 VSS.n2459 4.5005
R27245 VSS.n2640 VSS.n2459 4.5005
R27246 VSS.n2642 VSS.n2459 4.5005
R27247 VSS.n2643 VSS.n2459 4.5005
R27248 VSS.n2645 VSS.n2459 4.5005
R27249 VSS.n2648 VSS.n2459 4.5005
R27250 VSS.n2650 VSS.n2459 4.5005
R27251 VSS.n2651 VSS.n2459 4.5005
R27252 VSS.n2653 VSS.n2459 4.5005
R27253 VSS.n2656 VSS.n2459 4.5005
R27254 VSS.n2658 VSS.n2459 4.5005
R27255 VSS.n2659 VSS.n2459 4.5005
R27256 VSS.n2661 VSS.n2459 4.5005
R27257 VSS.n2664 VSS.n2459 4.5005
R27258 VSS.n2666 VSS.n2459 4.5005
R27259 VSS.n2667 VSS.n2459 4.5005
R27260 VSS.n2669 VSS.n2459 4.5005
R27261 VSS.n2672 VSS.n2459 4.5005
R27262 VSS.n2674 VSS.n2459 4.5005
R27263 VSS.n2675 VSS.n2459 4.5005
R27264 VSS.n2677 VSS.n2459 4.5005
R27265 VSS.n2680 VSS.n2459 4.5005
R27266 VSS.n2682 VSS.n2459 4.5005
R27267 VSS.n2683 VSS.n2459 4.5005
R27268 VSS.n2685 VSS.n2459 4.5005
R27269 VSS.n2688 VSS.n2459 4.5005
R27270 VSS.n2690 VSS.n2459 4.5005
R27271 VSS.n2691 VSS.n2459 4.5005
R27272 VSS.n2693 VSS.n2459 4.5005
R27273 VSS.n2696 VSS.n2459 4.5005
R27274 VSS.n2698 VSS.n2459 4.5005
R27275 VSS.n2699 VSS.n2459 4.5005
R27276 VSS.n2701 VSS.n2459 4.5005
R27277 VSS.n2704 VSS.n2459 4.5005
R27278 VSS.n2706 VSS.n2459 4.5005
R27279 VSS.n2707 VSS.n2459 4.5005
R27280 VSS.n2709 VSS.n2459 4.5005
R27281 VSS.n2712 VSS.n2459 4.5005
R27282 VSS.n2714 VSS.n2459 4.5005
R27283 VSS.n2715 VSS.n2459 4.5005
R27284 VSS.n2717 VSS.n2459 4.5005
R27285 VSS.n2720 VSS.n2459 4.5005
R27286 VSS.n2722 VSS.n2459 4.5005
R27287 VSS.n2723 VSS.n2459 4.5005
R27288 VSS.n2725 VSS.n2459 4.5005
R27289 VSS.n2793 VSS.n2459 4.5005
R27290 VSS.n2859 VSS.n2459 4.5005
R27291 VSS.n3051 VSS.n2372 4.5005
R27292 VSS.n2372 VSS.n2351 4.5005
R27293 VSS.n2483 VSS.n2372 4.5005
R27294 VSS.n2484 VSS.n2372 4.5005
R27295 VSS.n2486 VSS.n2372 4.5005
R27296 VSS.n2489 VSS.n2372 4.5005
R27297 VSS.n2491 VSS.n2372 4.5005
R27298 VSS.n2492 VSS.n2372 4.5005
R27299 VSS.n2494 VSS.n2372 4.5005
R27300 VSS.n2497 VSS.n2372 4.5005
R27301 VSS.n2499 VSS.n2372 4.5005
R27302 VSS.n2500 VSS.n2372 4.5005
R27303 VSS.n2502 VSS.n2372 4.5005
R27304 VSS.n2505 VSS.n2372 4.5005
R27305 VSS.n2507 VSS.n2372 4.5005
R27306 VSS.n2508 VSS.n2372 4.5005
R27307 VSS.n2510 VSS.n2372 4.5005
R27308 VSS.n2513 VSS.n2372 4.5005
R27309 VSS.n2515 VSS.n2372 4.5005
R27310 VSS.n2516 VSS.n2372 4.5005
R27311 VSS.n2518 VSS.n2372 4.5005
R27312 VSS.n2521 VSS.n2372 4.5005
R27313 VSS.n2523 VSS.n2372 4.5005
R27314 VSS.n2524 VSS.n2372 4.5005
R27315 VSS.n2526 VSS.n2372 4.5005
R27316 VSS.n2529 VSS.n2372 4.5005
R27317 VSS.n2531 VSS.n2372 4.5005
R27318 VSS.n2532 VSS.n2372 4.5005
R27319 VSS.n2534 VSS.n2372 4.5005
R27320 VSS.n2537 VSS.n2372 4.5005
R27321 VSS.n2539 VSS.n2372 4.5005
R27322 VSS.n2540 VSS.n2372 4.5005
R27323 VSS.n2542 VSS.n2372 4.5005
R27324 VSS.n2545 VSS.n2372 4.5005
R27325 VSS.n2547 VSS.n2372 4.5005
R27326 VSS.n2548 VSS.n2372 4.5005
R27327 VSS.n2550 VSS.n2372 4.5005
R27328 VSS.n2553 VSS.n2372 4.5005
R27329 VSS.n2555 VSS.n2372 4.5005
R27330 VSS.n2556 VSS.n2372 4.5005
R27331 VSS.n2558 VSS.n2372 4.5005
R27332 VSS.n2561 VSS.n2372 4.5005
R27333 VSS.n2563 VSS.n2372 4.5005
R27334 VSS.n2564 VSS.n2372 4.5005
R27335 VSS.n2566 VSS.n2372 4.5005
R27336 VSS.n2569 VSS.n2372 4.5005
R27337 VSS.n2571 VSS.n2372 4.5005
R27338 VSS.n2572 VSS.n2372 4.5005
R27339 VSS.n2574 VSS.n2372 4.5005
R27340 VSS.n2577 VSS.n2372 4.5005
R27341 VSS.n2579 VSS.n2372 4.5005
R27342 VSS.n2580 VSS.n2372 4.5005
R27343 VSS.n2582 VSS.n2372 4.5005
R27344 VSS.n2585 VSS.n2372 4.5005
R27345 VSS.n2587 VSS.n2372 4.5005
R27346 VSS.n2588 VSS.n2372 4.5005
R27347 VSS.n2590 VSS.n2372 4.5005
R27348 VSS.n2593 VSS.n2372 4.5005
R27349 VSS.n2595 VSS.n2372 4.5005
R27350 VSS.n2596 VSS.n2372 4.5005
R27351 VSS.n2598 VSS.n2372 4.5005
R27352 VSS.n2601 VSS.n2372 4.5005
R27353 VSS.n2603 VSS.n2372 4.5005
R27354 VSS.n2604 VSS.n2372 4.5005
R27355 VSS.n2606 VSS.n2372 4.5005
R27356 VSS.n2609 VSS.n2372 4.5005
R27357 VSS.n2611 VSS.n2372 4.5005
R27358 VSS.n2612 VSS.n2372 4.5005
R27359 VSS.n2614 VSS.n2372 4.5005
R27360 VSS.n2617 VSS.n2372 4.5005
R27361 VSS.n2619 VSS.n2372 4.5005
R27362 VSS.n2620 VSS.n2372 4.5005
R27363 VSS.n2622 VSS.n2372 4.5005
R27364 VSS.n2625 VSS.n2372 4.5005
R27365 VSS.n2627 VSS.n2372 4.5005
R27366 VSS.n2628 VSS.n2372 4.5005
R27367 VSS.n2630 VSS.n2372 4.5005
R27368 VSS.n2633 VSS.n2372 4.5005
R27369 VSS.n2635 VSS.n2372 4.5005
R27370 VSS.n2636 VSS.n2372 4.5005
R27371 VSS.n2638 VSS.n2372 4.5005
R27372 VSS.n2640 VSS.n2372 4.5005
R27373 VSS.n2642 VSS.n2372 4.5005
R27374 VSS.n2643 VSS.n2372 4.5005
R27375 VSS.n2645 VSS.n2372 4.5005
R27376 VSS.n2648 VSS.n2372 4.5005
R27377 VSS.n2650 VSS.n2372 4.5005
R27378 VSS.n2651 VSS.n2372 4.5005
R27379 VSS.n2653 VSS.n2372 4.5005
R27380 VSS.n2656 VSS.n2372 4.5005
R27381 VSS.n2658 VSS.n2372 4.5005
R27382 VSS.n2659 VSS.n2372 4.5005
R27383 VSS.n2661 VSS.n2372 4.5005
R27384 VSS.n2664 VSS.n2372 4.5005
R27385 VSS.n2666 VSS.n2372 4.5005
R27386 VSS.n2667 VSS.n2372 4.5005
R27387 VSS.n2669 VSS.n2372 4.5005
R27388 VSS.n2672 VSS.n2372 4.5005
R27389 VSS.n2674 VSS.n2372 4.5005
R27390 VSS.n2675 VSS.n2372 4.5005
R27391 VSS.n2677 VSS.n2372 4.5005
R27392 VSS.n2680 VSS.n2372 4.5005
R27393 VSS.n2682 VSS.n2372 4.5005
R27394 VSS.n2683 VSS.n2372 4.5005
R27395 VSS.n2685 VSS.n2372 4.5005
R27396 VSS.n2688 VSS.n2372 4.5005
R27397 VSS.n2690 VSS.n2372 4.5005
R27398 VSS.n2691 VSS.n2372 4.5005
R27399 VSS.n2693 VSS.n2372 4.5005
R27400 VSS.n2696 VSS.n2372 4.5005
R27401 VSS.n2698 VSS.n2372 4.5005
R27402 VSS.n2699 VSS.n2372 4.5005
R27403 VSS.n2701 VSS.n2372 4.5005
R27404 VSS.n2704 VSS.n2372 4.5005
R27405 VSS.n2706 VSS.n2372 4.5005
R27406 VSS.n2707 VSS.n2372 4.5005
R27407 VSS.n2709 VSS.n2372 4.5005
R27408 VSS.n2712 VSS.n2372 4.5005
R27409 VSS.n2714 VSS.n2372 4.5005
R27410 VSS.n2715 VSS.n2372 4.5005
R27411 VSS.n2717 VSS.n2372 4.5005
R27412 VSS.n2720 VSS.n2372 4.5005
R27413 VSS.n2722 VSS.n2372 4.5005
R27414 VSS.n2723 VSS.n2372 4.5005
R27415 VSS.n2725 VSS.n2372 4.5005
R27416 VSS.n2793 VSS.n2372 4.5005
R27417 VSS.n2859 VSS.n2372 4.5005
R27418 VSS.n3051 VSS.n2460 4.5005
R27419 VSS.n2460 VSS.n2351 4.5005
R27420 VSS.n2483 VSS.n2460 4.5005
R27421 VSS.n2484 VSS.n2460 4.5005
R27422 VSS.n2486 VSS.n2460 4.5005
R27423 VSS.n2489 VSS.n2460 4.5005
R27424 VSS.n2491 VSS.n2460 4.5005
R27425 VSS.n2492 VSS.n2460 4.5005
R27426 VSS.n2494 VSS.n2460 4.5005
R27427 VSS.n2497 VSS.n2460 4.5005
R27428 VSS.n2499 VSS.n2460 4.5005
R27429 VSS.n2500 VSS.n2460 4.5005
R27430 VSS.n2502 VSS.n2460 4.5005
R27431 VSS.n2505 VSS.n2460 4.5005
R27432 VSS.n2507 VSS.n2460 4.5005
R27433 VSS.n2508 VSS.n2460 4.5005
R27434 VSS.n2510 VSS.n2460 4.5005
R27435 VSS.n2513 VSS.n2460 4.5005
R27436 VSS.n2515 VSS.n2460 4.5005
R27437 VSS.n2516 VSS.n2460 4.5005
R27438 VSS.n2518 VSS.n2460 4.5005
R27439 VSS.n2521 VSS.n2460 4.5005
R27440 VSS.n2523 VSS.n2460 4.5005
R27441 VSS.n2524 VSS.n2460 4.5005
R27442 VSS.n2526 VSS.n2460 4.5005
R27443 VSS.n2529 VSS.n2460 4.5005
R27444 VSS.n2531 VSS.n2460 4.5005
R27445 VSS.n2532 VSS.n2460 4.5005
R27446 VSS.n2534 VSS.n2460 4.5005
R27447 VSS.n2537 VSS.n2460 4.5005
R27448 VSS.n2539 VSS.n2460 4.5005
R27449 VSS.n2540 VSS.n2460 4.5005
R27450 VSS.n2542 VSS.n2460 4.5005
R27451 VSS.n2545 VSS.n2460 4.5005
R27452 VSS.n2547 VSS.n2460 4.5005
R27453 VSS.n2548 VSS.n2460 4.5005
R27454 VSS.n2550 VSS.n2460 4.5005
R27455 VSS.n2553 VSS.n2460 4.5005
R27456 VSS.n2555 VSS.n2460 4.5005
R27457 VSS.n2556 VSS.n2460 4.5005
R27458 VSS.n2558 VSS.n2460 4.5005
R27459 VSS.n2561 VSS.n2460 4.5005
R27460 VSS.n2563 VSS.n2460 4.5005
R27461 VSS.n2564 VSS.n2460 4.5005
R27462 VSS.n2566 VSS.n2460 4.5005
R27463 VSS.n2569 VSS.n2460 4.5005
R27464 VSS.n2571 VSS.n2460 4.5005
R27465 VSS.n2572 VSS.n2460 4.5005
R27466 VSS.n2574 VSS.n2460 4.5005
R27467 VSS.n2577 VSS.n2460 4.5005
R27468 VSS.n2579 VSS.n2460 4.5005
R27469 VSS.n2580 VSS.n2460 4.5005
R27470 VSS.n2582 VSS.n2460 4.5005
R27471 VSS.n2585 VSS.n2460 4.5005
R27472 VSS.n2587 VSS.n2460 4.5005
R27473 VSS.n2588 VSS.n2460 4.5005
R27474 VSS.n2590 VSS.n2460 4.5005
R27475 VSS.n2593 VSS.n2460 4.5005
R27476 VSS.n2595 VSS.n2460 4.5005
R27477 VSS.n2596 VSS.n2460 4.5005
R27478 VSS.n2598 VSS.n2460 4.5005
R27479 VSS.n2601 VSS.n2460 4.5005
R27480 VSS.n2603 VSS.n2460 4.5005
R27481 VSS.n2604 VSS.n2460 4.5005
R27482 VSS.n2606 VSS.n2460 4.5005
R27483 VSS.n2609 VSS.n2460 4.5005
R27484 VSS.n2611 VSS.n2460 4.5005
R27485 VSS.n2612 VSS.n2460 4.5005
R27486 VSS.n2614 VSS.n2460 4.5005
R27487 VSS.n2617 VSS.n2460 4.5005
R27488 VSS.n2619 VSS.n2460 4.5005
R27489 VSS.n2620 VSS.n2460 4.5005
R27490 VSS.n2622 VSS.n2460 4.5005
R27491 VSS.n2625 VSS.n2460 4.5005
R27492 VSS.n2627 VSS.n2460 4.5005
R27493 VSS.n2628 VSS.n2460 4.5005
R27494 VSS.n2630 VSS.n2460 4.5005
R27495 VSS.n2633 VSS.n2460 4.5005
R27496 VSS.n2635 VSS.n2460 4.5005
R27497 VSS.n2636 VSS.n2460 4.5005
R27498 VSS.n2638 VSS.n2460 4.5005
R27499 VSS.n2640 VSS.n2460 4.5005
R27500 VSS.n2642 VSS.n2460 4.5005
R27501 VSS.n2643 VSS.n2460 4.5005
R27502 VSS.n2645 VSS.n2460 4.5005
R27503 VSS.n2648 VSS.n2460 4.5005
R27504 VSS.n2650 VSS.n2460 4.5005
R27505 VSS.n2651 VSS.n2460 4.5005
R27506 VSS.n2653 VSS.n2460 4.5005
R27507 VSS.n2656 VSS.n2460 4.5005
R27508 VSS.n2658 VSS.n2460 4.5005
R27509 VSS.n2659 VSS.n2460 4.5005
R27510 VSS.n2661 VSS.n2460 4.5005
R27511 VSS.n2664 VSS.n2460 4.5005
R27512 VSS.n2666 VSS.n2460 4.5005
R27513 VSS.n2667 VSS.n2460 4.5005
R27514 VSS.n2669 VSS.n2460 4.5005
R27515 VSS.n2672 VSS.n2460 4.5005
R27516 VSS.n2674 VSS.n2460 4.5005
R27517 VSS.n2675 VSS.n2460 4.5005
R27518 VSS.n2677 VSS.n2460 4.5005
R27519 VSS.n2680 VSS.n2460 4.5005
R27520 VSS.n2682 VSS.n2460 4.5005
R27521 VSS.n2683 VSS.n2460 4.5005
R27522 VSS.n2685 VSS.n2460 4.5005
R27523 VSS.n2688 VSS.n2460 4.5005
R27524 VSS.n2690 VSS.n2460 4.5005
R27525 VSS.n2691 VSS.n2460 4.5005
R27526 VSS.n2693 VSS.n2460 4.5005
R27527 VSS.n2696 VSS.n2460 4.5005
R27528 VSS.n2698 VSS.n2460 4.5005
R27529 VSS.n2699 VSS.n2460 4.5005
R27530 VSS.n2701 VSS.n2460 4.5005
R27531 VSS.n2704 VSS.n2460 4.5005
R27532 VSS.n2706 VSS.n2460 4.5005
R27533 VSS.n2707 VSS.n2460 4.5005
R27534 VSS.n2709 VSS.n2460 4.5005
R27535 VSS.n2712 VSS.n2460 4.5005
R27536 VSS.n2714 VSS.n2460 4.5005
R27537 VSS.n2715 VSS.n2460 4.5005
R27538 VSS.n2717 VSS.n2460 4.5005
R27539 VSS.n2720 VSS.n2460 4.5005
R27540 VSS.n2722 VSS.n2460 4.5005
R27541 VSS.n2723 VSS.n2460 4.5005
R27542 VSS.n2725 VSS.n2460 4.5005
R27543 VSS.n2793 VSS.n2460 4.5005
R27544 VSS.n2859 VSS.n2460 4.5005
R27545 VSS.n3051 VSS.n2371 4.5005
R27546 VSS.n2371 VSS.n2351 4.5005
R27547 VSS.n2483 VSS.n2371 4.5005
R27548 VSS.n2484 VSS.n2371 4.5005
R27549 VSS.n2486 VSS.n2371 4.5005
R27550 VSS.n2489 VSS.n2371 4.5005
R27551 VSS.n2491 VSS.n2371 4.5005
R27552 VSS.n2492 VSS.n2371 4.5005
R27553 VSS.n2494 VSS.n2371 4.5005
R27554 VSS.n2497 VSS.n2371 4.5005
R27555 VSS.n2499 VSS.n2371 4.5005
R27556 VSS.n2500 VSS.n2371 4.5005
R27557 VSS.n2502 VSS.n2371 4.5005
R27558 VSS.n2505 VSS.n2371 4.5005
R27559 VSS.n2507 VSS.n2371 4.5005
R27560 VSS.n2508 VSS.n2371 4.5005
R27561 VSS.n2510 VSS.n2371 4.5005
R27562 VSS.n2513 VSS.n2371 4.5005
R27563 VSS.n2515 VSS.n2371 4.5005
R27564 VSS.n2516 VSS.n2371 4.5005
R27565 VSS.n2518 VSS.n2371 4.5005
R27566 VSS.n2521 VSS.n2371 4.5005
R27567 VSS.n2523 VSS.n2371 4.5005
R27568 VSS.n2524 VSS.n2371 4.5005
R27569 VSS.n2526 VSS.n2371 4.5005
R27570 VSS.n2529 VSS.n2371 4.5005
R27571 VSS.n2531 VSS.n2371 4.5005
R27572 VSS.n2532 VSS.n2371 4.5005
R27573 VSS.n2534 VSS.n2371 4.5005
R27574 VSS.n2537 VSS.n2371 4.5005
R27575 VSS.n2539 VSS.n2371 4.5005
R27576 VSS.n2540 VSS.n2371 4.5005
R27577 VSS.n2542 VSS.n2371 4.5005
R27578 VSS.n2545 VSS.n2371 4.5005
R27579 VSS.n2547 VSS.n2371 4.5005
R27580 VSS.n2548 VSS.n2371 4.5005
R27581 VSS.n2550 VSS.n2371 4.5005
R27582 VSS.n2553 VSS.n2371 4.5005
R27583 VSS.n2555 VSS.n2371 4.5005
R27584 VSS.n2556 VSS.n2371 4.5005
R27585 VSS.n2558 VSS.n2371 4.5005
R27586 VSS.n2561 VSS.n2371 4.5005
R27587 VSS.n2563 VSS.n2371 4.5005
R27588 VSS.n2564 VSS.n2371 4.5005
R27589 VSS.n2566 VSS.n2371 4.5005
R27590 VSS.n2569 VSS.n2371 4.5005
R27591 VSS.n2571 VSS.n2371 4.5005
R27592 VSS.n2572 VSS.n2371 4.5005
R27593 VSS.n2574 VSS.n2371 4.5005
R27594 VSS.n2577 VSS.n2371 4.5005
R27595 VSS.n2579 VSS.n2371 4.5005
R27596 VSS.n2580 VSS.n2371 4.5005
R27597 VSS.n2582 VSS.n2371 4.5005
R27598 VSS.n2585 VSS.n2371 4.5005
R27599 VSS.n2587 VSS.n2371 4.5005
R27600 VSS.n2588 VSS.n2371 4.5005
R27601 VSS.n2590 VSS.n2371 4.5005
R27602 VSS.n2593 VSS.n2371 4.5005
R27603 VSS.n2595 VSS.n2371 4.5005
R27604 VSS.n2596 VSS.n2371 4.5005
R27605 VSS.n2598 VSS.n2371 4.5005
R27606 VSS.n2601 VSS.n2371 4.5005
R27607 VSS.n2603 VSS.n2371 4.5005
R27608 VSS.n2604 VSS.n2371 4.5005
R27609 VSS.n2606 VSS.n2371 4.5005
R27610 VSS.n2609 VSS.n2371 4.5005
R27611 VSS.n2611 VSS.n2371 4.5005
R27612 VSS.n2612 VSS.n2371 4.5005
R27613 VSS.n2614 VSS.n2371 4.5005
R27614 VSS.n2617 VSS.n2371 4.5005
R27615 VSS.n2619 VSS.n2371 4.5005
R27616 VSS.n2620 VSS.n2371 4.5005
R27617 VSS.n2622 VSS.n2371 4.5005
R27618 VSS.n2625 VSS.n2371 4.5005
R27619 VSS.n2627 VSS.n2371 4.5005
R27620 VSS.n2628 VSS.n2371 4.5005
R27621 VSS.n2630 VSS.n2371 4.5005
R27622 VSS.n2633 VSS.n2371 4.5005
R27623 VSS.n2635 VSS.n2371 4.5005
R27624 VSS.n2636 VSS.n2371 4.5005
R27625 VSS.n2638 VSS.n2371 4.5005
R27626 VSS.n2640 VSS.n2371 4.5005
R27627 VSS.n2642 VSS.n2371 4.5005
R27628 VSS.n2643 VSS.n2371 4.5005
R27629 VSS.n2645 VSS.n2371 4.5005
R27630 VSS.n2648 VSS.n2371 4.5005
R27631 VSS.n2650 VSS.n2371 4.5005
R27632 VSS.n2651 VSS.n2371 4.5005
R27633 VSS.n2653 VSS.n2371 4.5005
R27634 VSS.n2656 VSS.n2371 4.5005
R27635 VSS.n2658 VSS.n2371 4.5005
R27636 VSS.n2659 VSS.n2371 4.5005
R27637 VSS.n2661 VSS.n2371 4.5005
R27638 VSS.n2664 VSS.n2371 4.5005
R27639 VSS.n2666 VSS.n2371 4.5005
R27640 VSS.n2667 VSS.n2371 4.5005
R27641 VSS.n2669 VSS.n2371 4.5005
R27642 VSS.n2672 VSS.n2371 4.5005
R27643 VSS.n2674 VSS.n2371 4.5005
R27644 VSS.n2675 VSS.n2371 4.5005
R27645 VSS.n2677 VSS.n2371 4.5005
R27646 VSS.n2680 VSS.n2371 4.5005
R27647 VSS.n2682 VSS.n2371 4.5005
R27648 VSS.n2683 VSS.n2371 4.5005
R27649 VSS.n2685 VSS.n2371 4.5005
R27650 VSS.n2688 VSS.n2371 4.5005
R27651 VSS.n2690 VSS.n2371 4.5005
R27652 VSS.n2691 VSS.n2371 4.5005
R27653 VSS.n2693 VSS.n2371 4.5005
R27654 VSS.n2696 VSS.n2371 4.5005
R27655 VSS.n2698 VSS.n2371 4.5005
R27656 VSS.n2699 VSS.n2371 4.5005
R27657 VSS.n2701 VSS.n2371 4.5005
R27658 VSS.n2704 VSS.n2371 4.5005
R27659 VSS.n2706 VSS.n2371 4.5005
R27660 VSS.n2707 VSS.n2371 4.5005
R27661 VSS.n2709 VSS.n2371 4.5005
R27662 VSS.n2712 VSS.n2371 4.5005
R27663 VSS.n2714 VSS.n2371 4.5005
R27664 VSS.n2715 VSS.n2371 4.5005
R27665 VSS.n2717 VSS.n2371 4.5005
R27666 VSS.n2720 VSS.n2371 4.5005
R27667 VSS.n2722 VSS.n2371 4.5005
R27668 VSS.n2723 VSS.n2371 4.5005
R27669 VSS.n2725 VSS.n2371 4.5005
R27670 VSS.n2793 VSS.n2371 4.5005
R27671 VSS.n2859 VSS.n2371 4.5005
R27672 VSS.n3051 VSS.n2461 4.5005
R27673 VSS.n2461 VSS.n2351 4.5005
R27674 VSS.n2483 VSS.n2461 4.5005
R27675 VSS.n2484 VSS.n2461 4.5005
R27676 VSS.n2486 VSS.n2461 4.5005
R27677 VSS.n2489 VSS.n2461 4.5005
R27678 VSS.n2491 VSS.n2461 4.5005
R27679 VSS.n2492 VSS.n2461 4.5005
R27680 VSS.n2494 VSS.n2461 4.5005
R27681 VSS.n2497 VSS.n2461 4.5005
R27682 VSS.n2499 VSS.n2461 4.5005
R27683 VSS.n2500 VSS.n2461 4.5005
R27684 VSS.n2502 VSS.n2461 4.5005
R27685 VSS.n2505 VSS.n2461 4.5005
R27686 VSS.n2507 VSS.n2461 4.5005
R27687 VSS.n2508 VSS.n2461 4.5005
R27688 VSS.n2510 VSS.n2461 4.5005
R27689 VSS.n2513 VSS.n2461 4.5005
R27690 VSS.n2515 VSS.n2461 4.5005
R27691 VSS.n2516 VSS.n2461 4.5005
R27692 VSS.n2518 VSS.n2461 4.5005
R27693 VSS.n2521 VSS.n2461 4.5005
R27694 VSS.n2523 VSS.n2461 4.5005
R27695 VSS.n2524 VSS.n2461 4.5005
R27696 VSS.n2526 VSS.n2461 4.5005
R27697 VSS.n2529 VSS.n2461 4.5005
R27698 VSS.n2531 VSS.n2461 4.5005
R27699 VSS.n2532 VSS.n2461 4.5005
R27700 VSS.n2534 VSS.n2461 4.5005
R27701 VSS.n2537 VSS.n2461 4.5005
R27702 VSS.n2539 VSS.n2461 4.5005
R27703 VSS.n2540 VSS.n2461 4.5005
R27704 VSS.n2542 VSS.n2461 4.5005
R27705 VSS.n2545 VSS.n2461 4.5005
R27706 VSS.n2547 VSS.n2461 4.5005
R27707 VSS.n2548 VSS.n2461 4.5005
R27708 VSS.n2550 VSS.n2461 4.5005
R27709 VSS.n2553 VSS.n2461 4.5005
R27710 VSS.n2555 VSS.n2461 4.5005
R27711 VSS.n2556 VSS.n2461 4.5005
R27712 VSS.n2558 VSS.n2461 4.5005
R27713 VSS.n2561 VSS.n2461 4.5005
R27714 VSS.n2563 VSS.n2461 4.5005
R27715 VSS.n2564 VSS.n2461 4.5005
R27716 VSS.n2566 VSS.n2461 4.5005
R27717 VSS.n2569 VSS.n2461 4.5005
R27718 VSS.n2571 VSS.n2461 4.5005
R27719 VSS.n2572 VSS.n2461 4.5005
R27720 VSS.n2574 VSS.n2461 4.5005
R27721 VSS.n2577 VSS.n2461 4.5005
R27722 VSS.n2579 VSS.n2461 4.5005
R27723 VSS.n2580 VSS.n2461 4.5005
R27724 VSS.n2582 VSS.n2461 4.5005
R27725 VSS.n2585 VSS.n2461 4.5005
R27726 VSS.n2587 VSS.n2461 4.5005
R27727 VSS.n2588 VSS.n2461 4.5005
R27728 VSS.n2590 VSS.n2461 4.5005
R27729 VSS.n2593 VSS.n2461 4.5005
R27730 VSS.n2595 VSS.n2461 4.5005
R27731 VSS.n2596 VSS.n2461 4.5005
R27732 VSS.n2598 VSS.n2461 4.5005
R27733 VSS.n2601 VSS.n2461 4.5005
R27734 VSS.n2603 VSS.n2461 4.5005
R27735 VSS.n2604 VSS.n2461 4.5005
R27736 VSS.n2606 VSS.n2461 4.5005
R27737 VSS.n2609 VSS.n2461 4.5005
R27738 VSS.n2611 VSS.n2461 4.5005
R27739 VSS.n2612 VSS.n2461 4.5005
R27740 VSS.n2614 VSS.n2461 4.5005
R27741 VSS.n2617 VSS.n2461 4.5005
R27742 VSS.n2619 VSS.n2461 4.5005
R27743 VSS.n2620 VSS.n2461 4.5005
R27744 VSS.n2622 VSS.n2461 4.5005
R27745 VSS.n2625 VSS.n2461 4.5005
R27746 VSS.n2627 VSS.n2461 4.5005
R27747 VSS.n2628 VSS.n2461 4.5005
R27748 VSS.n2630 VSS.n2461 4.5005
R27749 VSS.n2633 VSS.n2461 4.5005
R27750 VSS.n2635 VSS.n2461 4.5005
R27751 VSS.n2636 VSS.n2461 4.5005
R27752 VSS.n2638 VSS.n2461 4.5005
R27753 VSS.n2640 VSS.n2461 4.5005
R27754 VSS.n2642 VSS.n2461 4.5005
R27755 VSS.n2643 VSS.n2461 4.5005
R27756 VSS.n2645 VSS.n2461 4.5005
R27757 VSS.n2648 VSS.n2461 4.5005
R27758 VSS.n2650 VSS.n2461 4.5005
R27759 VSS.n2651 VSS.n2461 4.5005
R27760 VSS.n2653 VSS.n2461 4.5005
R27761 VSS.n2656 VSS.n2461 4.5005
R27762 VSS.n2658 VSS.n2461 4.5005
R27763 VSS.n2659 VSS.n2461 4.5005
R27764 VSS.n2661 VSS.n2461 4.5005
R27765 VSS.n2664 VSS.n2461 4.5005
R27766 VSS.n2666 VSS.n2461 4.5005
R27767 VSS.n2667 VSS.n2461 4.5005
R27768 VSS.n2669 VSS.n2461 4.5005
R27769 VSS.n2672 VSS.n2461 4.5005
R27770 VSS.n2674 VSS.n2461 4.5005
R27771 VSS.n2675 VSS.n2461 4.5005
R27772 VSS.n2677 VSS.n2461 4.5005
R27773 VSS.n2680 VSS.n2461 4.5005
R27774 VSS.n2682 VSS.n2461 4.5005
R27775 VSS.n2683 VSS.n2461 4.5005
R27776 VSS.n2685 VSS.n2461 4.5005
R27777 VSS.n2688 VSS.n2461 4.5005
R27778 VSS.n2690 VSS.n2461 4.5005
R27779 VSS.n2691 VSS.n2461 4.5005
R27780 VSS.n2693 VSS.n2461 4.5005
R27781 VSS.n2696 VSS.n2461 4.5005
R27782 VSS.n2698 VSS.n2461 4.5005
R27783 VSS.n2699 VSS.n2461 4.5005
R27784 VSS.n2701 VSS.n2461 4.5005
R27785 VSS.n2704 VSS.n2461 4.5005
R27786 VSS.n2706 VSS.n2461 4.5005
R27787 VSS.n2707 VSS.n2461 4.5005
R27788 VSS.n2709 VSS.n2461 4.5005
R27789 VSS.n2712 VSS.n2461 4.5005
R27790 VSS.n2714 VSS.n2461 4.5005
R27791 VSS.n2715 VSS.n2461 4.5005
R27792 VSS.n2717 VSS.n2461 4.5005
R27793 VSS.n2720 VSS.n2461 4.5005
R27794 VSS.n2722 VSS.n2461 4.5005
R27795 VSS.n2723 VSS.n2461 4.5005
R27796 VSS.n2725 VSS.n2461 4.5005
R27797 VSS.n2793 VSS.n2461 4.5005
R27798 VSS.n2859 VSS.n2461 4.5005
R27799 VSS.n3051 VSS.n2370 4.5005
R27800 VSS.n2370 VSS.n2351 4.5005
R27801 VSS.n2483 VSS.n2370 4.5005
R27802 VSS.n2484 VSS.n2370 4.5005
R27803 VSS.n2486 VSS.n2370 4.5005
R27804 VSS.n2489 VSS.n2370 4.5005
R27805 VSS.n2491 VSS.n2370 4.5005
R27806 VSS.n2492 VSS.n2370 4.5005
R27807 VSS.n2494 VSS.n2370 4.5005
R27808 VSS.n2497 VSS.n2370 4.5005
R27809 VSS.n2499 VSS.n2370 4.5005
R27810 VSS.n2500 VSS.n2370 4.5005
R27811 VSS.n2502 VSS.n2370 4.5005
R27812 VSS.n2505 VSS.n2370 4.5005
R27813 VSS.n2507 VSS.n2370 4.5005
R27814 VSS.n2508 VSS.n2370 4.5005
R27815 VSS.n2510 VSS.n2370 4.5005
R27816 VSS.n2513 VSS.n2370 4.5005
R27817 VSS.n2515 VSS.n2370 4.5005
R27818 VSS.n2516 VSS.n2370 4.5005
R27819 VSS.n2518 VSS.n2370 4.5005
R27820 VSS.n2521 VSS.n2370 4.5005
R27821 VSS.n2523 VSS.n2370 4.5005
R27822 VSS.n2524 VSS.n2370 4.5005
R27823 VSS.n2526 VSS.n2370 4.5005
R27824 VSS.n2529 VSS.n2370 4.5005
R27825 VSS.n2531 VSS.n2370 4.5005
R27826 VSS.n2532 VSS.n2370 4.5005
R27827 VSS.n2534 VSS.n2370 4.5005
R27828 VSS.n2537 VSS.n2370 4.5005
R27829 VSS.n2539 VSS.n2370 4.5005
R27830 VSS.n2540 VSS.n2370 4.5005
R27831 VSS.n2542 VSS.n2370 4.5005
R27832 VSS.n2545 VSS.n2370 4.5005
R27833 VSS.n2547 VSS.n2370 4.5005
R27834 VSS.n2548 VSS.n2370 4.5005
R27835 VSS.n2550 VSS.n2370 4.5005
R27836 VSS.n2553 VSS.n2370 4.5005
R27837 VSS.n2555 VSS.n2370 4.5005
R27838 VSS.n2556 VSS.n2370 4.5005
R27839 VSS.n2558 VSS.n2370 4.5005
R27840 VSS.n2561 VSS.n2370 4.5005
R27841 VSS.n2563 VSS.n2370 4.5005
R27842 VSS.n2564 VSS.n2370 4.5005
R27843 VSS.n2566 VSS.n2370 4.5005
R27844 VSS.n2569 VSS.n2370 4.5005
R27845 VSS.n2571 VSS.n2370 4.5005
R27846 VSS.n2572 VSS.n2370 4.5005
R27847 VSS.n2574 VSS.n2370 4.5005
R27848 VSS.n2577 VSS.n2370 4.5005
R27849 VSS.n2579 VSS.n2370 4.5005
R27850 VSS.n2580 VSS.n2370 4.5005
R27851 VSS.n2582 VSS.n2370 4.5005
R27852 VSS.n2585 VSS.n2370 4.5005
R27853 VSS.n2587 VSS.n2370 4.5005
R27854 VSS.n2588 VSS.n2370 4.5005
R27855 VSS.n2590 VSS.n2370 4.5005
R27856 VSS.n2593 VSS.n2370 4.5005
R27857 VSS.n2595 VSS.n2370 4.5005
R27858 VSS.n2596 VSS.n2370 4.5005
R27859 VSS.n2598 VSS.n2370 4.5005
R27860 VSS.n2601 VSS.n2370 4.5005
R27861 VSS.n2603 VSS.n2370 4.5005
R27862 VSS.n2604 VSS.n2370 4.5005
R27863 VSS.n2606 VSS.n2370 4.5005
R27864 VSS.n2609 VSS.n2370 4.5005
R27865 VSS.n2611 VSS.n2370 4.5005
R27866 VSS.n2612 VSS.n2370 4.5005
R27867 VSS.n2614 VSS.n2370 4.5005
R27868 VSS.n2617 VSS.n2370 4.5005
R27869 VSS.n2619 VSS.n2370 4.5005
R27870 VSS.n2620 VSS.n2370 4.5005
R27871 VSS.n2622 VSS.n2370 4.5005
R27872 VSS.n2625 VSS.n2370 4.5005
R27873 VSS.n2627 VSS.n2370 4.5005
R27874 VSS.n2628 VSS.n2370 4.5005
R27875 VSS.n2630 VSS.n2370 4.5005
R27876 VSS.n2633 VSS.n2370 4.5005
R27877 VSS.n2635 VSS.n2370 4.5005
R27878 VSS.n2636 VSS.n2370 4.5005
R27879 VSS.n2638 VSS.n2370 4.5005
R27880 VSS.n2640 VSS.n2370 4.5005
R27881 VSS.n2642 VSS.n2370 4.5005
R27882 VSS.n2643 VSS.n2370 4.5005
R27883 VSS.n2645 VSS.n2370 4.5005
R27884 VSS.n2648 VSS.n2370 4.5005
R27885 VSS.n2650 VSS.n2370 4.5005
R27886 VSS.n2651 VSS.n2370 4.5005
R27887 VSS.n2653 VSS.n2370 4.5005
R27888 VSS.n2656 VSS.n2370 4.5005
R27889 VSS.n2658 VSS.n2370 4.5005
R27890 VSS.n2659 VSS.n2370 4.5005
R27891 VSS.n2661 VSS.n2370 4.5005
R27892 VSS.n2664 VSS.n2370 4.5005
R27893 VSS.n2666 VSS.n2370 4.5005
R27894 VSS.n2667 VSS.n2370 4.5005
R27895 VSS.n2669 VSS.n2370 4.5005
R27896 VSS.n2672 VSS.n2370 4.5005
R27897 VSS.n2674 VSS.n2370 4.5005
R27898 VSS.n2675 VSS.n2370 4.5005
R27899 VSS.n2677 VSS.n2370 4.5005
R27900 VSS.n2680 VSS.n2370 4.5005
R27901 VSS.n2682 VSS.n2370 4.5005
R27902 VSS.n2683 VSS.n2370 4.5005
R27903 VSS.n2685 VSS.n2370 4.5005
R27904 VSS.n2688 VSS.n2370 4.5005
R27905 VSS.n2690 VSS.n2370 4.5005
R27906 VSS.n2691 VSS.n2370 4.5005
R27907 VSS.n2693 VSS.n2370 4.5005
R27908 VSS.n2696 VSS.n2370 4.5005
R27909 VSS.n2698 VSS.n2370 4.5005
R27910 VSS.n2699 VSS.n2370 4.5005
R27911 VSS.n2701 VSS.n2370 4.5005
R27912 VSS.n2704 VSS.n2370 4.5005
R27913 VSS.n2706 VSS.n2370 4.5005
R27914 VSS.n2707 VSS.n2370 4.5005
R27915 VSS.n2709 VSS.n2370 4.5005
R27916 VSS.n2712 VSS.n2370 4.5005
R27917 VSS.n2714 VSS.n2370 4.5005
R27918 VSS.n2715 VSS.n2370 4.5005
R27919 VSS.n2717 VSS.n2370 4.5005
R27920 VSS.n2720 VSS.n2370 4.5005
R27921 VSS.n2722 VSS.n2370 4.5005
R27922 VSS.n2723 VSS.n2370 4.5005
R27923 VSS.n2725 VSS.n2370 4.5005
R27924 VSS.n2793 VSS.n2370 4.5005
R27925 VSS.n2859 VSS.n2370 4.5005
R27926 VSS.n3051 VSS.n2462 4.5005
R27927 VSS.n2462 VSS.n2351 4.5005
R27928 VSS.n2483 VSS.n2462 4.5005
R27929 VSS.n2484 VSS.n2462 4.5005
R27930 VSS.n2486 VSS.n2462 4.5005
R27931 VSS.n2489 VSS.n2462 4.5005
R27932 VSS.n2491 VSS.n2462 4.5005
R27933 VSS.n2492 VSS.n2462 4.5005
R27934 VSS.n2494 VSS.n2462 4.5005
R27935 VSS.n2497 VSS.n2462 4.5005
R27936 VSS.n2499 VSS.n2462 4.5005
R27937 VSS.n2500 VSS.n2462 4.5005
R27938 VSS.n2502 VSS.n2462 4.5005
R27939 VSS.n2505 VSS.n2462 4.5005
R27940 VSS.n2507 VSS.n2462 4.5005
R27941 VSS.n2508 VSS.n2462 4.5005
R27942 VSS.n2510 VSS.n2462 4.5005
R27943 VSS.n2513 VSS.n2462 4.5005
R27944 VSS.n2515 VSS.n2462 4.5005
R27945 VSS.n2516 VSS.n2462 4.5005
R27946 VSS.n2518 VSS.n2462 4.5005
R27947 VSS.n2521 VSS.n2462 4.5005
R27948 VSS.n2523 VSS.n2462 4.5005
R27949 VSS.n2524 VSS.n2462 4.5005
R27950 VSS.n2526 VSS.n2462 4.5005
R27951 VSS.n2529 VSS.n2462 4.5005
R27952 VSS.n2531 VSS.n2462 4.5005
R27953 VSS.n2532 VSS.n2462 4.5005
R27954 VSS.n2534 VSS.n2462 4.5005
R27955 VSS.n2537 VSS.n2462 4.5005
R27956 VSS.n2539 VSS.n2462 4.5005
R27957 VSS.n2540 VSS.n2462 4.5005
R27958 VSS.n2542 VSS.n2462 4.5005
R27959 VSS.n2545 VSS.n2462 4.5005
R27960 VSS.n2547 VSS.n2462 4.5005
R27961 VSS.n2548 VSS.n2462 4.5005
R27962 VSS.n2550 VSS.n2462 4.5005
R27963 VSS.n2553 VSS.n2462 4.5005
R27964 VSS.n2555 VSS.n2462 4.5005
R27965 VSS.n2556 VSS.n2462 4.5005
R27966 VSS.n2558 VSS.n2462 4.5005
R27967 VSS.n2561 VSS.n2462 4.5005
R27968 VSS.n2563 VSS.n2462 4.5005
R27969 VSS.n2564 VSS.n2462 4.5005
R27970 VSS.n2566 VSS.n2462 4.5005
R27971 VSS.n2569 VSS.n2462 4.5005
R27972 VSS.n2571 VSS.n2462 4.5005
R27973 VSS.n2572 VSS.n2462 4.5005
R27974 VSS.n2574 VSS.n2462 4.5005
R27975 VSS.n2577 VSS.n2462 4.5005
R27976 VSS.n2579 VSS.n2462 4.5005
R27977 VSS.n2580 VSS.n2462 4.5005
R27978 VSS.n2582 VSS.n2462 4.5005
R27979 VSS.n2585 VSS.n2462 4.5005
R27980 VSS.n2587 VSS.n2462 4.5005
R27981 VSS.n2588 VSS.n2462 4.5005
R27982 VSS.n2590 VSS.n2462 4.5005
R27983 VSS.n2593 VSS.n2462 4.5005
R27984 VSS.n2595 VSS.n2462 4.5005
R27985 VSS.n2596 VSS.n2462 4.5005
R27986 VSS.n2598 VSS.n2462 4.5005
R27987 VSS.n2601 VSS.n2462 4.5005
R27988 VSS.n2603 VSS.n2462 4.5005
R27989 VSS.n2604 VSS.n2462 4.5005
R27990 VSS.n2606 VSS.n2462 4.5005
R27991 VSS.n2609 VSS.n2462 4.5005
R27992 VSS.n2611 VSS.n2462 4.5005
R27993 VSS.n2612 VSS.n2462 4.5005
R27994 VSS.n2614 VSS.n2462 4.5005
R27995 VSS.n2617 VSS.n2462 4.5005
R27996 VSS.n2619 VSS.n2462 4.5005
R27997 VSS.n2620 VSS.n2462 4.5005
R27998 VSS.n2622 VSS.n2462 4.5005
R27999 VSS.n2625 VSS.n2462 4.5005
R28000 VSS.n2627 VSS.n2462 4.5005
R28001 VSS.n2628 VSS.n2462 4.5005
R28002 VSS.n2630 VSS.n2462 4.5005
R28003 VSS.n2633 VSS.n2462 4.5005
R28004 VSS.n2635 VSS.n2462 4.5005
R28005 VSS.n2636 VSS.n2462 4.5005
R28006 VSS.n2638 VSS.n2462 4.5005
R28007 VSS.n2640 VSS.n2462 4.5005
R28008 VSS.n2642 VSS.n2462 4.5005
R28009 VSS.n2643 VSS.n2462 4.5005
R28010 VSS.n2645 VSS.n2462 4.5005
R28011 VSS.n2648 VSS.n2462 4.5005
R28012 VSS.n2650 VSS.n2462 4.5005
R28013 VSS.n2651 VSS.n2462 4.5005
R28014 VSS.n2653 VSS.n2462 4.5005
R28015 VSS.n2656 VSS.n2462 4.5005
R28016 VSS.n2658 VSS.n2462 4.5005
R28017 VSS.n2659 VSS.n2462 4.5005
R28018 VSS.n2661 VSS.n2462 4.5005
R28019 VSS.n2664 VSS.n2462 4.5005
R28020 VSS.n2666 VSS.n2462 4.5005
R28021 VSS.n2667 VSS.n2462 4.5005
R28022 VSS.n2669 VSS.n2462 4.5005
R28023 VSS.n2672 VSS.n2462 4.5005
R28024 VSS.n2674 VSS.n2462 4.5005
R28025 VSS.n2675 VSS.n2462 4.5005
R28026 VSS.n2677 VSS.n2462 4.5005
R28027 VSS.n2680 VSS.n2462 4.5005
R28028 VSS.n2682 VSS.n2462 4.5005
R28029 VSS.n2683 VSS.n2462 4.5005
R28030 VSS.n2685 VSS.n2462 4.5005
R28031 VSS.n2688 VSS.n2462 4.5005
R28032 VSS.n2690 VSS.n2462 4.5005
R28033 VSS.n2691 VSS.n2462 4.5005
R28034 VSS.n2693 VSS.n2462 4.5005
R28035 VSS.n2696 VSS.n2462 4.5005
R28036 VSS.n2698 VSS.n2462 4.5005
R28037 VSS.n2699 VSS.n2462 4.5005
R28038 VSS.n2701 VSS.n2462 4.5005
R28039 VSS.n2704 VSS.n2462 4.5005
R28040 VSS.n2706 VSS.n2462 4.5005
R28041 VSS.n2707 VSS.n2462 4.5005
R28042 VSS.n2709 VSS.n2462 4.5005
R28043 VSS.n2712 VSS.n2462 4.5005
R28044 VSS.n2714 VSS.n2462 4.5005
R28045 VSS.n2715 VSS.n2462 4.5005
R28046 VSS.n2717 VSS.n2462 4.5005
R28047 VSS.n2720 VSS.n2462 4.5005
R28048 VSS.n2722 VSS.n2462 4.5005
R28049 VSS.n2723 VSS.n2462 4.5005
R28050 VSS.n2725 VSS.n2462 4.5005
R28051 VSS.n2793 VSS.n2462 4.5005
R28052 VSS.n2859 VSS.n2462 4.5005
R28053 VSS.n3051 VSS.n2369 4.5005
R28054 VSS.n2369 VSS.n2351 4.5005
R28055 VSS.n2483 VSS.n2369 4.5005
R28056 VSS.n2484 VSS.n2369 4.5005
R28057 VSS.n2486 VSS.n2369 4.5005
R28058 VSS.n2489 VSS.n2369 4.5005
R28059 VSS.n2491 VSS.n2369 4.5005
R28060 VSS.n2492 VSS.n2369 4.5005
R28061 VSS.n2494 VSS.n2369 4.5005
R28062 VSS.n2497 VSS.n2369 4.5005
R28063 VSS.n2499 VSS.n2369 4.5005
R28064 VSS.n2500 VSS.n2369 4.5005
R28065 VSS.n2502 VSS.n2369 4.5005
R28066 VSS.n2505 VSS.n2369 4.5005
R28067 VSS.n2507 VSS.n2369 4.5005
R28068 VSS.n2508 VSS.n2369 4.5005
R28069 VSS.n2510 VSS.n2369 4.5005
R28070 VSS.n2513 VSS.n2369 4.5005
R28071 VSS.n2515 VSS.n2369 4.5005
R28072 VSS.n2516 VSS.n2369 4.5005
R28073 VSS.n2518 VSS.n2369 4.5005
R28074 VSS.n2521 VSS.n2369 4.5005
R28075 VSS.n2523 VSS.n2369 4.5005
R28076 VSS.n2524 VSS.n2369 4.5005
R28077 VSS.n2526 VSS.n2369 4.5005
R28078 VSS.n2529 VSS.n2369 4.5005
R28079 VSS.n2531 VSS.n2369 4.5005
R28080 VSS.n2532 VSS.n2369 4.5005
R28081 VSS.n2534 VSS.n2369 4.5005
R28082 VSS.n2537 VSS.n2369 4.5005
R28083 VSS.n2539 VSS.n2369 4.5005
R28084 VSS.n2540 VSS.n2369 4.5005
R28085 VSS.n2542 VSS.n2369 4.5005
R28086 VSS.n2545 VSS.n2369 4.5005
R28087 VSS.n2547 VSS.n2369 4.5005
R28088 VSS.n2548 VSS.n2369 4.5005
R28089 VSS.n2550 VSS.n2369 4.5005
R28090 VSS.n2553 VSS.n2369 4.5005
R28091 VSS.n2555 VSS.n2369 4.5005
R28092 VSS.n2556 VSS.n2369 4.5005
R28093 VSS.n2558 VSS.n2369 4.5005
R28094 VSS.n2561 VSS.n2369 4.5005
R28095 VSS.n2563 VSS.n2369 4.5005
R28096 VSS.n2564 VSS.n2369 4.5005
R28097 VSS.n2566 VSS.n2369 4.5005
R28098 VSS.n2569 VSS.n2369 4.5005
R28099 VSS.n2571 VSS.n2369 4.5005
R28100 VSS.n2572 VSS.n2369 4.5005
R28101 VSS.n2574 VSS.n2369 4.5005
R28102 VSS.n2577 VSS.n2369 4.5005
R28103 VSS.n2579 VSS.n2369 4.5005
R28104 VSS.n2580 VSS.n2369 4.5005
R28105 VSS.n2582 VSS.n2369 4.5005
R28106 VSS.n2585 VSS.n2369 4.5005
R28107 VSS.n2587 VSS.n2369 4.5005
R28108 VSS.n2588 VSS.n2369 4.5005
R28109 VSS.n2590 VSS.n2369 4.5005
R28110 VSS.n2593 VSS.n2369 4.5005
R28111 VSS.n2595 VSS.n2369 4.5005
R28112 VSS.n2596 VSS.n2369 4.5005
R28113 VSS.n2598 VSS.n2369 4.5005
R28114 VSS.n2601 VSS.n2369 4.5005
R28115 VSS.n2603 VSS.n2369 4.5005
R28116 VSS.n2604 VSS.n2369 4.5005
R28117 VSS.n2606 VSS.n2369 4.5005
R28118 VSS.n2609 VSS.n2369 4.5005
R28119 VSS.n2611 VSS.n2369 4.5005
R28120 VSS.n2612 VSS.n2369 4.5005
R28121 VSS.n2614 VSS.n2369 4.5005
R28122 VSS.n2617 VSS.n2369 4.5005
R28123 VSS.n2619 VSS.n2369 4.5005
R28124 VSS.n2620 VSS.n2369 4.5005
R28125 VSS.n2622 VSS.n2369 4.5005
R28126 VSS.n2625 VSS.n2369 4.5005
R28127 VSS.n2627 VSS.n2369 4.5005
R28128 VSS.n2628 VSS.n2369 4.5005
R28129 VSS.n2630 VSS.n2369 4.5005
R28130 VSS.n2633 VSS.n2369 4.5005
R28131 VSS.n2635 VSS.n2369 4.5005
R28132 VSS.n2636 VSS.n2369 4.5005
R28133 VSS.n2638 VSS.n2369 4.5005
R28134 VSS.n2640 VSS.n2369 4.5005
R28135 VSS.n2642 VSS.n2369 4.5005
R28136 VSS.n2643 VSS.n2369 4.5005
R28137 VSS.n2645 VSS.n2369 4.5005
R28138 VSS.n2648 VSS.n2369 4.5005
R28139 VSS.n2650 VSS.n2369 4.5005
R28140 VSS.n2651 VSS.n2369 4.5005
R28141 VSS.n2653 VSS.n2369 4.5005
R28142 VSS.n2656 VSS.n2369 4.5005
R28143 VSS.n2658 VSS.n2369 4.5005
R28144 VSS.n2659 VSS.n2369 4.5005
R28145 VSS.n2661 VSS.n2369 4.5005
R28146 VSS.n2664 VSS.n2369 4.5005
R28147 VSS.n2666 VSS.n2369 4.5005
R28148 VSS.n2667 VSS.n2369 4.5005
R28149 VSS.n2669 VSS.n2369 4.5005
R28150 VSS.n2672 VSS.n2369 4.5005
R28151 VSS.n2674 VSS.n2369 4.5005
R28152 VSS.n2675 VSS.n2369 4.5005
R28153 VSS.n2677 VSS.n2369 4.5005
R28154 VSS.n2680 VSS.n2369 4.5005
R28155 VSS.n2682 VSS.n2369 4.5005
R28156 VSS.n2683 VSS.n2369 4.5005
R28157 VSS.n2685 VSS.n2369 4.5005
R28158 VSS.n2688 VSS.n2369 4.5005
R28159 VSS.n2690 VSS.n2369 4.5005
R28160 VSS.n2691 VSS.n2369 4.5005
R28161 VSS.n2693 VSS.n2369 4.5005
R28162 VSS.n2696 VSS.n2369 4.5005
R28163 VSS.n2698 VSS.n2369 4.5005
R28164 VSS.n2699 VSS.n2369 4.5005
R28165 VSS.n2701 VSS.n2369 4.5005
R28166 VSS.n2704 VSS.n2369 4.5005
R28167 VSS.n2706 VSS.n2369 4.5005
R28168 VSS.n2707 VSS.n2369 4.5005
R28169 VSS.n2709 VSS.n2369 4.5005
R28170 VSS.n2712 VSS.n2369 4.5005
R28171 VSS.n2714 VSS.n2369 4.5005
R28172 VSS.n2715 VSS.n2369 4.5005
R28173 VSS.n2717 VSS.n2369 4.5005
R28174 VSS.n2720 VSS.n2369 4.5005
R28175 VSS.n2722 VSS.n2369 4.5005
R28176 VSS.n2723 VSS.n2369 4.5005
R28177 VSS.n2725 VSS.n2369 4.5005
R28178 VSS.n2793 VSS.n2369 4.5005
R28179 VSS.n2859 VSS.n2369 4.5005
R28180 VSS.n3051 VSS.n2463 4.5005
R28181 VSS.n2463 VSS.n2351 4.5005
R28182 VSS.n2483 VSS.n2463 4.5005
R28183 VSS.n2484 VSS.n2463 4.5005
R28184 VSS.n2486 VSS.n2463 4.5005
R28185 VSS.n2489 VSS.n2463 4.5005
R28186 VSS.n2491 VSS.n2463 4.5005
R28187 VSS.n2492 VSS.n2463 4.5005
R28188 VSS.n2494 VSS.n2463 4.5005
R28189 VSS.n2497 VSS.n2463 4.5005
R28190 VSS.n2499 VSS.n2463 4.5005
R28191 VSS.n2500 VSS.n2463 4.5005
R28192 VSS.n2502 VSS.n2463 4.5005
R28193 VSS.n2505 VSS.n2463 4.5005
R28194 VSS.n2507 VSS.n2463 4.5005
R28195 VSS.n2508 VSS.n2463 4.5005
R28196 VSS.n2510 VSS.n2463 4.5005
R28197 VSS.n2513 VSS.n2463 4.5005
R28198 VSS.n2515 VSS.n2463 4.5005
R28199 VSS.n2516 VSS.n2463 4.5005
R28200 VSS.n2518 VSS.n2463 4.5005
R28201 VSS.n2521 VSS.n2463 4.5005
R28202 VSS.n2523 VSS.n2463 4.5005
R28203 VSS.n2524 VSS.n2463 4.5005
R28204 VSS.n2526 VSS.n2463 4.5005
R28205 VSS.n2529 VSS.n2463 4.5005
R28206 VSS.n2531 VSS.n2463 4.5005
R28207 VSS.n2532 VSS.n2463 4.5005
R28208 VSS.n2534 VSS.n2463 4.5005
R28209 VSS.n2537 VSS.n2463 4.5005
R28210 VSS.n2539 VSS.n2463 4.5005
R28211 VSS.n2540 VSS.n2463 4.5005
R28212 VSS.n2542 VSS.n2463 4.5005
R28213 VSS.n2545 VSS.n2463 4.5005
R28214 VSS.n2547 VSS.n2463 4.5005
R28215 VSS.n2548 VSS.n2463 4.5005
R28216 VSS.n2550 VSS.n2463 4.5005
R28217 VSS.n2553 VSS.n2463 4.5005
R28218 VSS.n2555 VSS.n2463 4.5005
R28219 VSS.n2556 VSS.n2463 4.5005
R28220 VSS.n2558 VSS.n2463 4.5005
R28221 VSS.n2561 VSS.n2463 4.5005
R28222 VSS.n2563 VSS.n2463 4.5005
R28223 VSS.n2564 VSS.n2463 4.5005
R28224 VSS.n2566 VSS.n2463 4.5005
R28225 VSS.n2569 VSS.n2463 4.5005
R28226 VSS.n2571 VSS.n2463 4.5005
R28227 VSS.n2572 VSS.n2463 4.5005
R28228 VSS.n2574 VSS.n2463 4.5005
R28229 VSS.n2577 VSS.n2463 4.5005
R28230 VSS.n2579 VSS.n2463 4.5005
R28231 VSS.n2580 VSS.n2463 4.5005
R28232 VSS.n2582 VSS.n2463 4.5005
R28233 VSS.n2585 VSS.n2463 4.5005
R28234 VSS.n2587 VSS.n2463 4.5005
R28235 VSS.n2588 VSS.n2463 4.5005
R28236 VSS.n2590 VSS.n2463 4.5005
R28237 VSS.n2593 VSS.n2463 4.5005
R28238 VSS.n2595 VSS.n2463 4.5005
R28239 VSS.n2596 VSS.n2463 4.5005
R28240 VSS.n2598 VSS.n2463 4.5005
R28241 VSS.n2601 VSS.n2463 4.5005
R28242 VSS.n2603 VSS.n2463 4.5005
R28243 VSS.n2604 VSS.n2463 4.5005
R28244 VSS.n2606 VSS.n2463 4.5005
R28245 VSS.n2609 VSS.n2463 4.5005
R28246 VSS.n2611 VSS.n2463 4.5005
R28247 VSS.n2612 VSS.n2463 4.5005
R28248 VSS.n2614 VSS.n2463 4.5005
R28249 VSS.n2617 VSS.n2463 4.5005
R28250 VSS.n2619 VSS.n2463 4.5005
R28251 VSS.n2620 VSS.n2463 4.5005
R28252 VSS.n2622 VSS.n2463 4.5005
R28253 VSS.n2625 VSS.n2463 4.5005
R28254 VSS.n2627 VSS.n2463 4.5005
R28255 VSS.n2628 VSS.n2463 4.5005
R28256 VSS.n2630 VSS.n2463 4.5005
R28257 VSS.n2633 VSS.n2463 4.5005
R28258 VSS.n2635 VSS.n2463 4.5005
R28259 VSS.n2636 VSS.n2463 4.5005
R28260 VSS.n2638 VSS.n2463 4.5005
R28261 VSS.n2640 VSS.n2463 4.5005
R28262 VSS.n2642 VSS.n2463 4.5005
R28263 VSS.n2643 VSS.n2463 4.5005
R28264 VSS.n2645 VSS.n2463 4.5005
R28265 VSS.n2648 VSS.n2463 4.5005
R28266 VSS.n2650 VSS.n2463 4.5005
R28267 VSS.n2651 VSS.n2463 4.5005
R28268 VSS.n2653 VSS.n2463 4.5005
R28269 VSS.n2656 VSS.n2463 4.5005
R28270 VSS.n2658 VSS.n2463 4.5005
R28271 VSS.n2659 VSS.n2463 4.5005
R28272 VSS.n2661 VSS.n2463 4.5005
R28273 VSS.n2664 VSS.n2463 4.5005
R28274 VSS.n2666 VSS.n2463 4.5005
R28275 VSS.n2667 VSS.n2463 4.5005
R28276 VSS.n2669 VSS.n2463 4.5005
R28277 VSS.n2672 VSS.n2463 4.5005
R28278 VSS.n2674 VSS.n2463 4.5005
R28279 VSS.n2675 VSS.n2463 4.5005
R28280 VSS.n2677 VSS.n2463 4.5005
R28281 VSS.n2680 VSS.n2463 4.5005
R28282 VSS.n2682 VSS.n2463 4.5005
R28283 VSS.n2683 VSS.n2463 4.5005
R28284 VSS.n2685 VSS.n2463 4.5005
R28285 VSS.n2688 VSS.n2463 4.5005
R28286 VSS.n2690 VSS.n2463 4.5005
R28287 VSS.n2691 VSS.n2463 4.5005
R28288 VSS.n2693 VSS.n2463 4.5005
R28289 VSS.n2696 VSS.n2463 4.5005
R28290 VSS.n2698 VSS.n2463 4.5005
R28291 VSS.n2699 VSS.n2463 4.5005
R28292 VSS.n2701 VSS.n2463 4.5005
R28293 VSS.n2704 VSS.n2463 4.5005
R28294 VSS.n2706 VSS.n2463 4.5005
R28295 VSS.n2707 VSS.n2463 4.5005
R28296 VSS.n2709 VSS.n2463 4.5005
R28297 VSS.n2712 VSS.n2463 4.5005
R28298 VSS.n2714 VSS.n2463 4.5005
R28299 VSS.n2715 VSS.n2463 4.5005
R28300 VSS.n2717 VSS.n2463 4.5005
R28301 VSS.n2720 VSS.n2463 4.5005
R28302 VSS.n2722 VSS.n2463 4.5005
R28303 VSS.n2723 VSS.n2463 4.5005
R28304 VSS.n2725 VSS.n2463 4.5005
R28305 VSS.n2793 VSS.n2463 4.5005
R28306 VSS.n2859 VSS.n2463 4.5005
R28307 VSS.n3051 VSS.n2368 4.5005
R28308 VSS.n2368 VSS.n2351 4.5005
R28309 VSS.n2483 VSS.n2368 4.5005
R28310 VSS.n2484 VSS.n2368 4.5005
R28311 VSS.n2486 VSS.n2368 4.5005
R28312 VSS.n2489 VSS.n2368 4.5005
R28313 VSS.n2491 VSS.n2368 4.5005
R28314 VSS.n2492 VSS.n2368 4.5005
R28315 VSS.n2494 VSS.n2368 4.5005
R28316 VSS.n2497 VSS.n2368 4.5005
R28317 VSS.n2499 VSS.n2368 4.5005
R28318 VSS.n2500 VSS.n2368 4.5005
R28319 VSS.n2502 VSS.n2368 4.5005
R28320 VSS.n2505 VSS.n2368 4.5005
R28321 VSS.n2507 VSS.n2368 4.5005
R28322 VSS.n2508 VSS.n2368 4.5005
R28323 VSS.n2510 VSS.n2368 4.5005
R28324 VSS.n2513 VSS.n2368 4.5005
R28325 VSS.n2515 VSS.n2368 4.5005
R28326 VSS.n2516 VSS.n2368 4.5005
R28327 VSS.n2518 VSS.n2368 4.5005
R28328 VSS.n2521 VSS.n2368 4.5005
R28329 VSS.n2523 VSS.n2368 4.5005
R28330 VSS.n2524 VSS.n2368 4.5005
R28331 VSS.n2526 VSS.n2368 4.5005
R28332 VSS.n2529 VSS.n2368 4.5005
R28333 VSS.n2531 VSS.n2368 4.5005
R28334 VSS.n2532 VSS.n2368 4.5005
R28335 VSS.n2534 VSS.n2368 4.5005
R28336 VSS.n2537 VSS.n2368 4.5005
R28337 VSS.n2539 VSS.n2368 4.5005
R28338 VSS.n2540 VSS.n2368 4.5005
R28339 VSS.n2542 VSS.n2368 4.5005
R28340 VSS.n2545 VSS.n2368 4.5005
R28341 VSS.n2547 VSS.n2368 4.5005
R28342 VSS.n2548 VSS.n2368 4.5005
R28343 VSS.n2550 VSS.n2368 4.5005
R28344 VSS.n2553 VSS.n2368 4.5005
R28345 VSS.n2555 VSS.n2368 4.5005
R28346 VSS.n2556 VSS.n2368 4.5005
R28347 VSS.n2558 VSS.n2368 4.5005
R28348 VSS.n2561 VSS.n2368 4.5005
R28349 VSS.n2563 VSS.n2368 4.5005
R28350 VSS.n2564 VSS.n2368 4.5005
R28351 VSS.n2566 VSS.n2368 4.5005
R28352 VSS.n2569 VSS.n2368 4.5005
R28353 VSS.n2571 VSS.n2368 4.5005
R28354 VSS.n2572 VSS.n2368 4.5005
R28355 VSS.n2574 VSS.n2368 4.5005
R28356 VSS.n2577 VSS.n2368 4.5005
R28357 VSS.n2579 VSS.n2368 4.5005
R28358 VSS.n2580 VSS.n2368 4.5005
R28359 VSS.n2582 VSS.n2368 4.5005
R28360 VSS.n2585 VSS.n2368 4.5005
R28361 VSS.n2587 VSS.n2368 4.5005
R28362 VSS.n2588 VSS.n2368 4.5005
R28363 VSS.n2590 VSS.n2368 4.5005
R28364 VSS.n2593 VSS.n2368 4.5005
R28365 VSS.n2595 VSS.n2368 4.5005
R28366 VSS.n2596 VSS.n2368 4.5005
R28367 VSS.n2598 VSS.n2368 4.5005
R28368 VSS.n2601 VSS.n2368 4.5005
R28369 VSS.n2603 VSS.n2368 4.5005
R28370 VSS.n2604 VSS.n2368 4.5005
R28371 VSS.n2606 VSS.n2368 4.5005
R28372 VSS.n2609 VSS.n2368 4.5005
R28373 VSS.n2611 VSS.n2368 4.5005
R28374 VSS.n2612 VSS.n2368 4.5005
R28375 VSS.n2614 VSS.n2368 4.5005
R28376 VSS.n2617 VSS.n2368 4.5005
R28377 VSS.n2619 VSS.n2368 4.5005
R28378 VSS.n2620 VSS.n2368 4.5005
R28379 VSS.n2622 VSS.n2368 4.5005
R28380 VSS.n2625 VSS.n2368 4.5005
R28381 VSS.n2627 VSS.n2368 4.5005
R28382 VSS.n2628 VSS.n2368 4.5005
R28383 VSS.n2630 VSS.n2368 4.5005
R28384 VSS.n2633 VSS.n2368 4.5005
R28385 VSS.n2635 VSS.n2368 4.5005
R28386 VSS.n2636 VSS.n2368 4.5005
R28387 VSS.n2638 VSS.n2368 4.5005
R28388 VSS.n2640 VSS.n2368 4.5005
R28389 VSS.n2642 VSS.n2368 4.5005
R28390 VSS.n2643 VSS.n2368 4.5005
R28391 VSS.n2645 VSS.n2368 4.5005
R28392 VSS.n2648 VSS.n2368 4.5005
R28393 VSS.n2650 VSS.n2368 4.5005
R28394 VSS.n2651 VSS.n2368 4.5005
R28395 VSS.n2653 VSS.n2368 4.5005
R28396 VSS.n2656 VSS.n2368 4.5005
R28397 VSS.n2658 VSS.n2368 4.5005
R28398 VSS.n2659 VSS.n2368 4.5005
R28399 VSS.n2661 VSS.n2368 4.5005
R28400 VSS.n2664 VSS.n2368 4.5005
R28401 VSS.n2666 VSS.n2368 4.5005
R28402 VSS.n2667 VSS.n2368 4.5005
R28403 VSS.n2669 VSS.n2368 4.5005
R28404 VSS.n2672 VSS.n2368 4.5005
R28405 VSS.n2674 VSS.n2368 4.5005
R28406 VSS.n2675 VSS.n2368 4.5005
R28407 VSS.n2677 VSS.n2368 4.5005
R28408 VSS.n2680 VSS.n2368 4.5005
R28409 VSS.n2682 VSS.n2368 4.5005
R28410 VSS.n2683 VSS.n2368 4.5005
R28411 VSS.n2685 VSS.n2368 4.5005
R28412 VSS.n2688 VSS.n2368 4.5005
R28413 VSS.n2690 VSS.n2368 4.5005
R28414 VSS.n2691 VSS.n2368 4.5005
R28415 VSS.n2693 VSS.n2368 4.5005
R28416 VSS.n2696 VSS.n2368 4.5005
R28417 VSS.n2698 VSS.n2368 4.5005
R28418 VSS.n2699 VSS.n2368 4.5005
R28419 VSS.n2701 VSS.n2368 4.5005
R28420 VSS.n2704 VSS.n2368 4.5005
R28421 VSS.n2706 VSS.n2368 4.5005
R28422 VSS.n2707 VSS.n2368 4.5005
R28423 VSS.n2709 VSS.n2368 4.5005
R28424 VSS.n2712 VSS.n2368 4.5005
R28425 VSS.n2714 VSS.n2368 4.5005
R28426 VSS.n2715 VSS.n2368 4.5005
R28427 VSS.n2717 VSS.n2368 4.5005
R28428 VSS.n2720 VSS.n2368 4.5005
R28429 VSS.n2722 VSS.n2368 4.5005
R28430 VSS.n2723 VSS.n2368 4.5005
R28431 VSS.n2725 VSS.n2368 4.5005
R28432 VSS.n2793 VSS.n2368 4.5005
R28433 VSS.n2859 VSS.n2368 4.5005
R28434 VSS.n3051 VSS.n2464 4.5005
R28435 VSS.n2464 VSS.n2351 4.5005
R28436 VSS.n2483 VSS.n2464 4.5005
R28437 VSS.n2484 VSS.n2464 4.5005
R28438 VSS.n2486 VSS.n2464 4.5005
R28439 VSS.n2489 VSS.n2464 4.5005
R28440 VSS.n2491 VSS.n2464 4.5005
R28441 VSS.n2492 VSS.n2464 4.5005
R28442 VSS.n2494 VSS.n2464 4.5005
R28443 VSS.n2497 VSS.n2464 4.5005
R28444 VSS.n2499 VSS.n2464 4.5005
R28445 VSS.n2500 VSS.n2464 4.5005
R28446 VSS.n2502 VSS.n2464 4.5005
R28447 VSS.n2505 VSS.n2464 4.5005
R28448 VSS.n2507 VSS.n2464 4.5005
R28449 VSS.n2508 VSS.n2464 4.5005
R28450 VSS.n2510 VSS.n2464 4.5005
R28451 VSS.n2513 VSS.n2464 4.5005
R28452 VSS.n2515 VSS.n2464 4.5005
R28453 VSS.n2516 VSS.n2464 4.5005
R28454 VSS.n2518 VSS.n2464 4.5005
R28455 VSS.n2521 VSS.n2464 4.5005
R28456 VSS.n2523 VSS.n2464 4.5005
R28457 VSS.n2524 VSS.n2464 4.5005
R28458 VSS.n2526 VSS.n2464 4.5005
R28459 VSS.n2529 VSS.n2464 4.5005
R28460 VSS.n2531 VSS.n2464 4.5005
R28461 VSS.n2532 VSS.n2464 4.5005
R28462 VSS.n2534 VSS.n2464 4.5005
R28463 VSS.n2537 VSS.n2464 4.5005
R28464 VSS.n2539 VSS.n2464 4.5005
R28465 VSS.n2540 VSS.n2464 4.5005
R28466 VSS.n2542 VSS.n2464 4.5005
R28467 VSS.n2545 VSS.n2464 4.5005
R28468 VSS.n2547 VSS.n2464 4.5005
R28469 VSS.n2548 VSS.n2464 4.5005
R28470 VSS.n2550 VSS.n2464 4.5005
R28471 VSS.n2553 VSS.n2464 4.5005
R28472 VSS.n2555 VSS.n2464 4.5005
R28473 VSS.n2556 VSS.n2464 4.5005
R28474 VSS.n2558 VSS.n2464 4.5005
R28475 VSS.n2561 VSS.n2464 4.5005
R28476 VSS.n2563 VSS.n2464 4.5005
R28477 VSS.n2564 VSS.n2464 4.5005
R28478 VSS.n2566 VSS.n2464 4.5005
R28479 VSS.n2569 VSS.n2464 4.5005
R28480 VSS.n2571 VSS.n2464 4.5005
R28481 VSS.n2572 VSS.n2464 4.5005
R28482 VSS.n2574 VSS.n2464 4.5005
R28483 VSS.n2577 VSS.n2464 4.5005
R28484 VSS.n2579 VSS.n2464 4.5005
R28485 VSS.n2580 VSS.n2464 4.5005
R28486 VSS.n2582 VSS.n2464 4.5005
R28487 VSS.n2585 VSS.n2464 4.5005
R28488 VSS.n2587 VSS.n2464 4.5005
R28489 VSS.n2588 VSS.n2464 4.5005
R28490 VSS.n2590 VSS.n2464 4.5005
R28491 VSS.n2593 VSS.n2464 4.5005
R28492 VSS.n2595 VSS.n2464 4.5005
R28493 VSS.n2596 VSS.n2464 4.5005
R28494 VSS.n2598 VSS.n2464 4.5005
R28495 VSS.n2601 VSS.n2464 4.5005
R28496 VSS.n2603 VSS.n2464 4.5005
R28497 VSS.n2604 VSS.n2464 4.5005
R28498 VSS.n2606 VSS.n2464 4.5005
R28499 VSS.n2609 VSS.n2464 4.5005
R28500 VSS.n2611 VSS.n2464 4.5005
R28501 VSS.n2612 VSS.n2464 4.5005
R28502 VSS.n2614 VSS.n2464 4.5005
R28503 VSS.n2617 VSS.n2464 4.5005
R28504 VSS.n2619 VSS.n2464 4.5005
R28505 VSS.n2620 VSS.n2464 4.5005
R28506 VSS.n2622 VSS.n2464 4.5005
R28507 VSS.n2625 VSS.n2464 4.5005
R28508 VSS.n2627 VSS.n2464 4.5005
R28509 VSS.n2628 VSS.n2464 4.5005
R28510 VSS.n2630 VSS.n2464 4.5005
R28511 VSS.n2633 VSS.n2464 4.5005
R28512 VSS.n2635 VSS.n2464 4.5005
R28513 VSS.n2636 VSS.n2464 4.5005
R28514 VSS.n2638 VSS.n2464 4.5005
R28515 VSS.n2640 VSS.n2464 4.5005
R28516 VSS.n2642 VSS.n2464 4.5005
R28517 VSS.n2643 VSS.n2464 4.5005
R28518 VSS.n2645 VSS.n2464 4.5005
R28519 VSS.n2648 VSS.n2464 4.5005
R28520 VSS.n2650 VSS.n2464 4.5005
R28521 VSS.n2651 VSS.n2464 4.5005
R28522 VSS.n2653 VSS.n2464 4.5005
R28523 VSS.n2656 VSS.n2464 4.5005
R28524 VSS.n2658 VSS.n2464 4.5005
R28525 VSS.n2659 VSS.n2464 4.5005
R28526 VSS.n2661 VSS.n2464 4.5005
R28527 VSS.n2664 VSS.n2464 4.5005
R28528 VSS.n2666 VSS.n2464 4.5005
R28529 VSS.n2667 VSS.n2464 4.5005
R28530 VSS.n2669 VSS.n2464 4.5005
R28531 VSS.n2672 VSS.n2464 4.5005
R28532 VSS.n2674 VSS.n2464 4.5005
R28533 VSS.n2675 VSS.n2464 4.5005
R28534 VSS.n2677 VSS.n2464 4.5005
R28535 VSS.n2680 VSS.n2464 4.5005
R28536 VSS.n2682 VSS.n2464 4.5005
R28537 VSS.n2683 VSS.n2464 4.5005
R28538 VSS.n2685 VSS.n2464 4.5005
R28539 VSS.n2688 VSS.n2464 4.5005
R28540 VSS.n2690 VSS.n2464 4.5005
R28541 VSS.n2691 VSS.n2464 4.5005
R28542 VSS.n2693 VSS.n2464 4.5005
R28543 VSS.n2696 VSS.n2464 4.5005
R28544 VSS.n2698 VSS.n2464 4.5005
R28545 VSS.n2699 VSS.n2464 4.5005
R28546 VSS.n2701 VSS.n2464 4.5005
R28547 VSS.n2704 VSS.n2464 4.5005
R28548 VSS.n2706 VSS.n2464 4.5005
R28549 VSS.n2707 VSS.n2464 4.5005
R28550 VSS.n2709 VSS.n2464 4.5005
R28551 VSS.n2712 VSS.n2464 4.5005
R28552 VSS.n2714 VSS.n2464 4.5005
R28553 VSS.n2715 VSS.n2464 4.5005
R28554 VSS.n2717 VSS.n2464 4.5005
R28555 VSS.n2720 VSS.n2464 4.5005
R28556 VSS.n2722 VSS.n2464 4.5005
R28557 VSS.n2723 VSS.n2464 4.5005
R28558 VSS.n2725 VSS.n2464 4.5005
R28559 VSS.n2793 VSS.n2464 4.5005
R28560 VSS.n2859 VSS.n2464 4.5005
R28561 VSS.n3051 VSS.n2367 4.5005
R28562 VSS.n2367 VSS.n2351 4.5005
R28563 VSS.n2483 VSS.n2367 4.5005
R28564 VSS.n2484 VSS.n2367 4.5005
R28565 VSS.n2486 VSS.n2367 4.5005
R28566 VSS.n2489 VSS.n2367 4.5005
R28567 VSS.n2491 VSS.n2367 4.5005
R28568 VSS.n2492 VSS.n2367 4.5005
R28569 VSS.n2494 VSS.n2367 4.5005
R28570 VSS.n2497 VSS.n2367 4.5005
R28571 VSS.n2499 VSS.n2367 4.5005
R28572 VSS.n2500 VSS.n2367 4.5005
R28573 VSS.n2502 VSS.n2367 4.5005
R28574 VSS.n2505 VSS.n2367 4.5005
R28575 VSS.n2507 VSS.n2367 4.5005
R28576 VSS.n2508 VSS.n2367 4.5005
R28577 VSS.n2510 VSS.n2367 4.5005
R28578 VSS.n2513 VSS.n2367 4.5005
R28579 VSS.n2515 VSS.n2367 4.5005
R28580 VSS.n2516 VSS.n2367 4.5005
R28581 VSS.n2518 VSS.n2367 4.5005
R28582 VSS.n2521 VSS.n2367 4.5005
R28583 VSS.n2523 VSS.n2367 4.5005
R28584 VSS.n2524 VSS.n2367 4.5005
R28585 VSS.n2526 VSS.n2367 4.5005
R28586 VSS.n2529 VSS.n2367 4.5005
R28587 VSS.n2531 VSS.n2367 4.5005
R28588 VSS.n2532 VSS.n2367 4.5005
R28589 VSS.n2534 VSS.n2367 4.5005
R28590 VSS.n2537 VSS.n2367 4.5005
R28591 VSS.n2539 VSS.n2367 4.5005
R28592 VSS.n2540 VSS.n2367 4.5005
R28593 VSS.n2542 VSS.n2367 4.5005
R28594 VSS.n2545 VSS.n2367 4.5005
R28595 VSS.n2547 VSS.n2367 4.5005
R28596 VSS.n2548 VSS.n2367 4.5005
R28597 VSS.n2550 VSS.n2367 4.5005
R28598 VSS.n2553 VSS.n2367 4.5005
R28599 VSS.n2555 VSS.n2367 4.5005
R28600 VSS.n2556 VSS.n2367 4.5005
R28601 VSS.n2558 VSS.n2367 4.5005
R28602 VSS.n2561 VSS.n2367 4.5005
R28603 VSS.n2563 VSS.n2367 4.5005
R28604 VSS.n2564 VSS.n2367 4.5005
R28605 VSS.n2566 VSS.n2367 4.5005
R28606 VSS.n2569 VSS.n2367 4.5005
R28607 VSS.n2571 VSS.n2367 4.5005
R28608 VSS.n2572 VSS.n2367 4.5005
R28609 VSS.n2574 VSS.n2367 4.5005
R28610 VSS.n2577 VSS.n2367 4.5005
R28611 VSS.n2579 VSS.n2367 4.5005
R28612 VSS.n2580 VSS.n2367 4.5005
R28613 VSS.n2582 VSS.n2367 4.5005
R28614 VSS.n2585 VSS.n2367 4.5005
R28615 VSS.n2587 VSS.n2367 4.5005
R28616 VSS.n2588 VSS.n2367 4.5005
R28617 VSS.n2590 VSS.n2367 4.5005
R28618 VSS.n2593 VSS.n2367 4.5005
R28619 VSS.n2595 VSS.n2367 4.5005
R28620 VSS.n2596 VSS.n2367 4.5005
R28621 VSS.n2598 VSS.n2367 4.5005
R28622 VSS.n2601 VSS.n2367 4.5005
R28623 VSS.n2603 VSS.n2367 4.5005
R28624 VSS.n2604 VSS.n2367 4.5005
R28625 VSS.n2606 VSS.n2367 4.5005
R28626 VSS.n2609 VSS.n2367 4.5005
R28627 VSS.n2611 VSS.n2367 4.5005
R28628 VSS.n2612 VSS.n2367 4.5005
R28629 VSS.n2614 VSS.n2367 4.5005
R28630 VSS.n2617 VSS.n2367 4.5005
R28631 VSS.n2619 VSS.n2367 4.5005
R28632 VSS.n2620 VSS.n2367 4.5005
R28633 VSS.n2622 VSS.n2367 4.5005
R28634 VSS.n2625 VSS.n2367 4.5005
R28635 VSS.n2627 VSS.n2367 4.5005
R28636 VSS.n2628 VSS.n2367 4.5005
R28637 VSS.n2630 VSS.n2367 4.5005
R28638 VSS.n2633 VSS.n2367 4.5005
R28639 VSS.n2635 VSS.n2367 4.5005
R28640 VSS.n2636 VSS.n2367 4.5005
R28641 VSS.n2638 VSS.n2367 4.5005
R28642 VSS.n2640 VSS.n2367 4.5005
R28643 VSS.n2642 VSS.n2367 4.5005
R28644 VSS.n2643 VSS.n2367 4.5005
R28645 VSS.n2645 VSS.n2367 4.5005
R28646 VSS.n2648 VSS.n2367 4.5005
R28647 VSS.n2650 VSS.n2367 4.5005
R28648 VSS.n2651 VSS.n2367 4.5005
R28649 VSS.n2653 VSS.n2367 4.5005
R28650 VSS.n2656 VSS.n2367 4.5005
R28651 VSS.n2658 VSS.n2367 4.5005
R28652 VSS.n2659 VSS.n2367 4.5005
R28653 VSS.n2661 VSS.n2367 4.5005
R28654 VSS.n2664 VSS.n2367 4.5005
R28655 VSS.n2666 VSS.n2367 4.5005
R28656 VSS.n2667 VSS.n2367 4.5005
R28657 VSS.n2669 VSS.n2367 4.5005
R28658 VSS.n2672 VSS.n2367 4.5005
R28659 VSS.n2674 VSS.n2367 4.5005
R28660 VSS.n2675 VSS.n2367 4.5005
R28661 VSS.n2677 VSS.n2367 4.5005
R28662 VSS.n2680 VSS.n2367 4.5005
R28663 VSS.n2682 VSS.n2367 4.5005
R28664 VSS.n2683 VSS.n2367 4.5005
R28665 VSS.n2685 VSS.n2367 4.5005
R28666 VSS.n2688 VSS.n2367 4.5005
R28667 VSS.n2690 VSS.n2367 4.5005
R28668 VSS.n2691 VSS.n2367 4.5005
R28669 VSS.n2693 VSS.n2367 4.5005
R28670 VSS.n2696 VSS.n2367 4.5005
R28671 VSS.n2698 VSS.n2367 4.5005
R28672 VSS.n2699 VSS.n2367 4.5005
R28673 VSS.n2701 VSS.n2367 4.5005
R28674 VSS.n2704 VSS.n2367 4.5005
R28675 VSS.n2706 VSS.n2367 4.5005
R28676 VSS.n2707 VSS.n2367 4.5005
R28677 VSS.n2709 VSS.n2367 4.5005
R28678 VSS.n2712 VSS.n2367 4.5005
R28679 VSS.n2714 VSS.n2367 4.5005
R28680 VSS.n2715 VSS.n2367 4.5005
R28681 VSS.n2717 VSS.n2367 4.5005
R28682 VSS.n2720 VSS.n2367 4.5005
R28683 VSS.n2722 VSS.n2367 4.5005
R28684 VSS.n2723 VSS.n2367 4.5005
R28685 VSS.n2725 VSS.n2367 4.5005
R28686 VSS.n2793 VSS.n2367 4.5005
R28687 VSS.n2859 VSS.n2367 4.5005
R28688 VSS.n3051 VSS.n2465 4.5005
R28689 VSS.n2465 VSS.n2351 4.5005
R28690 VSS.n2483 VSS.n2465 4.5005
R28691 VSS.n2484 VSS.n2465 4.5005
R28692 VSS.n2486 VSS.n2465 4.5005
R28693 VSS.n2489 VSS.n2465 4.5005
R28694 VSS.n2491 VSS.n2465 4.5005
R28695 VSS.n2492 VSS.n2465 4.5005
R28696 VSS.n2494 VSS.n2465 4.5005
R28697 VSS.n2497 VSS.n2465 4.5005
R28698 VSS.n2499 VSS.n2465 4.5005
R28699 VSS.n2500 VSS.n2465 4.5005
R28700 VSS.n2502 VSS.n2465 4.5005
R28701 VSS.n2505 VSS.n2465 4.5005
R28702 VSS.n2507 VSS.n2465 4.5005
R28703 VSS.n2508 VSS.n2465 4.5005
R28704 VSS.n2510 VSS.n2465 4.5005
R28705 VSS.n2513 VSS.n2465 4.5005
R28706 VSS.n2515 VSS.n2465 4.5005
R28707 VSS.n2516 VSS.n2465 4.5005
R28708 VSS.n2518 VSS.n2465 4.5005
R28709 VSS.n2521 VSS.n2465 4.5005
R28710 VSS.n2523 VSS.n2465 4.5005
R28711 VSS.n2524 VSS.n2465 4.5005
R28712 VSS.n2526 VSS.n2465 4.5005
R28713 VSS.n2529 VSS.n2465 4.5005
R28714 VSS.n2531 VSS.n2465 4.5005
R28715 VSS.n2532 VSS.n2465 4.5005
R28716 VSS.n2534 VSS.n2465 4.5005
R28717 VSS.n2537 VSS.n2465 4.5005
R28718 VSS.n2539 VSS.n2465 4.5005
R28719 VSS.n2540 VSS.n2465 4.5005
R28720 VSS.n2542 VSS.n2465 4.5005
R28721 VSS.n2545 VSS.n2465 4.5005
R28722 VSS.n2547 VSS.n2465 4.5005
R28723 VSS.n2548 VSS.n2465 4.5005
R28724 VSS.n2550 VSS.n2465 4.5005
R28725 VSS.n2553 VSS.n2465 4.5005
R28726 VSS.n2555 VSS.n2465 4.5005
R28727 VSS.n2556 VSS.n2465 4.5005
R28728 VSS.n2558 VSS.n2465 4.5005
R28729 VSS.n2561 VSS.n2465 4.5005
R28730 VSS.n2563 VSS.n2465 4.5005
R28731 VSS.n2564 VSS.n2465 4.5005
R28732 VSS.n2566 VSS.n2465 4.5005
R28733 VSS.n2569 VSS.n2465 4.5005
R28734 VSS.n2571 VSS.n2465 4.5005
R28735 VSS.n2572 VSS.n2465 4.5005
R28736 VSS.n2574 VSS.n2465 4.5005
R28737 VSS.n2577 VSS.n2465 4.5005
R28738 VSS.n2579 VSS.n2465 4.5005
R28739 VSS.n2580 VSS.n2465 4.5005
R28740 VSS.n2582 VSS.n2465 4.5005
R28741 VSS.n2585 VSS.n2465 4.5005
R28742 VSS.n2587 VSS.n2465 4.5005
R28743 VSS.n2588 VSS.n2465 4.5005
R28744 VSS.n2590 VSS.n2465 4.5005
R28745 VSS.n2593 VSS.n2465 4.5005
R28746 VSS.n2595 VSS.n2465 4.5005
R28747 VSS.n2596 VSS.n2465 4.5005
R28748 VSS.n2598 VSS.n2465 4.5005
R28749 VSS.n2601 VSS.n2465 4.5005
R28750 VSS.n2603 VSS.n2465 4.5005
R28751 VSS.n2604 VSS.n2465 4.5005
R28752 VSS.n2606 VSS.n2465 4.5005
R28753 VSS.n2609 VSS.n2465 4.5005
R28754 VSS.n2611 VSS.n2465 4.5005
R28755 VSS.n2612 VSS.n2465 4.5005
R28756 VSS.n2614 VSS.n2465 4.5005
R28757 VSS.n2617 VSS.n2465 4.5005
R28758 VSS.n2619 VSS.n2465 4.5005
R28759 VSS.n2620 VSS.n2465 4.5005
R28760 VSS.n2622 VSS.n2465 4.5005
R28761 VSS.n2625 VSS.n2465 4.5005
R28762 VSS.n2627 VSS.n2465 4.5005
R28763 VSS.n2628 VSS.n2465 4.5005
R28764 VSS.n2630 VSS.n2465 4.5005
R28765 VSS.n2633 VSS.n2465 4.5005
R28766 VSS.n2635 VSS.n2465 4.5005
R28767 VSS.n2636 VSS.n2465 4.5005
R28768 VSS.n2638 VSS.n2465 4.5005
R28769 VSS.n2640 VSS.n2465 4.5005
R28770 VSS.n2642 VSS.n2465 4.5005
R28771 VSS.n2643 VSS.n2465 4.5005
R28772 VSS.n2645 VSS.n2465 4.5005
R28773 VSS.n2648 VSS.n2465 4.5005
R28774 VSS.n2650 VSS.n2465 4.5005
R28775 VSS.n2651 VSS.n2465 4.5005
R28776 VSS.n2653 VSS.n2465 4.5005
R28777 VSS.n2656 VSS.n2465 4.5005
R28778 VSS.n2658 VSS.n2465 4.5005
R28779 VSS.n2659 VSS.n2465 4.5005
R28780 VSS.n2661 VSS.n2465 4.5005
R28781 VSS.n2664 VSS.n2465 4.5005
R28782 VSS.n2666 VSS.n2465 4.5005
R28783 VSS.n2667 VSS.n2465 4.5005
R28784 VSS.n2669 VSS.n2465 4.5005
R28785 VSS.n2672 VSS.n2465 4.5005
R28786 VSS.n2674 VSS.n2465 4.5005
R28787 VSS.n2675 VSS.n2465 4.5005
R28788 VSS.n2677 VSS.n2465 4.5005
R28789 VSS.n2680 VSS.n2465 4.5005
R28790 VSS.n2682 VSS.n2465 4.5005
R28791 VSS.n2683 VSS.n2465 4.5005
R28792 VSS.n2685 VSS.n2465 4.5005
R28793 VSS.n2688 VSS.n2465 4.5005
R28794 VSS.n2690 VSS.n2465 4.5005
R28795 VSS.n2691 VSS.n2465 4.5005
R28796 VSS.n2693 VSS.n2465 4.5005
R28797 VSS.n2696 VSS.n2465 4.5005
R28798 VSS.n2698 VSS.n2465 4.5005
R28799 VSS.n2699 VSS.n2465 4.5005
R28800 VSS.n2701 VSS.n2465 4.5005
R28801 VSS.n2704 VSS.n2465 4.5005
R28802 VSS.n2706 VSS.n2465 4.5005
R28803 VSS.n2707 VSS.n2465 4.5005
R28804 VSS.n2709 VSS.n2465 4.5005
R28805 VSS.n2712 VSS.n2465 4.5005
R28806 VSS.n2714 VSS.n2465 4.5005
R28807 VSS.n2715 VSS.n2465 4.5005
R28808 VSS.n2717 VSS.n2465 4.5005
R28809 VSS.n2720 VSS.n2465 4.5005
R28810 VSS.n2722 VSS.n2465 4.5005
R28811 VSS.n2723 VSS.n2465 4.5005
R28812 VSS.n2725 VSS.n2465 4.5005
R28813 VSS.n2793 VSS.n2465 4.5005
R28814 VSS.n2859 VSS.n2465 4.5005
R28815 VSS.n3051 VSS.n2366 4.5005
R28816 VSS.n2366 VSS.n2351 4.5005
R28817 VSS.n2483 VSS.n2366 4.5005
R28818 VSS.n2484 VSS.n2366 4.5005
R28819 VSS.n2486 VSS.n2366 4.5005
R28820 VSS.n2489 VSS.n2366 4.5005
R28821 VSS.n2491 VSS.n2366 4.5005
R28822 VSS.n2492 VSS.n2366 4.5005
R28823 VSS.n2494 VSS.n2366 4.5005
R28824 VSS.n2497 VSS.n2366 4.5005
R28825 VSS.n2499 VSS.n2366 4.5005
R28826 VSS.n2500 VSS.n2366 4.5005
R28827 VSS.n2502 VSS.n2366 4.5005
R28828 VSS.n2505 VSS.n2366 4.5005
R28829 VSS.n2507 VSS.n2366 4.5005
R28830 VSS.n2508 VSS.n2366 4.5005
R28831 VSS.n2510 VSS.n2366 4.5005
R28832 VSS.n2513 VSS.n2366 4.5005
R28833 VSS.n2515 VSS.n2366 4.5005
R28834 VSS.n2516 VSS.n2366 4.5005
R28835 VSS.n2518 VSS.n2366 4.5005
R28836 VSS.n2521 VSS.n2366 4.5005
R28837 VSS.n2523 VSS.n2366 4.5005
R28838 VSS.n2524 VSS.n2366 4.5005
R28839 VSS.n2526 VSS.n2366 4.5005
R28840 VSS.n2529 VSS.n2366 4.5005
R28841 VSS.n2531 VSS.n2366 4.5005
R28842 VSS.n2532 VSS.n2366 4.5005
R28843 VSS.n2534 VSS.n2366 4.5005
R28844 VSS.n2537 VSS.n2366 4.5005
R28845 VSS.n2539 VSS.n2366 4.5005
R28846 VSS.n2540 VSS.n2366 4.5005
R28847 VSS.n2542 VSS.n2366 4.5005
R28848 VSS.n2545 VSS.n2366 4.5005
R28849 VSS.n2547 VSS.n2366 4.5005
R28850 VSS.n2548 VSS.n2366 4.5005
R28851 VSS.n2550 VSS.n2366 4.5005
R28852 VSS.n2553 VSS.n2366 4.5005
R28853 VSS.n2555 VSS.n2366 4.5005
R28854 VSS.n2556 VSS.n2366 4.5005
R28855 VSS.n2558 VSS.n2366 4.5005
R28856 VSS.n2561 VSS.n2366 4.5005
R28857 VSS.n2563 VSS.n2366 4.5005
R28858 VSS.n2564 VSS.n2366 4.5005
R28859 VSS.n2566 VSS.n2366 4.5005
R28860 VSS.n2569 VSS.n2366 4.5005
R28861 VSS.n2571 VSS.n2366 4.5005
R28862 VSS.n2572 VSS.n2366 4.5005
R28863 VSS.n2574 VSS.n2366 4.5005
R28864 VSS.n2577 VSS.n2366 4.5005
R28865 VSS.n2579 VSS.n2366 4.5005
R28866 VSS.n2580 VSS.n2366 4.5005
R28867 VSS.n2582 VSS.n2366 4.5005
R28868 VSS.n2585 VSS.n2366 4.5005
R28869 VSS.n2587 VSS.n2366 4.5005
R28870 VSS.n2588 VSS.n2366 4.5005
R28871 VSS.n2590 VSS.n2366 4.5005
R28872 VSS.n2593 VSS.n2366 4.5005
R28873 VSS.n2595 VSS.n2366 4.5005
R28874 VSS.n2596 VSS.n2366 4.5005
R28875 VSS.n2598 VSS.n2366 4.5005
R28876 VSS.n2601 VSS.n2366 4.5005
R28877 VSS.n2603 VSS.n2366 4.5005
R28878 VSS.n2604 VSS.n2366 4.5005
R28879 VSS.n2606 VSS.n2366 4.5005
R28880 VSS.n2609 VSS.n2366 4.5005
R28881 VSS.n2611 VSS.n2366 4.5005
R28882 VSS.n2612 VSS.n2366 4.5005
R28883 VSS.n2614 VSS.n2366 4.5005
R28884 VSS.n2617 VSS.n2366 4.5005
R28885 VSS.n2619 VSS.n2366 4.5005
R28886 VSS.n2620 VSS.n2366 4.5005
R28887 VSS.n2622 VSS.n2366 4.5005
R28888 VSS.n2625 VSS.n2366 4.5005
R28889 VSS.n2627 VSS.n2366 4.5005
R28890 VSS.n2628 VSS.n2366 4.5005
R28891 VSS.n2630 VSS.n2366 4.5005
R28892 VSS.n2633 VSS.n2366 4.5005
R28893 VSS.n2635 VSS.n2366 4.5005
R28894 VSS.n2636 VSS.n2366 4.5005
R28895 VSS.n2638 VSS.n2366 4.5005
R28896 VSS.n2640 VSS.n2366 4.5005
R28897 VSS.n2642 VSS.n2366 4.5005
R28898 VSS.n2643 VSS.n2366 4.5005
R28899 VSS.n2645 VSS.n2366 4.5005
R28900 VSS.n2648 VSS.n2366 4.5005
R28901 VSS.n2650 VSS.n2366 4.5005
R28902 VSS.n2651 VSS.n2366 4.5005
R28903 VSS.n2653 VSS.n2366 4.5005
R28904 VSS.n2656 VSS.n2366 4.5005
R28905 VSS.n2658 VSS.n2366 4.5005
R28906 VSS.n2659 VSS.n2366 4.5005
R28907 VSS.n2661 VSS.n2366 4.5005
R28908 VSS.n2664 VSS.n2366 4.5005
R28909 VSS.n2666 VSS.n2366 4.5005
R28910 VSS.n2667 VSS.n2366 4.5005
R28911 VSS.n2669 VSS.n2366 4.5005
R28912 VSS.n2672 VSS.n2366 4.5005
R28913 VSS.n2674 VSS.n2366 4.5005
R28914 VSS.n2675 VSS.n2366 4.5005
R28915 VSS.n2677 VSS.n2366 4.5005
R28916 VSS.n2680 VSS.n2366 4.5005
R28917 VSS.n2682 VSS.n2366 4.5005
R28918 VSS.n2683 VSS.n2366 4.5005
R28919 VSS.n2685 VSS.n2366 4.5005
R28920 VSS.n2688 VSS.n2366 4.5005
R28921 VSS.n2690 VSS.n2366 4.5005
R28922 VSS.n2691 VSS.n2366 4.5005
R28923 VSS.n2693 VSS.n2366 4.5005
R28924 VSS.n2696 VSS.n2366 4.5005
R28925 VSS.n2698 VSS.n2366 4.5005
R28926 VSS.n2699 VSS.n2366 4.5005
R28927 VSS.n2701 VSS.n2366 4.5005
R28928 VSS.n2704 VSS.n2366 4.5005
R28929 VSS.n2706 VSS.n2366 4.5005
R28930 VSS.n2707 VSS.n2366 4.5005
R28931 VSS.n2709 VSS.n2366 4.5005
R28932 VSS.n2712 VSS.n2366 4.5005
R28933 VSS.n2714 VSS.n2366 4.5005
R28934 VSS.n2715 VSS.n2366 4.5005
R28935 VSS.n2717 VSS.n2366 4.5005
R28936 VSS.n2720 VSS.n2366 4.5005
R28937 VSS.n2722 VSS.n2366 4.5005
R28938 VSS.n2723 VSS.n2366 4.5005
R28939 VSS.n2725 VSS.n2366 4.5005
R28940 VSS.n2793 VSS.n2366 4.5005
R28941 VSS.n2859 VSS.n2366 4.5005
R28942 VSS.n3051 VSS.n2466 4.5005
R28943 VSS.n2466 VSS.n2351 4.5005
R28944 VSS.n2483 VSS.n2466 4.5005
R28945 VSS.n2484 VSS.n2466 4.5005
R28946 VSS.n2486 VSS.n2466 4.5005
R28947 VSS.n2489 VSS.n2466 4.5005
R28948 VSS.n2491 VSS.n2466 4.5005
R28949 VSS.n2492 VSS.n2466 4.5005
R28950 VSS.n2494 VSS.n2466 4.5005
R28951 VSS.n2497 VSS.n2466 4.5005
R28952 VSS.n2499 VSS.n2466 4.5005
R28953 VSS.n2500 VSS.n2466 4.5005
R28954 VSS.n2502 VSS.n2466 4.5005
R28955 VSS.n2505 VSS.n2466 4.5005
R28956 VSS.n2507 VSS.n2466 4.5005
R28957 VSS.n2508 VSS.n2466 4.5005
R28958 VSS.n2510 VSS.n2466 4.5005
R28959 VSS.n2513 VSS.n2466 4.5005
R28960 VSS.n2515 VSS.n2466 4.5005
R28961 VSS.n2516 VSS.n2466 4.5005
R28962 VSS.n2518 VSS.n2466 4.5005
R28963 VSS.n2521 VSS.n2466 4.5005
R28964 VSS.n2523 VSS.n2466 4.5005
R28965 VSS.n2524 VSS.n2466 4.5005
R28966 VSS.n2526 VSS.n2466 4.5005
R28967 VSS.n2529 VSS.n2466 4.5005
R28968 VSS.n2531 VSS.n2466 4.5005
R28969 VSS.n2532 VSS.n2466 4.5005
R28970 VSS.n2534 VSS.n2466 4.5005
R28971 VSS.n2537 VSS.n2466 4.5005
R28972 VSS.n2539 VSS.n2466 4.5005
R28973 VSS.n2540 VSS.n2466 4.5005
R28974 VSS.n2542 VSS.n2466 4.5005
R28975 VSS.n2545 VSS.n2466 4.5005
R28976 VSS.n2547 VSS.n2466 4.5005
R28977 VSS.n2548 VSS.n2466 4.5005
R28978 VSS.n2550 VSS.n2466 4.5005
R28979 VSS.n2553 VSS.n2466 4.5005
R28980 VSS.n2555 VSS.n2466 4.5005
R28981 VSS.n2556 VSS.n2466 4.5005
R28982 VSS.n2558 VSS.n2466 4.5005
R28983 VSS.n2561 VSS.n2466 4.5005
R28984 VSS.n2563 VSS.n2466 4.5005
R28985 VSS.n2564 VSS.n2466 4.5005
R28986 VSS.n2566 VSS.n2466 4.5005
R28987 VSS.n2569 VSS.n2466 4.5005
R28988 VSS.n2571 VSS.n2466 4.5005
R28989 VSS.n2572 VSS.n2466 4.5005
R28990 VSS.n2574 VSS.n2466 4.5005
R28991 VSS.n2577 VSS.n2466 4.5005
R28992 VSS.n2579 VSS.n2466 4.5005
R28993 VSS.n2580 VSS.n2466 4.5005
R28994 VSS.n2582 VSS.n2466 4.5005
R28995 VSS.n2585 VSS.n2466 4.5005
R28996 VSS.n2587 VSS.n2466 4.5005
R28997 VSS.n2588 VSS.n2466 4.5005
R28998 VSS.n2590 VSS.n2466 4.5005
R28999 VSS.n2593 VSS.n2466 4.5005
R29000 VSS.n2595 VSS.n2466 4.5005
R29001 VSS.n2596 VSS.n2466 4.5005
R29002 VSS.n2598 VSS.n2466 4.5005
R29003 VSS.n2601 VSS.n2466 4.5005
R29004 VSS.n2603 VSS.n2466 4.5005
R29005 VSS.n2604 VSS.n2466 4.5005
R29006 VSS.n2606 VSS.n2466 4.5005
R29007 VSS.n2609 VSS.n2466 4.5005
R29008 VSS.n2611 VSS.n2466 4.5005
R29009 VSS.n2612 VSS.n2466 4.5005
R29010 VSS.n2614 VSS.n2466 4.5005
R29011 VSS.n2617 VSS.n2466 4.5005
R29012 VSS.n2619 VSS.n2466 4.5005
R29013 VSS.n2620 VSS.n2466 4.5005
R29014 VSS.n2622 VSS.n2466 4.5005
R29015 VSS.n2625 VSS.n2466 4.5005
R29016 VSS.n2627 VSS.n2466 4.5005
R29017 VSS.n2628 VSS.n2466 4.5005
R29018 VSS.n2630 VSS.n2466 4.5005
R29019 VSS.n2633 VSS.n2466 4.5005
R29020 VSS.n2635 VSS.n2466 4.5005
R29021 VSS.n2636 VSS.n2466 4.5005
R29022 VSS.n2638 VSS.n2466 4.5005
R29023 VSS.n2640 VSS.n2466 4.5005
R29024 VSS.n2642 VSS.n2466 4.5005
R29025 VSS.n2643 VSS.n2466 4.5005
R29026 VSS.n2645 VSS.n2466 4.5005
R29027 VSS.n2648 VSS.n2466 4.5005
R29028 VSS.n2650 VSS.n2466 4.5005
R29029 VSS.n2651 VSS.n2466 4.5005
R29030 VSS.n2653 VSS.n2466 4.5005
R29031 VSS.n2656 VSS.n2466 4.5005
R29032 VSS.n2658 VSS.n2466 4.5005
R29033 VSS.n2659 VSS.n2466 4.5005
R29034 VSS.n2661 VSS.n2466 4.5005
R29035 VSS.n2664 VSS.n2466 4.5005
R29036 VSS.n2666 VSS.n2466 4.5005
R29037 VSS.n2667 VSS.n2466 4.5005
R29038 VSS.n2669 VSS.n2466 4.5005
R29039 VSS.n2672 VSS.n2466 4.5005
R29040 VSS.n2674 VSS.n2466 4.5005
R29041 VSS.n2675 VSS.n2466 4.5005
R29042 VSS.n2677 VSS.n2466 4.5005
R29043 VSS.n2680 VSS.n2466 4.5005
R29044 VSS.n2682 VSS.n2466 4.5005
R29045 VSS.n2683 VSS.n2466 4.5005
R29046 VSS.n2685 VSS.n2466 4.5005
R29047 VSS.n2688 VSS.n2466 4.5005
R29048 VSS.n2690 VSS.n2466 4.5005
R29049 VSS.n2691 VSS.n2466 4.5005
R29050 VSS.n2693 VSS.n2466 4.5005
R29051 VSS.n2696 VSS.n2466 4.5005
R29052 VSS.n2698 VSS.n2466 4.5005
R29053 VSS.n2699 VSS.n2466 4.5005
R29054 VSS.n2701 VSS.n2466 4.5005
R29055 VSS.n2704 VSS.n2466 4.5005
R29056 VSS.n2706 VSS.n2466 4.5005
R29057 VSS.n2707 VSS.n2466 4.5005
R29058 VSS.n2709 VSS.n2466 4.5005
R29059 VSS.n2712 VSS.n2466 4.5005
R29060 VSS.n2714 VSS.n2466 4.5005
R29061 VSS.n2715 VSS.n2466 4.5005
R29062 VSS.n2717 VSS.n2466 4.5005
R29063 VSS.n2720 VSS.n2466 4.5005
R29064 VSS.n2722 VSS.n2466 4.5005
R29065 VSS.n2723 VSS.n2466 4.5005
R29066 VSS.n2725 VSS.n2466 4.5005
R29067 VSS.n2793 VSS.n2466 4.5005
R29068 VSS.n2859 VSS.n2466 4.5005
R29069 VSS.n3051 VSS.n2365 4.5005
R29070 VSS.n2365 VSS.n2351 4.5005
R29071 VSS.n2483 VSS.n2365 4.5005
R29072 VSS.n2484 VSS.n2365 4.5005
R29073 VSS.n2486 VSS.n2365 4.5005
R29074 VSS.n2489 VSS.n2365 4.5005
R29075 VSS.n2491 VSS.n2365 4.5005
R29076 VSS.n2492 VSS.n2365 4.5005
R29077 VSS.n2494 VSS.n2365 4.5005
R29078 VSS.n2497 VSS.n2365 4.5005
R29079 VSS.n2499 VSS.n2365 4.5005
R29080 VSS.n2500 VSS.n2365 4.5005
R29081 VSS.n2502 VSS.n2365 4.5005
R29082 VSS.n2505 VSS.n2365 4.5005
R29083 VSS.n2507 VSS.n2365 4.5005
R29084 VSS.n2508 VSS.n2365 4.5005
R29085 VSS.n2510 VSS.n2365 4.5005
R29086 VSS.n2513 VSS.n2365 4.5005
R29087 VSS.n2515 VSS.n2365 4.5005
R29088 VSS.n2516 VSS.n2365 4.5005
R29089 VSS.n2518 VSS.n2365 4.5005
R29090 VSS.n2521 VSS.n2365 4.5005
R29091 VSS.n2523 VSS.n2365 4.5005
R29092 VSS.n2524 VSS.n2365 4.5005
R29093 VSS.n2526 VSS.n2365 4.5005
R29094 VSS.n2529 VSS.n2365 4.5005
R29095 VSS.n2531 VSS.n2365 4.5005
R29096 VSS.n2532 VSS.n2365 4.5005
R29097 VSS.n2534 VSS.n2365 4.5005
R29098 VSS.n2537 VSS.n2365 4.5005
R29099 VSS.n2539 VSS.n2365 4.5005
R29100 VSS.n2540 VSS.n2365 4.5005
R29101 VSS.n2542 VSS.n2365 4.5005
R29102 VSS.n2545 VSS.n2365 4.5005
R29103 VSS.n2547 VSS.n2365 4.5005
R29104 VSS.n2548 VSS.n2365 4.5005
R29105 VSS.n2550 VSS.n2365 4.5005
R29106 VSS.n2553 VSS.n2365 4.5005
R29107 VSS.n2555 VSS.n2365 4.5005
R29108 VSS.n2556 VSS.n2365 4.5005
R29109 VSS.n2558 VSS.n2365 4.5005
R29110 VSS.n2561 VSS.n2365 4.5005
R29111 VSS.n2563 VSS.n2365 4.5005
R29112 VSS.n2564 VSS.n2365 4.5005
R29113 VSS.n2566 VSS.n2365 4.5005
R29114 VSS.n2569 VSS.n2365 4.5005
R29115 VSS.n2571 VSS.n2365 4.5005
R29116 VSS.n2572 VSS.n2365 4.5005
R29117 VSS.n2574 VSS.n2365 4.5005
R29118 VSS.n2577 VSS.n2365 4.5005
R29119 VSS.n2579 VSS.n2365 4.5005
R29120 VSS.n2580 VSS.n2365 4.5005
R29121 VSS.n2582 VSS.n2365 4.5005
R29122 VSS.n2585 VSS.n2365 4.5005
R29123 VSS.n2587 VSS.n2365 4.5005
R29124 VSS.n2588 VSS.n2365 4.5005
R29125 VSS.n2590 VSS.n2365 4.5005
R29126 VSS.n2593 VSS.n2365 4.5005
R29127 VSS.n2595 VSS.n2365 4.5005
R29128 VSS.n2596 VSS.n2365 4.5005
R29129 VSS.n2598 VSS.n2365 4.5005
R29130 VSS.n2601 VSS.n2365 4.5005
R29131 VSS.n2603 VSS.n2365 4.5005
R29132 VSS.n2604 VSS.n2365 4.5005
R29133 VSS.n2606 VSS.n2365 4.5005
R29134 VSS.n2609 VSS.n2365 4.5005
R29135 VSS.n2611 VSS.n2365 4.5005
R29136 VSS.n2612 VSS.n2365 4.5005
R29137 VSS.n2614 VSS.n2365 4.5005
R29138 VSS.n2617 VSS.n2365 4.5005
R29139 VSS.n2619 VSS.n2365 4.5005
R29140 VSS.n2620 VSS.n2365 4.5005
R29141 VSS.n2622 VSS.n2365 4.5005
R29142 VSS.n2625 VSS.n2365 4.5005
R29143 VSS.n2627 VSS.n2365 4.5005
R29144 VSS.n2628 VSS.n2365 4.5005
R29145 VSS.n2630 VSS.n2365 4.5005
R29146 VSS.n2633 VSS.n2365 4.5005
R29147 VSS.n2635 VSS.n2365 4.5005
R29148 VSS.n2636 VSS.n2365 4.5005
R29149 VSS.n2638 VSS.n2365 4.5005
R29150 VSS.n2640 VSS.n2365 4.5005
R29151 VSS.n2642 VSS.n2365 4.5005
R29152 VSS.n2643 VSS.n2365 4.5005
R29153 VSS.n2645 VSS.n2365 4.5005
R29154 VSS.n2648 VSS.n2365 4.5005
R29155 VSS.n2650 VSS.n2365 4.5005
R29156 VSS.n2651 VSS.n2365 4.5005
R29157 VSS.n2653 VSS.n2365 4.5005
R29158 VSS.n2656 VSS.n2365 4.5005
R29159 VSS.n2658 VSS.n2365 4.5005
R29160 VSS.n2659 VSS.n2365 4.5005
R29161 VSS.n2661 VSS.n2365 4.5005
R29162 VSS.n2664 VSS.n2365 4.5005
R29163 VSS.n2666 VSS.n2365 4.5005
R29164 VSS.n2667 VSS.n2365 4.5005
R29165 VSS.n2669 VSS.n2365 4.5005
R29166 VSS.n2672 VSS.n2365 4.5005
R29167 VSS.n2674 VSS.n2365 4.5005
R29168 VSS.n2675 VSS.n2365 4.5005
R29169 VSS.n2677 VSS.n2365 4.5005
R29170 VSS.n2680 VSS.n2365 4.5005
R29171 VSS.n2682 VSS.n2365 4.5005
R29172 VSS.n2683 VSS.n2365 4.5005
R29173 VSS.n2685 VSS.n2365 4.5005
R29174 VSS.n2688 VSS.n2365 4.5005
R29175 VSS.n2690 VSS.n2365 4.5005
R29176 VSS.n2691 VSS.n2365 4.5005
R29177 VSS.n2693 VSS.n2365 4.5005
R29178 VSS.n2696 VSS.n2365 4.5005
R29179 VSS.n2698 VSS.n2365 4.5005
R29180 VSS.n2699 VSS.n2365 4.5005
R29181 VSS.n2701 VSS.n2365 4.5005
R29182 VSS.n2704 VSS.n2365 4.5005
R29183 VSS.n2706 VSS.n2365 4.5005
R29184 VSS.n2707 VSS.n2365 4.5005
R29185 VSS.n2709 VSS.n2365 4.5005
R29186 VSS.n2712 VSS.n2365 4.5005
R29187 VSS.n2714 VSS.n2365 4.5005
R29188 VSS.n2715 VSS.n2365 4.5005
R29189 VSS.n2717 VSS.n2365 4.5005
R29190 VSS.n2720 VSS.n2365 4.5005
R29191 VSS.n2722 VSS.n2365 4.5005
R29192 VSS.n2723 VSS.n2365 4.5005
R29193 VSS.n2725 VSS.n2365 4.5005
R29194 VSS.n2793 VSS.n2365 4.5005
R29195 VSS.n2859 VSS.n2365 4.5005
R29196 VSS.n3051 VSS.n2467 4.5005
R29197 VSS.n2467 VSS.n2351 4.5005
R29198 VSS.n2483 VSS.n2467 4.5005
R29199 VSS.n2484 VSS.n2467 4.5005
R29200 VSS.n2486 VSS.n2467 4.5005
R29201 VSS.n2489 VSS.n2467 4.5005
R29202 VSS.n2491 VSS.n2467 4.5005
R29203 VSS.n2492 VSS.n2467 4.5005
R29204 VSS.n2494 VSS.n2467 4.5005
R29205 VSS.n2497 VSS.n2467 4.5005
R29206 VSS.n2499 VSS.n2467 4.5005
R29207 VSS.n2500 VSS.n2467 4.5005
R29208 VSS.n2502 VSS.n2467 4.5005
R29209 VSS.n2505 VSS.n2467 4.5005
R29210 VSS.n2507 VSS.n2467 4.5005
R29211 VSS.n2508 VSS.n2467 4.5005
R29212 VSS.n2510 VSS.n2467 4.5005
R29213 VSS.n2513 VSS.n2467 4.5005
R29214 VSS.n2515 VSS.n2467 4.5005
R29215 VSS.n2516 VSS.n2467 4.5005
R29216 VSS.n2518 VSS.n2467 4.5005
R29217 VSS.n2521 VSS.n2467 4.5005
R29218 VSS.n2523 VSS.n2467 4.5005
R29219 VSS.n2524 VSS.n2467 4.5005
R29220 VSS.n2526 VSS.n2467 4.5005
R29221 VSS.n2529 VSS.n2467 4.5005
R29222 VSS.n2531 VSS.n2467 4.5005
R29223 VSS.n2532 VSS.n2467 4.5005
R29224 VSS.n2534 VSS.n2467 4.5005
R29225 VSS.n2537 VSS.n2467 4.5005
R29226 VSS.n2539 VSS.n2467 4.5005
R29227 VSS.n2540 VSS.n2467 4.5005
R29228 VSS.n2542 VSS.n2467 4.5005
R29229 VSS.n2545 VSS.n2467 4.5005
R29230 VSS.n2547 VSS.n2467 4.5005
R29231 VSS.n2548 VSS.n2467 4.5005
R29232 VSS.n2550 VSS.n2467 4.5005
R29233 VSS.n2553 VSS.n2467 4.5005
R29234 VSS.n2555 VSS.n2467 4.5005
R29235 VSS.n2556 VSS.n2467 4.5005
R29236 VSS.n2558 VSS.n2467 4.5005
R29237 VSS.n2561 VSS.n2467 4.5005
R29238 VSS.n2563 VSS.n2467 4.5005
R29239 VSS.n2564 VSS.n2467 4.5005
R29240 VSS.n2566 VSS.n2467 4.5005
R29241 VSS.n2569 VSS.n2467 4.5005
R29242 VSS.n2571 VSS.n2467 4.5005
R29243 VSS.n2572 VSS.n2467 4.5005
R29244 VSS.n2574 VSS.n2467 4.5005
R29245 VSS.n2577 VSS.n2467 4.5005
R29246 VSS.n2579 VSS.n2467 4.5005
R29247 VSS.n2580 VSS.n2467 4.5005
R29248 VSS.n2582 VSS.n2467 4.5005
R29249 VSS.n2585 VSS.n2467 4.5005
R29250 VSS.n2587 VSS.n2467 4.5005
R29251 VSS.n2588 VSS.n2467 4.5005
R29252 VSS.n2590 VSS.n2467 4.5005
R29253 VSS.n2593 VSS.n2467 4.5005
R29254 VSS.n2595 VSS.n2467 4.5005
R29255 VSS.n2596 VSS.n2467 4.5005
R29256 VSS.n2598 VSS.n2467 4.5005
R29257 VSS.n2601 VSS.n2467 4.5005
R29258 VSS.n2603 VSS.n2467 4.5005
R29259 VSS.n2604 VSS.n2467 4.5005
R29260 VSS.n2606 VSS.n2467 4.5005
R29261 VSS.n2609 VSS.n2467 4.5005
R29262 VSS.n2611 VSS.n2467 4.5005
R29263 VSS.n2612 VSS.n2467 4.5005
R29264 VSS.n2614 VSS.n2467 4.5005
R29265 VSS.n2617 VSS.n2467 4.5005
R29266 VSS.n2619 VSS.n2467 4.5005
R29267 VSS.n2620 VSS.n2467 4.5005
R29268 VSS.n2622 VSS.n2467 4.5005
R29269 VSS.n2625 VSS.n2467 4.5005
R29270 VSS.n2627 VSS.n2467 4.5005
R29271 VSS.n2628 VSS.n2467 4.5005
R29272 VSS.n2630 VSS.n2467 4.5005
R29273 VSS.n2633 VSS.n2467 4.5005
R29274 VSS.n2635 VSS.n2467 4.5005
R29275 VSS.n2636 VSS.n2467 4.5005
R29276 VSS.n2638 VSS.n2467 4.5005
R29277 VSS.n2640 VSS.n2467 4.5005
R29278 VSS.n2642 VSS.n2467 4.5005
R29279 VSS.n2643 VSS.n2467 4.5005
R29280 VSS.n2645 VSS.n2467 4.5005
R29281 VSS.n2648 VSS.n2467 4.5005
R29282 VSS.n2650 VSS.n2467 4.5005
R29283 VSS.n2651 VSS.n2467 4.5005
R29284 VSS.n2653 VSS.n2467 4.5005
R29285 VSS.n2656 VSS.n2467 4.5005
R29286 VSS.n2658 VSS.n2467 4.5005
R29287 VSS.n2659 VSS.n2467 4.5005
R29288 VSS.n2661 VSS.n2467 4.5005
R29289 VSS.n2664 VSS.n2467 4.5005
R29290 VSS.n2666 VSS.n2467 4.5005
R29291 VSS.n2667 VSS.n2467 4.5005
R29292 VSS.n2669 VSS.n2467 4.5005
R29293 VSS.n2672 VSS.n2467 4.5005
R29294 VSS.n2674 VSS.n2467 4.5005
R29295 VSS.n2675 VSS.n2467 4.5005
R29296 VSS.n2677 VSS.n2467 4.5005
R29297 VSS.n2680 VSS.n2467 4.5005
R29298 VSS.n2682 VSS.n2467 4.5005
R29299 VSS.n2683 VSS.n2467 4.5005
R29300 VSS.n2685 VSS.n2467 4.5005
R29301 VSS.n2688 VSS.n2467 4.5005
R29302 VSS.n2690 VSS.n2467 4.5005
R29303 VSS.n2691 VSS.n2467 4.5005
R29304 VSS.n2693 VSS.n2467 4.5005
R29305 VSS.n2696 VSS.n2467 4.5005
R29306 VSS.n2698 VSS.n2467 4.5005
R29307 VSS.n2699 VSS.n2467 4.5005
R29308 VSS.n2701 VSS.n2467 4.5005
R29309 VSS.n2704 VSS.n2467 4.5005
R29310 VSS.n2706 VSS.n2467 4.5005
R29311 VSS.n2707 VSS.n2467 4.5005
R29312 VSS.n2709 VSS.n2467 4.5005
R29313 VSS.n2712 VSS.n2467 4.5005
R29314 VSS.n2714 VSS.n2467 4.5005
R29315 VSS.n2715 VSS.n2467 4.5005
R29316 VSS.n2717 VSS.n2467 4.5005
R29317 VSS.n2720 VSS.n2467 4.5005
R29318 VSS.n2722 VSS.n2467 4.5005
R29319 VSS.n2723 VSS.n2467 4.5005
R29320 VSS.n2725 VSS.n2467 4.5005
R29321 VSS.n2793 VSS.n2467 4.5005
R29322 VSS.n2859 VSS.n2467 4.5005
R29323 VSS.n3051 VSS.n2364 4.5005
R29324 VSS.n2364 VSS.n2351 4.5005
R29325 VSS.n2483 VSS.n2364 4.5005
R29326 VSS.n2484 VSS.n2364 4.5005
R29327 VSS.n2486 VSS.n2364 4.5005
R29328 VSS.n2489 VSS.n2364 4.5005
R29329 VSS.n2491 VSS.n2364 4.5005
R29330 VSS.n2492 VSS.n2364 4.5005
R29331 VSS.n2494 VSS.n2364 4.5005
R29332 VSS.n2497 VSS.n2364 4.5005
R29333 VSS.n2499 VSS.n2364 4.5005
R29334 VSS.n2500 VSS.n2364 4.5005
R29335 VSS.n2502 VSS.n2364 4.5005
R29336 VSS.n2505 VSS.n2364 4.5005
R29337 VSS.n2507 VSS.n2364 4.5005
R29338 VSS.n2508 VSS.n2364 4.5005
R29339 VSS.n2510 VSS.n2364 4.5005
R29340 VSS.n2513 VSS.n2364 4.5005
R29341 VSS.n2515 VSS.n2364 4.5005
R29342 VSS.n2516 VSS.n2364 4.5005
R29343 VSS.n2518 VSS.n2364 4.5005
R29344 VSS.n2521 VSS.n2364 4.5005
R29345 VSS.n2523 VSS.n2364 4.5005
R29346 VSS.n2524 VSS.n2364 4.5005
R29347 VSS.n2526 VSS.n2364 4.5005
R29348 VSS.n2529 VSS.n2364 4.5005
R29349 VSS.n2531 VSS.n2364 4.5005
R29350 VSS.n2532 VSS.n2364 4.5005
R29351 VSS.n2534 VSS.n2364 4.5005
R29352 VSS.n2537 VSS.n2364 4.5005
R29353 VSS.n2539 VSS.n2364 4.5005
R29354 VSS.n2540 VSS.n2364 4.5005
R29355 VSS.n2542 VSS.n2364 4.5005
R29356 VSS.n2545 VSS.n2364 4.5005
R29357 VSS.n2547 VSS.n2364 4.5005
R29358 VSS.n2548 VSS.n2364 4.5005
R29359 VSS.n2550 VSS.n2364 4.5005
R29360 VSS.n2553 VSS.n2364 4.5005
R29361 VSS.n2555 VSS.n2364 4.5005
R29362 VSS.n2556 VSS.n2364 4.5005
R29363 VSS.n2558 VSS.n2364 4.5005
R29364 VSS.n2561 VSS.n2364 4.5005
R29365 VSS.n2563 VSS.n2364 4.5005
R29366 VSS.n2564 VSS.n2364 4.5005
R29367 VSS.n2566 VSS.n2364 4.5005
R29368 VSS.n2569 VSS.n2364 4.5005
R29369 VSS.n2571 VSS.n2364 4.5005
R29370 VSS.n2572 VSS.n2364 4.5005
R29371 VSS.n2574 VSS.n2364 4.5005
R29372 VSS.n2577 VSS.n2364 4.5005
R29373 VSS.n2579 VSS.n2364 4.5005
R29374 VSS.n2580 VSS.n2364 4.5005
R29375 VSS.n2582 VSS.n2364 4.5005
R29376 VSS.n2585 VSS.n2364 4.5005
R29377 VSS.n2587 VSS.n2364 4.5005
R29378 VSS.n2588 VSS.n2364 4.5005
R29379 VSS.n2590 VSS.n2364 4.5005
R29380 VSS.n2593 VSS.n2364 4.5005
R29381 VSS.n2595 VSS.n2364 4.5005
R29382 VSS.n2596 VSS.n2364 4.5005
R29383 VSS.n2598 VSS.n2364 4.5005
R29384 VSS.n2601 VSS.n2364 4.5005
R29385 VSS.n2603 VSS.n2364 4.5005
R29386 VSS.n2604 VSS.n2364 4.5005
R29387 VSS.n2606 VSS.n2364 4.5005
R29388 VSS.n2609 VSS.n2364 4.5005
R29389 VSS.n2611 VSS.n2364 4.5005
R29390 VSS.n2612 VSS.n2364 4.5005
R29391 VSS.n2614 VSS.n2364 4.5005
R29392 VSS.n2617 VSS.n2364 4.5005
R29393 VSS.n2619 VSS.n2364 4.5005
R29394 VSS.n2620 VSS.n2364 4.5005
R29395 VSS.n2622 VSS.n2364 4.5005
R29396 VSS.n2625 VSS.n2364 4.5005
R29397 VSS.n2627 VSS.n2364 4.5005
R29398 VSS.n2628 VSS.n2364 4.5005
R29399 VSS.n2630 VSS.n2364 4.5005
R29400 VSS.n2633 VSS.n2364 4.5005
R29401 VSS.n2635 VSS.n2364 4.5005
R29402 VSS.n2636 VSS.n2364 4.5005
R29403 VSS.n2638 VSS.n2364 4.5005
R29404 VSS.n2640 VSS.n2364 4.5005
R29405 VSS.n2642 VSS.n2364 4.5005
R29406 VSS.n2643 VSS.n2364 4.5005
R29407 VSS.n2645 VSS.n2364 4.5005
R29408 VSS.n2648 VSS.n2364 4.5005
R29409 VSS.n2650 VSS.n2364 4.5005
R29410 VSS.n2651 VSS.n2364 4.5005
R29411 VSS.n2653 VSS.n2364 4.5005
R29412 VSS.n2656 VSS.n2364 4.5005
R29413 VSS.n2658 VSS.n2364 4.5005
R29414 VSS.n2659 VSS.n2364 4.5005
R29415 VSS.n2661 VSS.n2364 4.5005
R29416 VSS.n2664 VSS.n2364 4.5005
R29417 VSS.n2666 VSS.n2364 4.5005
R29418 VSS.n2667 VSS.n2364 4.5005
R29419 VSS.n2669 VSS.n2364 4.5005
R29420 VSS.n2672 VSS.n2364 4.5005
R29421 VSS.n2674 VSS.n2364 4.5005
R29422 VSS.n2675 VSS.n2364 4.5005
R29423 VSS.n2677 VSS.n2364 4.5005
R29424 VSS.n2680 VSS.n2364 4.5005
R29425 VSS.n2682 VSS.n2364 4.5005
R29426 VSS.n2683 VSS.n2364 4.5005
R29427 VSS.n2685 VSS.n2364 4.5005
R29428 VSS.n2688 VSS.n2364 4.5005
R29429 VSS.n2690 VSS.n2364 4.5005
R29430 VSS.n2691 VSS.n2364 4.5005
R29431 VSS.n2693 VSS.n2364 4.5005
R29432 VSS.n2696 VSS.n2364 4.5005
R29433 VSS.n2698 VSS.n2364 4.5005
R29434 VSS.n2699 VSS.n2364 4.5005
R29435 VSS.n2701 VSS.n2364 4.5005
R29436 VSS.n2704 VSS.n2364 4.5005
R29437 VSS.n2706 VSS.n2364 4.5005
R29438 VSS.n2707 VSS.n2364 4.5005
R29439 VSS.n2709 VSS.n2364 4.5005
R29440 VSS.n2712 VSS.n2364 4.5005
R29441 VSS.n2714 VSS.n2364 4.5005
R29442 VSS.n2715 VSS.n2364 4.5005
R29443 VSS.n2717 VSS.n2364 4.5005
R29444 VSS.n2720 VSS.n2364 4.5005
R29445 VSS.n2722 VSS.n2364 4.5005
R29446 VSS.n2723 VSS.n2364 4.5005
R29447 VSS.n2725 VSS.n2364 4.5005
R29448 VSS.n2793 VSS.n2364 4.5005
R29449 VSS.n2859 VSS.n2364 4.5005
R29450 VSS.n3051 VSS.n2468 4.5005
R29451 VSS.n2468 VSS.n2351 4.5005
R29452 VSS.n2483 VSS.n2468 4.5005
R29453 VSS.n2484 VSS.n2468 4.5005
R29454 VSS.n2486 VSS.n2468 4.5005
R29455 VSS.n2489 VSS.n2468 4.5005
R29456 VSS.n2491 VSS.n2468 4.5005
R29457 VSS.n2492 VSS.n2468 4.5005
R29458 VSS.n2494 VSS.n2468 4.5005
R29459 VSS.n2497 VSS.n2468 4.5005
R29460 VSS.n2499 VSS.n2468 4.5005
R29461 VSS.n2500 VSS.n2468 4.5005
R29462 VSS.n2502 VSS.n2468 4.5005
R29463 VSS.n2505 VSS.n2468 4.5005
R29464 VSS.n2507 VSS.n2468 4.5005
R29465 VSS.n2508 VSS.n2468 4.5005
R29466 VSS.n2510 VSS.n2468 4.5005
R29467 VSS.n2513 VSS.n2468 4.5005
R29468 VSS.n2515 VSS.n2468 4.5005
R29469 VSS.n2516 VSS.n2468 4.5005
R29470 VSS.n2518 VSS.n2468 4.5005
R29471 VSS.n2521 VSS.n2468 4.5005
R29472 VSS.n2523 VSS.n2468 4.5005
R29473 VSS.n2524 VSS.n2468 4.5005
R29474 VSS.n2526 VSS.n2468 4.5005
R29475 VSS.n2529 VSS.n2468 4.5005
R29476 VSS.n2531 VSS.n2468 4.5005
R29477 VSS.n2532 VSS.n2468 4.5005
R29478 VSS.n2534 VSS.n2468 4.5005
R29479 VSS.n2537 VSS.n2468 4.5005
R29480 VSS.n2539 VSS.n2468 4.5005
R29481 VSS.n2540 VSS.n2468 4.5005
R29482 VSS.n2542 VSS.n2468 4.5005
R29483 VSS.n2545 VSS.n2468 4.5005
R29484 VSS.n2547 VSS.n2468 4.5005
R29485 VSS.n2548 VSS.n2468 4.5005
R29486 VSS.n2550 VSS.n2468 4.5005
R29487 VSS.n2553 VSS.n2468 4.5005
R29488 VSS.n2555 VSS.n2468 4.5005
R29489 VSS.n2556 VSS.n2468 4.5005
R29490 VSS.n2558 VSS.n2468 4.5005
R29491 VSS.n2561 VSS.n2468 4.5005
R29492 VSS.n2563 VSS.n2468 4.5005
R29493 VSS.n2564 VSS.n2468 4.5005
R29494 VSS.n2566 VSS.n2468 4.5005
R29495 VSS.n2569 VSS.n2468 4.5005
R29496 VSS.n2571 VSS.n2468 4.5005
R29497 VSS.n2572 VSS.n2468 4.5005
R29498 VSS.n2574 VSS.n2468 4.5005
R29499 VSS.n2577 VSS.n2468 4.5005
R29500 VSS.n2579 VSS.n2468 4.5005
R29501 VSS.n2580 VSS.n2468 4.5005
R29502 VSS.n2582 VSS.n2468 4.5005
R29503 VSS.n2585 VSS.n2468 4.5005
R29504 VSS.n2587 VSS.n2468 4.5005
R29505 VSS.n2588 VSS.n2468 4.5005
R29506 VSS.n2590 VSS.n2468 4.5005
R29507 VSS.n2593 VSS.n2468 4.5005
R29508 VSS.n2595 VSS.n2468 4.5005
R29509 VSS.n2596 VSS.n2468 4.5005
R29510 VSS.n2598 VSS.n2468 4.5005
R29511 VSS.n2601 VSS.n2468 4.5005
R29512 VSS.n2603 VSS.n2468 4.5005
R29513 VSS.n2604 VSS.n2468 4.5005
R29514 VSS.n2606 VSS.n2468 4.5005
R29515 VSS.n2609 VSS.n2468 4.5005
R29516 VSS.n2611 VSS.n2468 4.5005
R29517 VSS.n2612 VSS.n2468 4.5005
R29518 VSS.n2614 VSS.n2468 4.5005
R29519 VSS.n2617 VSS.n2468 4.5005
R29520 VSS.n2619 VSS.n2468 4.5005
R29521 VSS.n2620 VSS.n2468 4.5005
R29522 VSS.n2622 VSS.n2468 4.5005
R29523 VSS.n2625 VSS.n2468 4.5005
R29524 VSS.n2627 VSS.n2468 4.5005
R29525 VSS.n2628 VSS.n2468 4.5005
R29526 VSS.n2630 VSS.n2468 4.5005
R29527 VSS.n2633 VSS.n2468 4.5005
R29528 VSS.n2635 VSS.n2468 4.5005
R29529 VSS.n2636 VSS.n2468 4.5005
R29530 VSS.n2638 VSS.n2468 4.5005
R29531 VSS.n2640 VSS.n2468 4.5005
R29532 VSS.n2642 VSS.n2468 4.5005
R29533 VSS.n2643 VSS.n2468 4.5005
R29534 VSS.n2645 VSS.n2468 4.5005
R29535 VSS.n2648 VSS.n2468 4.5005
R29536 VSS.n2650 VSS.n2468 4.5005
R29537 VSS.n2651 VSS.n2468 4.5005
R29538 VSS.n2653 VSS.n2468 4.5005
R29539 VSS.n2656 VSS.n2468 4.5005
R29540 VSS.n2658 VSS.n2468 4.5005
R29541 VSS.n2659 VSS.n2468 4.5005
R29542 VSS.n2661 VSS.n2468 4.5005
R29543 VSS.n2664 VSS.n2468 4.5005
R29544 VSS.n2666 VSS.n2468 4.5005
R29545 VSS.n2667 VSS.n2468 4.5005
R29546 VSS.n2669 VSS.n2468 4.5005
R29547 VSS.n2672 VSS.n2468 4.5005
R29548 VSS.n2674 VSS.n2468 4.5005
R29549 VSS.n2675 VSS.n2468 4.5005
R29550 VSS.n2677 VSS.n2468 4.5005
R29551 VSS.n2680 VSS.n2468 4.5005
R29552 VSS.n2682 VSS.n2468 4.5005
R29553 VSS.n2683 VSS.n2468 4.5005
R29554 VSS.n2685 VSS.n2468 4.5005
R29555 VSS.n2688 VSS.n2468 4.5005
R29556 VSS.n2690 VSS.n2468 4.5005
R29557 VSS.n2691 VSS.n2468 4.5005
R29558 VSS.n2693 VSS.n2468 4.5005
R29559 VSS.n2696 VSS.n2468 4.5005
R29560 VSS.n2698 VSS.n2468 4.5005
R29561 VSS.n2699 VSS.n2468 4.5005
R29562 VSS.n2701 VSS.n2468 4.5005
R29563 VSS.n2704 VSS.n2468 4.5005
R29564 VSS.n2706 VSS.n2468 4.5005
R29565 VSS.n2707 VSS.n2468 4.5005
R29566 VSS.n2709 VSS.n2468 4.5005
R29567 VSS.n2712 VSS.n2468 4.5005
R29568 VSS.n2714 VSS.n2468 4.5005
R29569 VSS.n2715 VSS.n2468 4.5005
R29570 VSS.n2717 VSS.n2468 4.5005
R29571 VSS.n2720 VSS.n2468 4.5005
R29572 VSS.n2722 VSS.n2468 4.5005
R29573 VSS.n2723 VSS.n2468 4.5005
R29574 VSS.n2725 VSS.n2468 4.5005
R29575 VSS.n2793 VSS.n2468 4.5005
R29576 VSS.n2859 VSS.n2468 4.5005
R29577 VSS.n3051 VSS.n2363 4.5005
R29578 VSS.n2363 VSS.n2351 4.5005
R29579 VSS.n2483 VSS.n2363 4.5005
R29580 VSS.n2484 VSS.n2363 4.5005
R29581 VSS.n2486 VSS.n2363 4.5005
R29582 VSS.n2489 VSS.n2363 4.5005
R29583 VSS.n2491 VSS.n2363 4.5005
R29584 VSS.n2492 VSS.n2363 4.5005
R29585 VSS.n2494 VSS.n2363 4.5005
R29586 VSS.n2497 VSS.n2363 4.5005
R29587 VSS.n2499 VSS.n2363 4.5005
R29588 VSS.n2500 VSS.n2363 4.5005
R29589 VSS.n2502 VSS.n2363 4.5005
R29590 VSS.n2505 VSS.n2363 4.5005
R29591 VSS.n2507 VSS.n2363 4.5005
R29592 VSS.n2508 VSS.n2363 4.5005
R29593 VSS.n2510 VSS.n2363 4.5005
R29594 VSS.n2513 VSS.n2363 4.5005
R29595 VSS.n2515 VSS.n2363 4.5005
R29596 VSS.n2516 VSS.n2363 4.5005
R29597 VSS.n2518 VSS.n2363 4.5005
R29598 VSS.n2521 VSS.n2363 4.5005
R29599 VSS.n2523 VSS.n2363 4.5005
R29600 VSS.n2524 VSS.n2363 4.5005
R29601 VSS.n2526 VSS.n2363 4.5005
R29602 VSS.n2529 VSS.n2363 4.5005
R29603 VSS.n2531 VSS.n2363 4.5005
R29604 VSS.n2532 VSS.n2363 4.5005
R29605 VSS.n2534 VSS.n2363 4.5005
R29606 VSS.n2537 VSS.n2363 4.5005
R29607 VSS.n2539 VSS.n2363 4.5005
R29608 VSS.n2540 VSS.n2363 4.5005
R29609 VSS.n2542 VSS.n2363 4.5005
R29610 VSS.n2545 VSS.n2363 4.5005
R29611 VSS.n2547 VSS.n2363 4.5005
R29612 VSS.n2548 VSS.n2363 4.5005
R29613 VSS.n2550 VSS.n2363 4.5005
R29614 VSS.n2553 VSS.n2363 4.5005
R29615 VSS.n2555 VSS.n2363 4.5005
R29616 VSS.n2556 VSS.n2363 4.5005
R29617 VSS.n2558 VSS.n2363 4.5005
R29618 VSS.n2561 VSS.n2363 4.5005
R29619 VSS.n2563 VSS.n2363 4.5005
R29620 VSS.n2564 VSS.n2363 4.5005
R29621 VSS.n2566 VSS.n2363 4.5005
R29622 VSS.n2569 VSS.n2363 4.5005
R29623 VSS.n2571 VSS.n2363 4.5005
R29624 VSS.n2572 VSS.n2363 4.5005
R29625 VSS.n2574 VSS.n2363 4.5005
R29626 VSS.n2577 VSS.n2363 4.5005
R29627 VSS.n2579 VSS.n2363 4.5005
R29628 VSS.n2580 VSS.n2363 4.5005
R29629 VSS.n2582 VSS.n2363 4.5005
R29630 VSS.n2585 VSS.n2363 4.5005
R29631 VSS.n2587 VSS.n2363 4.5005
R29632 VSS.n2588 VSS.n2363 4.5005
R29633 VSS.n2590 VSS.n2363 4.5005
R29634 VSS.n2593 VSS.n2363 4.5005
R29635 VSS.n2595 VSS.n2363 4.5005
R29636 VSS.n2596 VSS.n2363 4.5005
R29637 VSS.n2598 VSS.n2363 4.5005
R29638 VSS.n2601 VSS.n2363 4.5005
R29639 VSS.n2603 VSS.n2363 4.5005
R29640 VSS.n2604 VSS.n2363 4.5005
R29641 VSS.n2606 VSS.n2363 4.5005
R29642 VSS.n2609 VSS.n2363 4.5005
R29643 VSS.n2611 VSS.n2363 4.5005
R29644 VSS.n2612 VSS.n2363 4.5005
R29645 VSS.n2614 VSS.n2363 4.5005
R29646 VSS.n2617 VSS.n2363 4.5005
R29647 VSS.n2619 VSS.n2363 4.5005
R29648 VSS.n2620 VSS.n2363 4.5005
R29649 VSS.n2622 VSS.n2363 4.5005
R29650 VSS.n2625 VSS.n2363 4.5005
R29651 VSS.n2627 VSS.n2363 4.5005
R29652 VSS.n2628 VSS.n2363 4.5005
R29653 VSS.n2630 VSS.n2363 4.5005
R29654 VSS.n2633 VSS.n2363 4.5005
R29655 VSS.n2635 VSS.n2363 4.5005
R29656 VSS.n2636 VSS.n2363 4.5005
R29657 VSS.n2638 VSS.n2363 4.5005
R29658 VSS.n2640 VSS.n2363 4.5005
R29659 VSS.n2642 VSS.n2363 4.5005
R29660 VSS.n2643 VSS.n2363 4.5005
R29661 VSS.n2645 VSS.n2363 4.5005
R29662 VSS.n2648 VSS.n2363 4.5005
R29663 VSS.n2650 VSS.n2363 4.5005
R29664 VSS.n2651 VSS.n2363 4.5005
R29665 VSS.n2653 VSS.n2363 4.5005
R29666 VSS.n2656 VSS.n2363 4.5005
R29667 VSS.n2658 VSS.n2363 4.5005
R29668 VSS.n2659 VSS.n2363 4.5005
R29669 VSS.n2661 VSS.n2363 4.5005
R29670 VSS.n2664 VSS.n2363 4.5005
R29671 VSS.n2666 VSS.n2363 4.5005
R29672 VSS.n2667 VSS.n2363 4.5005
R29673 VSS.n2669 VSS.n2363 4.5005
R29674 VSS.n2672 VSS.n2363 4.5005
R29675 VSS.n2674 VSS.n2363 4.5005
R29676 VSS.n2675 VSS.n2363 4.5005
R29677 VSS.n2677 VSS.n2363 4.5005
R29678 VSS.n2680 VSS.n2363 4.5005
R29679 VSS.n2682 VSS.n2363 4.5005
R29680 VSS.n2683 VSS.n2363 4.5005
R29681 VSS.n2685 VSS.n2363 4.5005
R29682 VSS.n2688 VSS.n2363 4.5005
R29683 VSS.n2690 VSS.n2363 4.5005
R29684 VSS.n2691 VSS.n2363 4.5005
R29685 VSS.n2693 VSS.n2363 4.5005
R29686 VSS.n2696 VSS.n2363 4.5005
R29687 VSS.n2698 VSS.n2363 4.5005
R29688 VSS.n2699 VSS.n2363 4.5005
R29689 VSS.n2701 VSS.n2363 4.5005
R29690 VSS.n2704 VSS.n2363 4.5005
R29691 VSS.n2706 VSS.n2363 4.5005
R29692 VSS.n2707 VSS.n2363 4.5005
R29693 VSS.n2709 VSS.n2363 4.5005
R29694 VSS.n2712 VSS.n2363 4.5005
R29695 VSS.n2714 VSS.n2363 4.5005
R29696 VSS.n2715 VSS.n2363 4.5005
R29697 VSS.n2717 VSS.n2363 4.5005
R29698 VSS.n2720 VSS.n2363 4.5005
R29699 VSS.n2722 VSS.n2363 4.5005
R29700 VSS.n2723 VSS.n2363 4.5005
R29701 VSS.n2725 VSS.n2363 4.5005
R29702 VSS.n2793 VSS.n2363 4.5005
R29703 VSS.n2859 VSS.n2363 4.5005
R29704 VSS.n3051 VSS.n2469 4.5005
R29705 VSS.n2469 VSS.n2351 4.5005
R29706 VSS.n2483 VSS.n2469 4.5005
R29707 VSS.n2484 VSS.n2469 4.5005
R29708 VSS.n2486 VSS.n2469 4.5005
R29709 VSS.n2489 VSS.n2469 4.5005
R29710 VSS.n2491 VSS.n2469 4.5005
R29711 VSS.n2492 VSS.n2469 4.5005
R29712 VSS.n2494 VSS.n2469 4.5005
R29713 VSS.n2497 VSS.n2469 4.5005
R29714 VSS.n2499 VSS.n2469 4.5005
R29715 VSS.n2500 VSS.n2469 4.5005
R29716 VSS.n2502 VSS.n2469 4.5005
R29717 VSS.n2505 VSS.n2469 4.5005
R29718 VSS.n2507 VSS.n2469 4.5005
R29719 VSS.n2508 VSS.n2469 4.5005
R29720 VSS.n2510 VSS.n2469 4.5005
R29721 VSS.n2513 VSS.n2469 4.5005
R29722 VSS.n2515 VSS.n2469 4.5005
R29723 VSS.n2516 VSS.n2469 4.5005
R29724 VSS.n2518 VSS.n2469 4.5005
R29725 VSS.n2521 VSS.n2469 4.5005
R29726 VSS.n2523 VSS.n2469 4.5005
R29727 VSS.n2524 VSS.n2469 4.5005
R29728 VSS.n2526 VSS.n2469 4.5005
R29729 VSS.n2529 VSS.n2469 4.5005
R29730 VSS.n2531 VSS.n2469 4.5005
R29731 VSS.n2532 VSS.n2469 4.5005
R29732 VSS.n2534 VSS.n2469 4.5005
R29733 VSS.n2537 VSS.n2469 4.5005
R29734 VSS.n2539 VSS.n2469 4.5005
R29735 VSS.n2540 VSS.n2469 4.5005
R29736 VSS.n2542 VSS.n2469 4.5005
R29737 VSS.n2545 VSS.n2469 4.5005
R29738 VSS.n2547 VSS.n2469 4.5005
R29739 VSS.n2548 VSS.n2469 4.5005
R29740 VSS.n2550 VSS.n2469 4.5005
R29741 VSS.n2553 VSS.n2469 4.5005
R29742 VSS.n2555 VSS.n2469 4.5005
R29743 VSS.n2556 VSS.n2469 4.5005
R29744 VSS.n2558 VSS.n2469 4.5005
R29745 VSS.n2561 VSS.n2469 4.5005
R29746 VSS.n2563 VSS.n2469 4.5005
R29747 VSS.n2564 VSS.n2469 4.5005
R29748 VSS.n2566 VSS.n2469 4.5005
R29749 VSS.n2569 VSS.n2469 4.5005
R29750 VSS.n2571 VSS.n2469 4.5005
R29751 VSS.n2572 VSS.n2469 4.5005
R29752 VSS.n2574 VSS.n2469 4.5005
R29753 VSS.n2577 VSS.n2469 4.5005
R29754 VSS.n2579 VSS.n2469 4.5005
R29755 VSS.n2580 VSS.n2469 4.5005
R29756 VSS.n2582 VSS.n2469 4.5005
R29757 VSS.n2585 VSS.n2469 4.5005
R29758 VSS.n2587 VSS.n2469 4.5005
R29759 VSS.n2588 VSS.n2469 4.5005
R29760 VSS.n2590 VSS.n2469 4.5005
R29761 VSS.n2593 VSS.n2469 4.5005
R29762 VSS.n2595 VSS.n2469 4.5005
R29763 VSS.n2596 VSS.n2469 4.5005
R29764 VSS.n2598 VSS.n2469 4.5005
R29765 VSS.n2601 VSS.n2469 4.5005
R29766 VSS.n2603 VSS.n2469 4.5005
R29767 VSS.n2604 VSS.n2469 4.5005
R29768 VSS.n2606 VSS.n2469 4.5005
R29769 VSS.n2609 VSS.n2469 4.5005
R29770 VSS.n2611 VSS.n2469 4.5005
R29771 VSS.n2612 VSS.n2469 4.5005
R29772 VSS.n2614 VSS.n2469 4.5005
R29773 VSS.n2617 VSS.n2469 4.5005
R29774 VSS.n2619 VSS.n2469 4.5005
R29775 VSS.n2620 VSS.n2469 4.5005
R29776 VSS.n2622 VSS.n2469 4.5005
R29777 VSS.n2625 VSS.n2469 4.5005
R29778 VSS.n2627 VSS.n2469 4.5005
R29779 VSS.n2628 VSS.n2469 4.5005
R29780 VSS.n2630 VSS.n2469 4.5005
R29781 VSS.n2633 VSS.n2469 4.5005
R29782 VSS.n2635 VSS.n2469 4.5005
R29783 VSS.n2636 VSS.n2469 4.5005
R29784 VSS.n2638 VSS.n2469 4.5005
R29785 VSS.n2640 VSS.n2469 4.5005
R29786 VSS.n2642 VSS.n2469 4.5005
R29787 VSS.n2643 VSS.n2469 4.5005
R29788 VSS.n2645 VSS.n2469 4.5005
R29789 VSS.n2648 VSS.n2469 4.5005
R29790 VSS.n2650 VSS.n2469 4.5005
R29791 VSS.n2651 VSS.n2469 4.5005
R29792 VSS.n2653 VSS.n2469 4.5005
R29793 VSS.n2656 VSS.n2469 4.5005
R29794 VSS.n2658 VSS.n2469 4.5005
R29795 VSS.n2659 VSS.n2469 4.5005
R29796 VSS.n2661 VSS.n2469 4.5005
R29797 VSS.n2664 VSS.n2469 4.5005
R29798 VSS.n2666 VSS.n2469 4.5005
R29799 VSS.n2667 VSS.n2469 4.5005
R29800 VSS.n2669 VSS.n2469 4.5005
R29801 VSS.n2672 VSS.n2469 4.5005
R29802 VSS.n2674 VSS.n2469 4.5005
R29803 VSS.n2675 VSS.n2469 4.5005
R29804 VSS.n2677 VSS.n2469 4.5005
R29805 VSS.n2680 VSS.n2469 4.5005
R29806 VSS.n2682 VSS.n2469 4.5005
R29807 VSS.n2683 VSS.n2469 4.5005
R29808 VSS.n2685 VSS.n2469 4.5005
R29809 VSS.n2688 VSS.n2469 4.5005
R29810 VSS.n2690 VSS.n2469 4.5005
R29811 VSS.n2691 VSS.n2469 4.5005
R29812 VSS.n2693 VSS.n2469 4.5005
R29813 VSS.n2696 VSS.n2469 4.5005
R29814 VSS.n2698 VSS.n2469 4.5005
R29815 VSS.n2699 VSS.n2469 4.5005
R29816 VSS.n2701 VSS.n2469 4.5005
R29817 VSS.n2704 VSS.n2469 4.5005
R29818 VSS.n2706 VSS.n2469 4.5005
R29819 VSS.n2707 VSS.n2469 4.5005
R29820 VSS.n2709 VSS.n2469 4.5005
R29821 VSS.n2712 VSS.n2469 4.5005
R29822 VSS.n2714 VSS.n2469 4.5005
R29823 VSS.n2715 VSS.n2469 4.5005
R29824 VSS.n2717 VSS.n2469 4.5005
R29825 VSS.n2720 VSS.n2469 4.5005
R29826 VSS.n2722 VSS.n2469 4.5005
R29827 VSS.n2723 VSS.n2469 4.5005
R29828 VSS.n2725 VSS.n2469 4.5005
R29829 VSS.n2793 VSS.n2469 4.5005
R29830 VSS.n2859 VSS.n2469 4.5005
R29831 VSS.n3051 VSS.n2362 4.5005
R29832 VSS.n2362 VSS.n2351 4.5005
R29833 VSS.n2483 VSS.n2362 4.5005
R29834 VSS.n2484 VSS.n2362 4.5005
R29835 VSS.n2486 VSS.n2362 4.5005
R29836 VSS.n2489 VSS.n2362 4.5005
R29837 VSS.n2491 VSS.n2362 4.5005
R29838 VSS.n2492 VSS.n2362 4.5005
R29839 VSS.n2494 VSS.n2362 4.5005
R29840 VSS.n2497 VSS.n2362 4.5005
R29841 VSS.n2499 VSS.n2362 4.5005
R29842 VSS.n2500 VSS.n2362 4.5005
R29843 VSS.n2502 VSS.n2362 4.5005
R29844 VSS.n2505 VSS.n2362 4.5005
R29845 VSS.n2507 VSS.n2362 4.5005
R29846 VSS.n2508 VSS.n2362 4.5005
R29847 VSS.n2510 VSS.n2362 4.5005
R29848 VSS.n2513 VSS.n2362 4.5005
R29849 VSS.n2515 VSS.n2362 4.5005
R29850 VSS.n2516 VSS.n2362 4.5005
R29851 VSS.n2518 VSS.n2362 4.5005
R29852 VSS.n2521 VSS.n2362 4.5005
R29853 VSS.n2523 VSS.n2362 4.5005
R29854 VSS.n2524 VSS.n2362 4.5005
R29855 VSS.n2526 VSS.n2362 4.5005
R29856 VSS.n2529 VSS.n2362 4.5005
R29857 VSS.n2531 VSS.n2362 4.5005
R29858 VSS.n2532 VSS.n2362 4.5005
R29859 VSS.n2534 VSS.n2362 4.5005
R29860 VSS.n2537 VSS.n2362 4.5005
R29861 VSS.n2539 VSS.n2362 4.5005
R29862 VSS.n2540 VSS.n2362 4.5005
R29863 VSS.n2542 VSS.n2362 4.5005
R29864 VSS.n2545 VSS.n2362 4.5005
R29865 VSS.n2547 VSS.n2362 4.5005
R29866 VSS.n2548 VSS.n2362 4.5005
R29867 VSS.n2550 VSS.n2362 4.5005
R29868 VSS.n2553 VSS.n2362 4.5005
R29869 VSS.n2555 VSS.n2362 4.5005
R29870 VSS.n2556 VSS.n2362 4.5005
R29871 VSS.n2558 VSS.n2362 4.5005
R29872 VSS.n2561 VSS.n2362 4.5005
R29873 VSS.n2563 VSS.n2362 4.5005
R29874 VSS.n2564 VSS.n2362 4.5005
R29875 VSS.n2566 VSS.n2362 4.5005
R29876 VSS.n2569 VSS.n2362 4.5005
R29877 VSS.n2571 VSS.n2362 4.5005
R29878 VSS.n2572 VSS.n2362 4.5005
R29879 VSS.n2574 VSS.n2362 4.5005
R29880 VSS.n2577 VSS.n2362 4.5005
R29881 VSS.n2579 VSS.n2362 4.5005
R29882 VSS.n2580 VSS.n2362 4.5005
R29883 VSS.n2582 VSS.n2362 4.5005
R29884 VSS.n2585 VSS.n2362 4.5005
R29885 VSS.n2587 VSS.n2362 4.5005
R29886 VSS.n2588 VSS.n2362 4.5005
R29887 VSS.n2590 VSS.n2362 4.5005
R29888 VSS.n2593 VSS.n2362 4.5005
R29889 VSS.n2595 VSS.n2362 4.5005
R29890 VSS.n2596 VSS.n2362 4.5005
R29891 VSS.n2598 VSS.n2362 4.5005
R29892 VSS.n2601 VSS.n2362 4.5005
R29893 VSS.n2603 VSS.n2362 4.5005
R29894 VSS.n2604 VSS.n2362 4.5005
R29895 VSS.n2606 VSS.n2362 4.5005
R29896 VSS.n2609 VSS.n2362 4.5005
R29897 VSS.n2611 VSS.n2362 4.5005
R29898 VSS.n2612 VSS.n2362 4.5005
R29899 VSS.n2614 VSS.n2362 4.5005
R29900 VSS.n2617 VSS.n2362 4.5005
R29901 VSS.n2619 VSS.n2362 4.5005
R29902 VSS.n2620 VSS.n2362 4.5005
R29903 VSS.n2622 VSS.n2362 4.5005
R29904 VSS.n2625 VSS.n2362 4.5005
R29905 VSS.n2627 VSS.n2362 4.5005
R29906 VSS.n2628 VSS.n2362 4.5005
R29907 VSS.n2630 VSS.n2362 4.5005
R29908 VSS.n2633 VSS.n2362 4.5005
R29909 VSS.n2635 VSS.n2362 4.5005
R29910 VSS.n2636 VSS.n2362 4.5005
R29911 VSS.n2638 VSS.n2362 4.5005
R29912 VSS.n2640 VSS.n2362 4.5005
R29913 VSS.n2642 VSS.n2362 4.5005
R29914 VSS.n2643 VSS.n2362 4.5005
R29915 VSS.n2645 VSS.n2362 4.5005
R29916 VSS.n2648 VSS.n2362 4.5005
R29917 VSS.n2650 VSS.n2362 4.5005
R29918 VSS.n2651 VSS.n2362 4.5005
R29919 VSS.n2653 VSS.n2362 4.5005
R29920 VSS.n2656 VSS.n2362 4.5005
R29921 VSS.n2658 VSS.n2362 4.5005
R29922 VSS.n2659 VSS.n2362 4.5005
R29923 VSS.n2661 VSS.n2362 4.5005
R29924 VSS.n2664 VSS.n2362 4.5005
R29925 VSS.n2666 VSS.n2362 4.5005
R29926 VSS.n2667 VSS.n2362 4.5005
R29927 VSS.n2669 VSS.n2362 4.5005
R29928 VSS.n2672 VSS.n2362 4.5005
R29929 VSS.n2674 VSS.n2362 4.5005
R29930 VSS.n2675 VSS.n2362 4.5005
R29931 VSS.n2677 VSS.n2362 4.5005
R29932 VSS.n2680 VSS.n2362 4.5005
R29933 VSS.n2682 VSS.n2362 4.5005
R29934 VSS.n2683 VSS.n2362 4.5005
R29935 VSS.n2685 VSS.n2362 4.5005
R29936 VSS.n2688 VSS.n2362 4.5005
R29937 VSS.n2690 VSS.n2362 4.5005
R29938 VSS.n2691 VSS.n2362 4.5005
R29939 VSS.n2693 VSS.n2362 4.5005
R29940 VSS.n2696 VSS.n2362 4.5005
R29941 VSS.n2698 VSS.n2362 4.5005
R29942 VSS.n2699 VSS.n2362 4.5005
R29943 VSS.n2701 VSS.n2362 4.5005
R29944 VSS.n2704 VSS.n2362 4.5005
R29945 VSS.n2706 VSS.n2362 4.5005
R29946 VSS.n2707 VSS.n2362 4.5005
R29947 VSS.n2709 VSS.n2362 4.5005
R29948 VSS.n2712 VSS.n2362 4.5005
R29949 VSS.n2714 VSS.n2362 4.5005
R29950 VSS.n2715 VSS.n2362 4.5005
R29951 VSS.n2717 VSS.n2362 4.5005
R29952 VSS.n2720 VSS.n2362 4.5005
R29953 VSS.n2722 VSS.n2362 4.5005
R29954 VSS.n2723 VSS.n2362 4.5005
R29955 VSS.n2725 VSS.n2362 4.5005
R29956 VSS.n2793 VSS.n2362 4.5005
R29957 VSS.n2859 VSS.n2362 4.5005
R29958 VSS.n3051 VSS.n2470 4.5005
R29959 VSS.n2470 VSS.n2351 4.5005
R29960 VSS.n2483 VSS.n2470 4.5005
R29961 VSS.n2484 VSS.n2470 4.5005
R29962 VSS.n2486 VSS.n2470 4.5005
R29963 VSS.n2489 VSS.n2470 4.5005
R29964 VSS.n2491 VSS.n2470 4.5005
R29965 VSS.n2492 VSS.n2470 4.5005
R29966 VSS.n2494 VSS.n2470 4.5005
R29967 VSS.n2497 VSS.n2470 4.5005
R29968 VSS.n2499 VSS.n2470 4.5005
R29969 VSS.n2500 VSS.n2470 4.5005
R29970 VSS.n2502 VSS.n2470 4.5005
R29971 VSS.n2505 VSS.n2470 4.5005
R29972 VSS.n2507 VSS.n2470 4.5005
R29973 VSS.n2508 VSS.n2470 4.5005
R29974 VSS.n2510 VSS.n2470 4.5005
R29975 VSS.n2513 VSS.n2470 4.5005
R29976 VSS.n2515 VSS.n2470 4.5005
R29977 VSS.n2516 VSS.n2470 4.5005
R29978 VSS.n2518 VSS.n2470 4.5005
R29979 VSS.n2521 VSS.n2470 4.5005
R29980 VSS.n2523 VSS.n2470 4.5005
R29981 VSS.n2524 VSS.n2470 4.5005
R29982 VSS.n2526 VSS.n2470 4.5005
R29983 VSS.n2529 VSS.n2470 4.5005
R29984 VSS.n2531 VSS.n2470 4.5005
R29985 VSS.n2532 VSS.n2470 4.5005
R29986 VSS.n2534 VSS.n2470 4.5005
R29987 VSS.n2537 VSS.n2470 4.5005
R29988 VSS.n2539 VSS.n2470 4.5005
R29989 VSS.n2540 VSS.n2470 4.5005
R29990 VSS.n2542 VSS.n2470 4.5005
R29991 VSS.n2545 VSS.n2470 4.5005
R29992 VSS.n2547 VSS.n2470 4.5005
R29993 VSS.n2548 VSS.n2470 4.5005
R29994 VSS.n2550 VSS.n2470 4.5005
R29995 VSS.n2553 VSS.n2470 4.5005
R29996 VSS.n2555 VSS.n2470 4.5005
R29997 VSS.n2556 VSS.n2470 4.5005
R29998 VSS.n2558 VSS.n2470 4.5005
R29999 VSS.n2561 VSS.n2470 4.5005
R30000 VSS.n2563 VSS.n2470 4.5005
R30001 VSS.n2564 VSS.n2470 4.5005
R30002 VSS.n2566 VSS.n2470 4.5005
R30003 VSS.n2569 VSS.n2470 4.5005
R30004 VSS.n2571 VSS.n2470 4.5005
R30005 VSS.n2572 VSS.n2470 4.5005
R30006 VSS.n2574 VSS.n2470 4.5005
R30007 VSS.n2577 VSS.n2470 4.5005
R30008 VSS.n2579 VSS.n2470 4.5005
R30009 VSS.n2580 VSS.n2470 4.5005
R30010 VSS.n2582 VSS.n2470 4.5005
R30011 VSS.n2585 VSS.n2470 4.5005
R30012 VSS.n2587 VSS.n2470 4.5005
R30013 VSS.n2588 VSS.n2470 4.5005
R30014 VSS.n2590 VSS.n2470 4.5005
R30015 VSS.n2593 VSS.n2470 4.5005
R30016 VSS.n2595 VSS.n2470 4.5005
R30017 VSS.n2596 VSS.n2470 4.5005
R30018 VSS.n2598 VSS.n2470 4.5005
R30019 VSS.n2601 VSS.n2470 4.5005
R30020 VSS.n2603 VSS.n2470 4.5005
R30021 VSS.n2604 VSS.n2470 4.5005
R30022 VSS.n2606 VSS.n2470 4.5005
R30023 VSS.n2609 VSS.n2470 4.5005
R30024 VSS.n2611 VSS.n2470 4.5005
R30025 VSS.n2612 VSS.n2470 4.5005
R30026 VSS.n2614 VSS.n2470 4.5005
R30027 VSS.n2617 VSS.n2470 4.5005
R30028 VSS.n2619 VSS.n2470 4.5005
R30029 VSS.n2620 VSS.n2470 4.5005
R30030 VSS.n2622 VSS.n2470 4.5005
R30031 VSS.n2625 VSS.n2470 4.5005
R30032 VSS.n2627 VSS.n2470 4.5005
R30033 VSS.n2628 VSS.n2470 4.5005
R30034 VSS.n2630 VSS.n2470 4.5005
R30035 VSS.n2633 VSS.n2470 4.5005
R30036 VSS.n2635 VSS.n2470 4.5005
R30037 VSS.n2636 VSS.n2470 4.5005
R30038 VSS.n2638 VSS.n2470 4.5005
R30039 VSS.n2640 VSS.n2470 4.5005
R30040 VSS.n2642 VSS.n2470 4.5005
R30041 VSS.n2643 VSS.n2470 4.5005
R30042 VSS.n2645 VSS.n2470 4.5005
R30043 VSS.n2648 VSS.n2470 4.5005
R30044 VSS.n2650 VSS.n2470 4.5005
R30045 VSS.n2651 VSS.n2470 4.5005
R30046 VSS.n2653 VSS.n2470 4.5005
R30047 VSS.n2656 VSS.n2470 4.5005
R30048 VSS.n2658 VSS.n2470 4.5005
R30049 VSS.n2659 VSS.n2470 4.5005
R30050 VSS.n2661 VSS.n2470 4.5005
R30051 VSS.n2664 VSS.n2470 4.5005
R30052 VSS.n2666 VSS.n2470 4.5005
R30053 VSS.n2667 VSS.n2470 4.5005
R30054 VSS.n2669 VSS.n2470 4.5005
R30055 VSS.n2672 VSS.n2470 4.5005
R30056 VSS.n2674 VSS.n2470 4.5005
R30057 VSS.n2675 VSS.n2470 4.5005
R30058 VSS.n2677 VSS.n2470 4.5005
R30059 VSS.n2680 VSS.n2470 4.5005
R30060 VSS.n2682 VSS.n2470 4.5005
R30061 VSS.n2683 VSS.n2470 4.5005
R30062 VSS.n2685 VSS.n2470 4.5005
R30063 VSS.n2688 VSS.n2470 4.5005
R30064 VSS.n2690 VSS.n2470 4.5005
R30065 VSS.n2691 VSS.n2470 4.5005
R30066 VSS.n2693 VSS.n2470 4.5005
R30067 VSS.n2696 VSS.n2470 4.5005
R30068 VSS.n2698 VSS.n2470 4.5005
R30069 VSS.n2699 VSS.n2470 4.5005
R30070 VSS.n2701 VSS.n2470 4.5005
R30071 VSS.n2704 VSS.n2470 4.5005
R30072 VSS.n2706 VSS.n2470 4.5005
R30073 VSS.n2707 VSS.n2470 4.5005
R30074 VSS.n2709 VSS.n2470 4.5005
R30075 VSS.n2712 VSS.n2470 4.5005
R30076 VSS.n2714 VSS.n2470 4.5005
R30077 VSS.n2715 VSS.n2470 4.5005
R30078 VSS.n2717 VSS.n2470 4.5005
R30079 VSS.n2720 VSS.n2470 4.5005
R30080 VSS.n2722 VSS.n2470 4.5005
R30081 VSS.n2723 VSS.n2470 4.5005
R30082 VSS.n2725 VSS.n2470 4.5005
R30083 VSS.n2793 VSS.n2470 4.5005
R30084 VSS.n2859 VSS.n2470 4.5005
R30085 VSS.n3051 VSS.n2361 4.5005
R30086 VSS.n2361 VSS.n2351 4.5005
R30087 VSS.n2483 VSS.n2361 4.5005
R30088 VSS.n2484 VSS.n2361 4.5005
R30089 VSS.n2486 VSS.n2361 4.5005
R30090 VSS.n2489 VSS.n2361 4.5005
R30091 VSS.n2491 VSS.n2361 4.5005
R30092 VSS.n2492 VSS.n2361 4.5005
R30093 VSS.n2494 VSS.n2361 4.5005
R30094 VSS.n2497 VSS.n2361 4.5005
R30095 VSS.n2499 VSS.n2361 4.5005
R30096 VSS.n2500 VSS.n2361 4.5005
R30097 VSS.n2502 VSS.n2361 4.5005
R30098 VSS.n2505 VSS.n2361 4.5005
R30099 VSS.n2507 VSS.n2361 4.5005
R30100 VSS.n2508 VSS.n2361 4.5005
R30101 VSS.n2510 VSS.n2361 4.5005
R30102 VSS.n2513 VSS.n2361 4.5005
R30103 VSS.n2515 VSS.n2361 4.5005
R30104 VSS.n2516 VSS.n2361 4.5005
R30105 VSS.n2518 VSS.n2361 4.5005
R30106 VSS.n2521 VSS.n2361 4.5005
R30107 VSS.n2523 VSS.n2361 4.5005
R30108 VSS.n2524 VSS.n2361 4.5005
R30109 VSS.n2526 VSS.n2361 4.5005
R30110 VSS.n2529 VSS.n2361 4.5005
R30111 VSS.n2531 VSS.n2361 4.5005
R30112 VSS.n2532 VSS.n2361 4.5005
R30113 VSS.n2534 VSS.n2361 4.5005
R30114 VSS.n2537 VSS.n2361 4.5005
R30115 VSS.n2539 VSS.n2361 4.5005
R30116 VSS.n2540 VSS.n2361 4.5005
R30117 VSS.n2542 VSS.n2361 4.5005
R30118 VSS.n2545 VSS.n2361 4.5005
R30119 VSS.n2547 VSS.n2361 4.5005
R30120 VSS.n2548 VSS.n2361 4.5005
R30121 VSS.n2550 VSS.n2361 4.5005
R30122 VSS.n2553 VSS.n2361 4.5005
R30123 VSS.n2555 VSS.n2361 4.5005
R30124 VSS.n2556 VSS.n2361 4.5005
R30125 VSS.n2558 VSS.n2361 4.5005
R30126 VSS.n2561 VSS.n2361 4.5005
R30127 VSS.n2563 VSS.n2361 4.5005
R30128 VSS.n2564 VSS.n2361 4.5005
R30129 VSS.n2566 VSS.n2361 4.5005
R30130 VSS.n2569 VSS.n2361 4.5005
R30131 VSS.n2571 VSS.n2361 4.5005
R30132 VSS.n2572 VSS.n2361 4.5005
R30133 VSS.n2574 VSS.n2361 4.5005
R30134 VSS.n2577 VSS.n2361 4.5005
R30135 VSS.n2579 VSS.n2361 4.5005
R30136 VSS.n2580 VSS.n2361 4.5005
R30137 VSS.n2582 VSS.n2361 4.5005
R30138 VSS.n2585 VSS.n2361 4.5005
R30139 VSS.n2587 VSS.n2361 4.5005
R30140 VSS.n2588 VSS.n2361 4.5005
R30141 VSS.n2590 VSS.n2361 4.5005
R30142 VSS.n2593 VSS.n2361 4.5005
R30143 VSS.n2595 VSS.n2361 4.5005
R30144 VSS.n2596 VSS.n2361 4.5005
R30145 VSS.n2598 VSS.n2361 4.5005
R30146 VSS.n2601 VSS.n2361 4.5005
R30147 VSS.n2603 VSS.n2361 4.5005
R30148 VSS.n2604 VSS.n2361 4.5005
R30149 VSS.n2606 VSS.n2361 4.5005
R30150 VSS.n2609 VSS.n2361 4.5005
R30151 VSS.n2611 VSS.n2361 4.5005
R30152 VSS.n2612 VSS.n2361 4.5005
R30153 VSS.n2614 VSS.n2361 4.5005
R30154 VSS.n2617 VSS.n2361 4.5005
R30155 VSS.n2619 VSS.n2361 4.5005
R30156 VSS.n2620 VSS.n2361 4.5005
R30157 VSS.n2622 VSS.n2361 4.5005
R30158 VSS.n2625 VSS.n2361 4.5005
R30159 VSS.n2627 VSS.n2361 4.5005
R30160 VSS.n2628 VSS.n2361 4.5005
R30161 VSS.n2630 VSS.n2361 4.5005
R30162 VSS.n2633 VSS.n2361 4.5005
R30163 VSS.n2635 VSS.n2361 4.5005
R30164 VSS.n2636 VSS.n2361 4.5005
R30165 VSS.n2638 VSS.n2361 4.5005
R30166 VSS.n2640 VSS.n2361 4.5005
R30167 VSS.n2642 VSS.n2361 4.5005
R30168 VSS.n2643 VSS.n2361 4.5005
R30169 VSS.n2645 VSS.n2361 4.5005
R30170 VSS.n2648 VSS.n2361 4.5005
R30171 VSS.n2650 VSS.n2361 4.5005
R30172 VSS.n2651 VSS.n2361 4.5005
R30173 VSS.n2653 VSS.n2361 4.5005
R30174 VSS.n2656 VSS.n2361 4.5005
R30175 VSS.n2658 VSS.n2361 4.5005
R30176 VSS.n2659 VSS.n2361 4.5005
R30177 VSS.n2661 VSS.n2361 4.5005
R30178 VSS.n2664 VSS.n2361 4.5005
R30179 VSS.n2666 VSS.n2361 4.5005
R30180 VSS.n2667 VSS.n2361 4.5005
R30181 VSS.n2669 VSS.n2361 4.5005
R30182 VSS.n2672 VSS.n2361 4.5005
R30183 VSS.n2674 VSS.n2361 4.5005
R30184 VSS.n2675 VSS.n2361 4.5005
R30185 VSS.n2677 VSS.n2361 4.5005
R30186 VSS.n2680 VSS.n2361 4.5005
R30187 VSS.n2682 VSS.n2361 4.5005
R30188 VSS.n2683 VSS.n2361 4.5005
R30189 VSS.n2685 VSS.n2361 4.5005
R30190 VSS.n2688 VSS.n2361 4.5005
R30191 VSS.n2690 VSS.n2361 4.5005
R30192 VSS.n2691 VSS.n2361 4.5005
R30193 VSS.n2693 VSS.n2361 4.5005
R30194 VSS.n2696 VSS.n2361 4.5005
R30195 VSS.n2698 VSS.n2361 4.5005
R30196 VSS.n2699 VSS.n2361 4.5005
R30197 VSS.n2701 VSS.n2361 4.5005
R30198 VSS.n2704 VSS.n2361 4.5005
R30199 VSS.n2706 VSS.n2361 4.5005
R30200 VSS.n2707 VSS.n2361 4.5005
R30201 VSS.n2709 VSS.n2361 4.5005
R30202 VSS.n2712 VSS.n2361 4.5005
R30203 VSS.n2714 VSS.n2361 4.5005
R30204 VSS.n2715 VSS.n2361 4.5005
R30205 VSS.n2717 VSS.n2361 4.5005
R30206 VSS.n2720 VSS.n2361 4.5005
R30207 VSS.n2722 VSS.n2361 4.5005
R30208 VSS.n2723 VSS.n2361 4.5005
R30209 VSS.n2725 VSS.n2361 4.5005
R30210 VSS.n2793 VSS.n2361 4.5005
R30211 VSS.n2859 VSS.n2361 4.5005
R30212 VSS.n3051 VSS.n2471 4.5005
R30213 VSS.n2471 VSS.n2351 4.5005
R30214 VSS.n2483 VSS.n2471 4.5005
R30215 VSS.n2484 VSS.n2471 4.5005
R30216 VSS.n2486 VSS.n2471 4.5005
R30217 VSS.n2489 VSS.n2471 4.5005
R30218 VSS.n2491 VSS.n2471 4.5005
R30219 VSS.n2492 VSS.n2471 4.5005
R30220 VSS.n2494 VSS.n2471 4.5005
R30221 VSS.n2497 VSS.n2471 4.5005
R30222 VSS.n2499 VSS.n2471 4.5005
R30223 VSS.n2500 VSS.n2471 4.5005
R30224 VSS.n2502 VSS.n2471 4.5005
R30225 VSS.n2505 VSS.n2471 4.5005
R30226 VSS.n2507 VSS.n2471 4.5005
R30227 VSS.n2508 VSS.n2471 4.5005
R30228 VSS.n2510 VSS.n2471 4.5005
R30229 VSS.n2513 VSS.n2471 4.5005
R30230 VSS.n2515 VSS.n2471 4.5005
R30231 VSS.n2516 VSS.n2471 4.5005
R30232 VSS.n2518 VSS.n2471 4.5005
R30233 VSS.n2521 VSS.n2471 4.5005
R30234 VSS.n2523 VSS.n2471 4.5005
R30235 VSS.n2524 VSS.n2471 4.5005
R30236 VSS.n2526 VSS.n2471 4.5005
R30237 VSS.n2529 VSS.n2471 4.5005
R30238 VSS.n2531 VSS.n2471 4.5005
R30239 VSS.n2532 VSS.n2471 4.5005
R30240 VSS.n2534 VSS.n2471 4.5005
R30241 VSS.n2537 VSS.n2471 4.5005
R30242 VSS.n2539 VSS.n2471 4.5005
R30243 VSS.n2540 VSS.n2471 4.5005
R30244 VSS.n2542 VSS.n2471 4.5005
R30245 VSS.n2545 VSS.n2471 4.5005
R30246 VSS.n2547 VSS.n2471 4.5005
R30247 VSS.n2548 VSS.n2471 4.5005
R30248 VSS.n2550 VSS.n2471 4.5005
R30249 VSS.n2553 VSS.n2471 4.5005
R30250 VSS.n2555 VSS.n2471 4.5005
R30251 VSS.n2556 VSS.n2471 4.5005
R30252 VSS.n2558 VSS.n2471 4.5005
R30253 VSS.n2561 VSS.n2471 4.5005
R30254 VSS.n2563 VSS.n2471 4.5005
R30255 VSS.n2564 VSS.n2471 4.5005
R30256 VSS.n2566 VSS.n2471 4.5005
R30257 VSS.n2569 VSS.n2471 4.5005
R30258 VSS.n2571 VSS.n2471 4.5005
R30259 VSS.n2572 VSS.n2471 4.5005
R30260 VSS.n2574 VSS.n2471 4.5005
R30261 VSS.n2577 VSS.n2471 4.5005
R30262 VSS.n2579 VSS.n2471 4.5005
R30263 VSS.n2580 VSS.n2471 4.5005
R30264 VSS.n2582 VSS.n2471 4.5005
R30265 VSS.n2585 VSS.n2471 4.5005
R30266 VSS.n2587 VSS.n2471 4.5005
R30267 VSS.n2588 VSS.n2471 4.5005
R30268 VSS.n2590 VSS.n2471 4.5005
R30269 VSS.n2593 VSS.n2471 4.5005
R30270 VSS.n2595 VSS.n2471 4.5005
R30271 VSS.n2596 VSS.n2471 4.5005
R30272 VSS.n2598 VSS.n2471 4.5005
R30273 VSS.n2601 VSS.n2471 4.5005
R30274 VSS.n2603 VSS.n2471 4.5005
R30275 VSS.n2604 VSS.n2471 4.5005
R30276 VSS.n2606 VSS.n2471 4.5005
R30277 VSS.n2609 VSS.n2471 4.5005
R30278 VSS.n2611 VSS.n2471 4.5005
R30279 VSS.n2612 VSS.n2471 4.5005
R30280 VSS.n2614 VSS.n2471 4.5005
R30281 VSS.n2617 VSS.n2471 4.5005
R30282 VSS.n2619 VSS.n2471 4.5005
R30283 VSS.n2620 VSS.n2471 4.5005
R30284 VSS.n2622 VSS.n2471 4.5005
R30285 VSS.n2625 VSS.n2471 4.5005
R30286 VSS.n2627 VSS.n2471 4.5005
R30287 VSS.n2628 VSS.n2471 4.5005
R30288 VSS.n2630 VSS.n2471 4.5005
R30289 VSS.n2633 VSS.n2471 4.5005
R30290 VSS.n2635 VSS.n2471 4.5005
R30291 VSS.n2636 VSS.n2471 4.5005
R30292 VSS.n2638 VSS.n2471 4.5005
R30293 VSS.n2640 VSS.n2471 4.5005
R30294 VSS.n2642 VSS.n2471 4.5005
R30295 VSS.n2643 VSS.n2471 4.5005
R30296 VSS.n2645 VSS.n2471 4.5005
R30297 VSS.n2648 VSS.n2471 4.5005
R30298 VSS.n2650 VSS.n2471 4.5005
R30299 VSS.n2651 VSS.n2471 4.5005
R30300 VSS.n2653 VSS.n2471 4.5005
R30301 VSS.n2656 VSS.n2471 4.5005
R30302 VSS.n2658 VSS.n2471 4.5005
R30303 VSS.n2659 VSS.n2471 4.5005
R30304 VSS.n2661 VSS.n2471 4.5005
R30305 VSS.n2664 VSS.n2471 4.5005
R30306 VSS.n2666 VSS.n2471 4.5005
R30307 VSS.n2667 VSS.n2471 4.5005
R30308 VSS.n2669 VSS.n2471 4.5005
R30309 VSS.n2672 VSS.n2471 4.5005
R30310 VSS.n2674 VSS.n2471 4.5005
R30311 VSS.n2675 VSS.n2471 4.5005
R30312 VSS.n2677 VSS.n2471 4.5005
R30313 VSS.n2680 VSS.n2471 4.5005
R30314 VSS.n2682 VSS.n2471 4.5005
R30315 VSS.n2683 VSS.n2471 4.5005
R30316 VSS.n2685 VSS.n2471 4.5005
R30317 VSS.n2688 VSS.n2471 4.5005
R30318 VSS.n2690 VSS.n2471 4.5005
R30319 VSS.n2691 VSS.n2471 4.5005
R30320 VSS.n2693 VSS.n2471 4.5005
R30321 VSS.n2696 VSS.n2471 4.5005
R30322 VSS.n2698 VSS.n2471 4.5005
R30323 VSS.n2699 VSS.n2471 4.5005
R30324 VSS.n2701 VSS.n2471 4.5005
R30325 VSS.n2704 VSS.n2471 4.5005
R30326 VSS.n2706 VSS.n2471 4.5005
R30327 VSS.n2707 VSS.n2471 4.5005
R30328 VSS.n2709 VSS.n2471 4.5005
R30329 VSS.n2712 VSS.n2471 4.5005
R30330 VSS.n2714 VSS.n2471 4.5005
R30331 VSS.n2715 VSS.n2471 4.5005
R30332 VSS.n2717 VSS.n2471 4.5005
R30333 VSS.n2720 VSS.n2471 4.5005
R30334 VSS.n2722 VSS.n2471 4.5005
R30335 VSS.n2723 VSS.n2471 4.5005
R30336 VSS.n2725 VSS.n2471 4.5005
R30337 VSS.n2793 VSS.n2471 4.5005
R30338 VSS.n2859 VSS.n2471 4.5005
R30339 VSS.n3051 VSS.n2360 4.5005
R30340 VSS.n2360 VSS.n2351 4.5005
R30341 VSS.n2483 VSS.n2360 4.5005
R30342 VSS.n2484 VSS.n2360 4.5005
R30343 VSS.n2486 VSS.n2360 4.5005
R30344 VSS.n2489 VSS.n2360 4.5005
R30345 VSS.n2491 VSS.n2360 4.5005
R30346 VSS.n2492 VSS.n2360 4.5005
R30347 VSS.n2494 VSS.n2360 4.5005
R30348 VSS.n2497 VSS.n2360 4.5005
R30349 VSS.n2499 VSS.n2360 4.5005
R30350 VSS.n2500 VSS.n2360 4.5005
R30351 VSS.n2502 VSS.n2360 4.5005
R30352 VSS.n2505 VSS.n2360 4.5005
R30353 VSS.n2507 VSS.n2360 4.5005
R30354 VSS.n2508 VSS.n2360 4.5005
R30355 VSS.n2510 VSS.n2360 4.5005
R30356 VSS.n2513 VSS.n2360 4.5005
R30357 VSS.n2515 VSS.n2360 4.5005
R30358 VSS.n2516 VSS.n2360 4.5005
R30359 VSS.n2518 VSS.n2360 4.5005
R30360 VSS.n2521 VSS.n2360 4.5005
R30361 VSS.n2523 VSS.n2360 4.5005
R30362 VSS.n2524 VSS.n2360 4.5005
R30363 VSS.n2526 VSS.n2360 4.5005
R30364 VSS.n2529 VSS.n2360 4.5005
R30365 VSS.n2531 VSS.n2360 4.5005
R30366 VSS.n2532 VSS.n2360 4.5005
R30367 VSS.n2534 VSS.n2360 4.5005
R30368 VSS.n2537 VSS.n2360 4.5005
R30369 VSS.n2539 VSS.n2360 4.5005
R30370 VSS.n2540 VSS.n2360 4.5005
R30371 VSS.n2542 VSS.n2360 4.5005
R30372 VSS.n2545 VSS.n2360 4.5005
R30373 VSS.n2547 VSS.n2360 4.5005
R30374 VSS.n2548 VSS.n2360 4.5005
R30375 VSS.n2550 VSS.n2360 4.5005
R30376 VSS.n2553 VSS.n2360 4.5005
R30377 VSS.n2555 VSS.n2360 4.5005
R30378 VSS.n2556 VSS.n2360 4.5005
R30379 VSS.n2558 VSS.n2360 4.5005
R30380 VSS.n2561 VSS.n2360 4.5005
R30381 VSS.n2563 VSS.n2360 4.5005
R30382 VSS.n2564 VSS.n2360 4.5005
R30383 VSS.n2566 VSS.n2360 4.5005
R30384 VSS.n2569 VSS.n2360 4.5005
R30385 VSS.n2571 VSS.n2360 4.5005
R30386 VSS.n2572 VSS.n2360 4.5005
R30387 VSS.n2574 VSS.n2360 4.5005
R30388 VSS.n2577 VSS.n2360 4.5005
R30389 VSS.n2579 VSS.n2360 4.5005
R30390 VSS.n2580 VSS.n2360 4.5005
R30391 VSS.n2582 VSS.n2360 4.5005
R30392 VSS.n2585 VSS.n2360 4.5005
R30393 VSS.n2587 VSS.n2360 4.5005
R30394 VSS.n2588 VSS.n2360 4.5005
R30395 VSS.n2590 VSS.n2360 4.5005
R30396 VSS.n2593 VSS.n2360 4.5005
R30397 VSS.n2595 VSS.n2360 4.5005
R30398 VSS.n2596 VSS.n2360 4.5005
R30399 VSS.n2598 VSS.n2360 4.5005
R30400 VSS.n2601 VSS.n2360 4.5005
R30401 VSS.n2603 VSS.n2360 4.5005
R30402 VSS.n2604 VSS.n2360 4.5005
R30403 VSS.n2606 VSS.n2360 4.5005
R30404 VSS.n2609 VSS.n2360 4.5005
R30405 VSS.n2611 VSS.n2360 4.5005
R30406 VSS.n2612 VSS.n2360 4.5005
R30407 VSS.n2614 VSS.n2360 4.5005
R30408 VSS.n2617 VSS.n2360 4.5005
R30409 VSS.n2619 VSS.n2360 4.5005
R30410 VSS.n2620 VSS.n2360 4.5005
R30411 VSS.n2622 VSS.n2360 4.5005
R30412 VSS.n2625 VSS.n2360 4.5005
R30413 VSS.n2627 VSS.n2360 4.5005
R30414 VSS.n2628 VSS.n2360 4.5005
R30415 VSS.n2630 VSS.n2360 4.5005
R30416 VSS.n2633 VSS.n2360 4.5005
R30417 VSS.n2635 VSS.n2360 4.5005
R30418 VSS.n2636 VSS.n2360 4.5005
R30419 VSS.n2638 VSS.n2360 4.5005
R30420 VSS.n2640 VSS.n2360 4.5005
R30421 VSS.n2642 VSS.n2360 4.5005
R30422 VSS.n2643 VSS.n2360 4.5005
R30423 VSS.n2645 VSS.n2360 4.5005
R30424 VSS.n2648 VSS.n2360 4.5005
R30425 VSS.n2650 VSS.n2360 4.5005
R30426 VSS.n2651 VSS.n2360 4.5005
R30427 VSS.n2653 VSS.n2360 4.5005
R30428 VSS.n2656 VSS.n2360 4.5005
R30429 VSS.n2658 VSS.n2360 4.5005
R30430 VSS.n2659 VSS.n2360 4.5005
R30431 VSS.n2661 VSS.n2360 4.5005
R30432 VSS.n2664 VSS.n2360 4.5005
R30433 VSS.n2666 VSS.n2360 4.5005
R30434 VSS.n2667 VSS.n2360 4.5005
R30435 VSS.n2669 VSS.n2360 4.5005
R30436 VSS.n2672 VSS.n2360 4.5005
R30437 VSS.n2674 VSS.n2360 4.5005
R30438 VSS.n2675 VSS.n2360 4.5005
R30439 VSS.n2677 VSS.n2360 4.5005
R30440 VSS.n2680 VSS.n2360 4.5005
R30441 VSS.n2682 VSS.n2360 4.5005
R30442 VSS.n2683 VSS.n2360 4.5005
R30443 VSS.n2685 VSS.n2360 4.5005
R30444 VSS.n2688 VSS.n2360 4.5005
R30445 VSS.n2690 VSS.n2360 4.5005
R30446 VSS.n2691 VSS.n2360 4.5005
R30447 VSS.n2693 VSS.n2360 4.5005
R30448 VSS.n2696 VSS.n2360 4.5005
R30449 VSS.n2698 VSS.n2360 4.5005
R30450 VSS.n2699 VSS.n2360 4.5005
R30451 VSS.n2701 VSS.n2360 4.5005
R30452 VSS.n2704 VSS.n2360 4.5005
R30453 VSS.n2706 VSS.n2360 4.5005
R30454 VSS.n2707 VSS.n2360 4.5005
R30455 VSS.n2709 VSS.n2360 4.5005
R30456 VSS.n2712 VSS.n2360 4.5005
R30457 VSS.n2714 VSS.n2360 4.5005
R30458 VSS.n2715 VSS.n2360 4.5005
R30459 VSS.n2717 VSS.n2360 4.5005
R30460 VSS.n2720 VSS.n2360 4.5005
R30461 VSS.n2722 VSS.n2360 4.5005
R30462 VSS.n2723 VSS.n2360 4.5005
R30463 VSS.n2725 VSS.n2360 4.5005
R30464 VSS.n2793 VSS.n2360 4.5005
R30465 VSS.n2859 VSS.n2360 4.5005
R30466 VSS.n3051 VSS.n2472 4.5005
R30467 VSS.n2472 VSS.n2351 4.5005
R30468 VSS.n2483 VSS.n2472 4.5005
R30469 VSS.n2484 VSS.n2472 4.5005
R30470 VSS.n2486 VSS.n2472 4.5005
R30471 VSS.n2489 VSS.n2472 4.5005
R30472 VSS.n2491 VSS.n2472 4.5005
R30473 VSS.n2492 VSS.n2472 4.5005
R30474 VSS.n2494 VSS.n2472 4.5005
R30475 VSS.n2497 VSS.n2472 4.5005
R30476 VSS.n2499 VSS.n2472 4.5005
R30477 VSS.n2500 VSS.n2472 4.5005
R30478 VSS.n2502 VSS.n2472 4.5005
R30479 VSS.n2505 VSS.n2472 4.5005
R30480 VSS.n2507 VSS.n2472 4.5005
R30481 VSS.n2508 VSS.n2472 4.5005
R30482 VSS.n2510 VSS.n2472 4.5005
R30483 VSS.n2513 VSS.n2472 4.5005
R30484 VSS.n2515 VSS.n2472 4.5005
R30485 VSS.n2516 VSS.n2472 4.5005
R30486 VSS.n2518 VSS.n2472 4.5005
R30487 VSS.n2521 VSS.n2472 4.5005
R30488 VSS.n2523 VSS.n2472 4.5005
R30489 VSS.n2524 VSS.n2472 4.5005
R30490 VSS.n2526 VSS.n2472 4.5005
R30491 VSS.n2529 VSS.n2472 4.5005
R30492 VSS.n2531 VSS.n2472 4.5005
R30493 VSS.n2532 VSS.n2472 4.5005
R30494 VSS.n2534 VSS.n2472 4.5005
R30495 VSS.n2537 VSS.n2472 4.5005
R30496 VSS.n2539 VSS.n2472 4.5005
R30497 VSS.n2540 VSS.n2472 4.5005
R30498 VSS.n2542 VSS.n2472 4.5005
R30499 VSS.n2545 VSS.n2472 4.5005
R30500 VSS.n2547 VSS.n2472 4.5005
R30501 VSS.n2548 VSS.n2472 4.5005
R30502 VSS.n2550 VSS.n2472 4.5005
R30503 VSS.n2553 VSS.n2472 4.5005
R30504 VSS.n2555 VSS.n2472 4.5005
R30505 VSS.n2556 VSS.n2472 4.5005
R30506 VSS.n2558 VSS.n2472 4.5005
R30507 VSS.n2561 VSS.n2472 4.5005
R30508 VSS.n2563 VSS.n2472 4.5005
R30509 VSS.n2564 VSS.n2472 4.5005
R30510 VSS.n2566 VSS.n2472 4.5005
R30511 VSS.n2569 VSS.n2472 4.5005
R30512 VSS.n2571 VSS.n2472 4.5005
R30513 VSS.n2572 VSS.n2472 4.5005
R30514 VSS.n2574 VSS.n2472 4.5005
R30515 VSS.n2577 VSS.n2472 4.5005
R30516 VSS.n2579 VSS.n2472 4.5005
R30517 VSS.n2580 VSS.n2472 4.5005
R30518 VSS.n2582 VSS.n2472 4.5005
R30519 VSS.n2585 VSS.n2472 4.5005
R30520 VSS.n2587 VSS.n2472 4.5005
R30521 VSS.n2588 VSS.n2472 4.5005
R30522 VSS.n2590 VSS.n2472 4.5005
R30523 VSS.n2593 VSS.n2472 4.5005
R30524 VSS.n2595 VSS.n2472 4.5005
R30525 VSS.n2596 VSS.n2472 4.5005
R30526 VSS.n2598 VSS.n2472 4.5005
R30527 VSS.n2601 VSS.n2472 4.5005
R30528 VSS.n2603 VSS.n2472 4.5005
R30529 VSS.n2604 VSS.n2472 4.5005
R30530 VSS.n2606 VSS.n2472 4.5005
R30531 VSS.n2609 VSS.n2472 4.5005
R30532 VSS.n2611 VSS.n2472 4.5005
R30533 VSS.n2612 VSS.n2472 4.5005
R30534 VSS.n2614 VSS.n2472 4.5005
R30535 VSS.n2617 VSS.n2472 4.5005
R30536 VSS.n2619 VSS.n2472 4.5005
R30537 VSS.n2620 VSS.n2472 4.5005
R30538 VSS.n2622 VSS.n2472 4.5005
R30539 VSS.n2625 VSS.n2472 4.5005
R30540 VSS.n2627 VSS.n2472 4.5005
R30541 VSS.n2628 VSS.n2472 4.5005
R30542 VSS.n2630 VSS.n2472 4.5005
R30543 VSS.n2633 VSS.n2472 4.5005
R30544 VSS.n2635 VSS.n2472 4.5005
R30545 VSS.n2636 VSS.n2472 4.5005
R30546 VSS.n2638 VSS.n2472 4.5005
R30547 VSS.n2640 VSS.n2472 4.5005
R30548 VSS.n2642 VSS.n2472 4.5005
R30549 VSS.n2643 VSS.n2472 4.5005
R30550 VSS.n2645 VSS.n2472 4.5005
R30551 VSS.n2648 VSS.n2472 4.5005
R30552 VSS.n2650 VSS.n2472 4.5005
R30553 VSS.n2651 VSS.n2472 4.5005
R30554 VSS.n2653 VSS.n2472 4.5005
R30555 VSS.n2656 VSS.n2472 4.5005
R30556 VSS.n2658 VSS.n2472 4.5005
R30557 VSS.n2659 VSS.n2472 4.5005
R30558 VSS.n2661 VSS.n2472 4.5005
R30559 VSS.n2664 VSS.n2472 4.5005
R30560 VSS.n2666 VSS.n2472 4.5005
R30561 VSS.n2667 VSS.n2472 4.5005
R30562 VSS.n2669 VSS.n2472 4.5005
R30563 VSS.n2672 VSS.n2472 4.5005
R30564 VSS.n2674 VSS.n2472 4.5005
R30565 VSS.n2675 VSS.n2472 4.5005
R30566 VSS.n2677 VSS.n2472 4.5005
R30567 VSS.n2680 VSS.n2472 4.5005
R30568 VSS.n2682 VSS.n2472 4.5005
R30569 VSS.n2683 VSS.n2472 4.5005
R30570 VSS.n2685 VSS.n2472 4.5005
R30571 VSS.n2688 VSS.n2472 4.5005
R30572 VSS.n2690 VSS.n2472 4.5005
R30573 VSS.n2691 VSS.n2472 4.5005
R30574 VSS.n2693 VSS.n2472 4.5005
R30575 VSS.n2696 VSS.n2472 4.5005
R30576 VSS.n2698 VSS.n2472 4.5005
R30577 VSS.n2699 VSS.n2472 4.5005
R30578 VSS.n2701 VSS.n2472 4.5005
R30579 VSS.n2704 VSS.n2472 4.5005
R30580 VSS.n2706 VSS.n2472 4.5005
R30581 VSS.n2707 VSS.n2472 4.5005
R30582 VSS.n2709 VSS.n2472 4.5005
R30583 VSS.n2712 VSS.n2472 4.5005
R30584 VSS.n2714 VSS.n2472 4.5005
R30585 VSS.n2715 VSS.n2472 4.5005
R30586 VSS.n2717 VSS.n2472 4.5005
R30587 VSS.n2720 VSS.n2472 4.5005
R30588 VSS.n2722 VSS.n2472 4.5005
R30589 VSS.n2723 VSS.n2472 4.5005
R30590 VSS.n2725 VSS.n2472 4.5005
R30591 VSS.n2793 VSS.n2472 4.5005
R30592 VSS.n2859 VSS.n2472 4.5005
R30593 VSS.n3051 VSS.n2359 4.5005
R30594 VSS.n2359 VSS.n2351 4.5005
R30595 VSS.n2483 VSS.n2359 4.5005
R30596 VSS.n2484 VSS.n2359 4.5005
R30597 VSS.n2486 VSS.n2359 4.5005
R30598 VSS.n2489 VSS.n2359 4.5005
R30599 VSS.n2491 VSS.n2359 4.5005
R30600 VSS.n2492 VSS.n2359 4.5005
R30601 VSS.n2494 VSS.n2359 4.5005
R30602 VSS.n2497 VSS.n2359 4.5005
R30603 VSS.n2499 VSS.n2359 4.5005
R30604 VSS.n2500 VSS.n2359 4.5005
R30605 VSS.n2502 VSS.n2359 4.5005
R30606 VSS.n2505 VSS.n2359 4.5005
R30607 VSS.n2507 VSS.n2359 4.5005
R30608 VSS.n2508 VSS.n2359 4.5005
R30609 VSS.n2510 VSS.n2359 4.5005
R30610 VSS.n2513 VSS.n2359 4.5005
R30611 VSS.n2515 VSS.n2359 4.5005
R30612 VSS.n2516 VSS.n2359 4.5005
R30613 VSS.n2518 VSS.n2359 4.5005
R30614 VSS.n2521 VSS.n2359 4.5005
R30615 VSS.n2523 VSS.n2359 4.5005
R30616 VSS.n2524 VSS.n2359 4.5005
R30617 VSS.n2526 VSS.n2359 4.5005
R30618 VSS.n2529 VSS.n2359 4.5005
R30619 VSS.n2531 VSS.n2359 4.5005
R30620 VSS.n2532 VSS.n2359 4.5005
R30621 VSS.n2534 VSS.n2359 4.5005
R30622 VSS.n2537 VSS.n2359 4.5005
R30623 VSS.n2539 VSS.n2359 4.5005
R30624 VSS.n2540 VSS.n2359 4.5005
R30625 VSS.n2542 VSS.n2359 4.5005
R30626 VSS.n2545 VSS.n2359 4.5005
R30627 VSS.n2547 VSS.n2359 4.5005
R30628 VSS.n2548 VSS.n2359 4.5005
R30629 VSS.n2550 VSS.n2359 4.5005
R30630 VSS.n2553 VSS.n2359 4.5005
R30631 VSS.n2555 VSS.n2359 4.5005
R30632 VSS.n2556 VSS.n2359 4.5005
R30633 VSS.n2558 VSS.n2359 4.5005
R30634 VSS.n2561 VSS.n2359 4.5005
R30635 VSS.n2563 VSS.n2359 4.5005
R30636 VSS.n2564 VSS.n2359 4.5005
R30637 VSS.n2566 VSS.n2359 4.5005
R30638 VSS.n2569 VSS.n2359 4.5005
R30639 VSS.n2571 VSS.n2359 4.5005
R30640 VSS.n2572 VSS.n2359 4.5005
R30641 VSS.n2574 VSS.n2359 4.5005
R30642 VSS.n2577 VSS.n2359 4.5005
R30643 VSS.n2579 VSS.n2359 4.5005
R30644 VSS.n2580 VSS.n2359 4.5005
R30645 VSS.n2582 VSS.n2359 4.5005
R30646 VSS.n2585 VSS.n2359 4.5005
R30647 VSS.n2587 VSS.n2359 4.5005
R30648 VSS.n2588 VSS.n2359 4.5005
R30649 VSS.n2590 VSS.n2359 4.5005
R30650 VSS.n2593 VSS.n2359 4.5005
R30651 VSS.n2595 VSS.n2359 4.5005
R30652 VSS.n2596 VSS.n2359 4.5005
R30653 VSS.n2598 VSS.n2359 4.5005
R30654 VSS.n2601 VSS.n2359 4.5005
R30655 VSS.n2603 VSS.n2359 4.5005
R30656 VSS.n2604 VSS.n2359 4.5005
R30657 VSS.n2606 VSS.n2359 4.5005
R30658 VSS.n2609 VSS.n2359 4.5005
R30659 VSS.n2611 VSS.n2359 4.5005
R30660 VSS.n2612 VSS.n2359 4.5005
R30661 VSS.n2614 VSS.n2359 4.5005
R30662 VSS.n2617 VSS.n2359 4.5005
R30663 VSS.n2619 VSS.n2359 4.5005
R30664 VSS.n2620 VSS.n2359 4.5005
R30665 VSS.n2622 VSS.n2359 4.5005
R30666 VSS.n2625 VSS.n2359 4.5005
R30667 VSS.n2627 VSS.n2359 4.5005
R30668 VSS.n2628 VSS.n2359 4.5005
R30669 VSS.n2630 VSS.n2359 4.5005
R30670 VSS.n2633 VSS.n2359 4.5005
R30671 VSS.n2635 VSS.n2359 4.5005
R30672 VSS.n2636 VSS.n2359 4.5005
R30673 VSS.n2638 VSS.n2359 4.5005
R30674 VSS.n2640 VSS.n2359 4.5005
R30675 VSS.n2642 VSS.n2359 4.5005
R30676 VSS.n2643 VSS.n2359 4.5005
R30677 VSS.n2645 VSS.n2359 4.5005
R30678 VSS.n2648 VSS.n2359 4.5005
R30679 VSS.n2650 VSS.n2359 4.5005
R30680 VSS.n2651 VSS.n2359 4.5005
R30681 VSS.n2653 VSS.n2359 4.5005
R30682 VSS.n2656 VSS.n2359 4.5005
R30683 VSS.n2658 VSS.n2359 4.5005
R30684 VSS.n2659 VSS.n2359 4.5005
R30685 VSS.n2661 VSS.n2359 4.5005
R30686 VSS.n2664 VSS.n2359 4.5005
R30687 VSS.n2666 VSS.n2359 4.5005
R30688 VSS.n2667 VSS.n2359 4.5005
R30689 VSS.n2669 VSS.n2359 4.5005
R30690 VSS.n2672 VSS.n2359 4.5005
R30691 VSS.n2674 VSS.n2359 4.5005
R30692 VSS.n2675 VSS.n2359 4.5005
R30693 VSS.n2677 VSS.n2359 4.5005
R30694 VSS.n2680 VSS.n2359 4.5005
R30695 VSS.n2682 VSS.n2359 4.5005
R30696 VSS.n2683 VSS.n2359 4.5005
R30697 VSS.n2685 VSS.n2359 4.5005
R30698 VSS.n2688 VSS.n2359 4.5005
R30699 VSS.n2690 VSS.n2359 4.5005
R30700 VSS.n2691 VSS.n2359 4.5005
R30701 VSS.n2693 VSS.n2359 4.5005
R30702 VSS.n2696 VSS.n2359 4.5005
R30703 VSS.n2698 VSS.n2359 4.5005
R30704 VSS.n2699 VSS.n2359 4.5005
R30705 VSS.n2701 VSS.n2359 4.5005
R30706 VSS.n2704 VSS.n2359 4.5005
R30707 VSS.n2706 VSS.n2359 4.5005
R30708 VSS.n2707 VSS.n2359 4.5005
R30709 VSS.n2709 VSS.n2359 4.5005
R30710 VSS.n2712 VSS.n2359 4.5005
R30711 VSS.n2714 VSS.n2359 4.5005
R30712 VSS.n2715 VSS.n2359 4.5005
R30713 VSS.n2717 VSS.n2359 4.5005
R30714 VSS.n2720 VSS.n2359 4.5005
R30715 VSS.n2722 VSS.n2359 4.5005
R30716 VSS.n2723 VSS.n2359 4.5005
R30717 VSS.n2725 VSS.n2359 4.5005
R30718 VSS.n2793 VSS.n2359 4.5005
R30719 VSS.n2859 VSS.n2359 4.5005
R30720 VSS.n3051 VSS.n2473 4.5005
R30721 VSS.n2473 VSS.n2351 4.5005
R30722 VSS.n2483 VSS.n2473 4.5005
R30723 VSS.n2484 VSS.n2473 4.5005
R30724 VSS.n2486 VSS.n2473 4.5005
R30725 VSS.n2489 VSS.n2473 4.5005
R30726 VSS.n2491 VSS.n2473 4.5005
R30727 VSS.n2492 VSS.n2473 4.5005
R30728 VSS.n2494 VSS.n2473 4.5005
R30729 VSS.n2497 VSS.n2473 4.5005
R30730 VSS.n2499 VSS.n2473 4.5005
R30731 VSS.n2500 VSS.n2473 4.5005
R30732 VSS.n2502 VSS.n2473 4.5005
R30733 VSS.n2505 VSS.n2473 4.5005
R30734 VSS.n2507 VSS.n2473 4.5005
R30735 VSS.n2508 VSS.n2473 4.5005
R30736 VSS.n2510 VSS.n2473 4.5005
R30737 VSS.n2513 VSS.n2473 4.5005
R30738 VSS.n2515 VSS.n2473 4.5005
R30739 VSS.n2516 VSS.n2473 4.5005
R30740 VSS.n2518 VSS.n2473 4.5005
R30741 VSS.n2521 VSS.n2473 4.5005
R30742 VSS.n2523 VSS.n2473 4.5005
R30743 VSS.n2524 VSS.n2473 4.5005
R30744 VSS.n2526 VSS.n2473 4.5005
R30745 VSS.n2529 VSS.n2473 4.5005
R30746 VSS.n2531 VSS.n2473 4.5005
R30747 VSS.n2532 VSS.n2473 4.5005
R30748 VSS.n2534 VSS.n2473 4.5005
R30749 VSS.n2537 VSS.n2473 4.5005
R30750 VSS.n2539 VSS.n2473 4.5005
R30751 VSS.n2540 VSS.n2473 4.5005
R30752 VSS.n2542 VSS.n2473 4.5005
R30753 VSS.n2545 VSS.n2473 4.5005
R30754 VSS.n2547 VSS.n2473 4.5005
R30755 VSS.n2548 VSS.n2473 4.5005
R30756 VSS.n2550 VSS.n2473 4.5005
R30757 VSS.n2553 VSS.n2473 4.5005
R30758 VSS.n2555 VSS.n2473 4.5005
R30759 VSS.n2556 VSS.n2473 4.5005
R30760 VSS.n2558 VSS.n2473 4.5005
R30761 VSS.n2561 VSS.n2473 4.5005
R30762 VSS.n2563 VSS.n2473 4.5005
R30763 VSS.n2564 VSS.n2473 4.5005
R30764 VSS.n2566 VSS.n2473 4.5005
R30765 VSS.n2569 VSS.n2473 4.5005
R30766 VSS.n2571 VSS.n2473 4.5005
R30767 VSS.n2572 VSS.n2473 4.5005
R30768 VSS.n2574 VSS.n2473 4.5005
R30769 VSS.n2577 VSS.n2473 4.5005
R30770 VSS.n2579 VSS.n2473 4.5005
R30771 VSS.n2580 VSS.n2473 4.5005
R30772 VSS.n2582 VSS.n2473 4.5005
R30773 VSS.n2585 VSS.n2473 4.5005
R30774 VSS.n2587 VSS.n2473 4.5005
R30775 VSS.n2588 VSS.n2473 4.5005
R30776 VSS.n2590 VSS.n2473 4.5005
R30777 VSS.n2593 VSS.n2473 4.5005
R30778 VSS.n2595 VSS.n2473 4.5005
R30779 VSS.n2596 VSS.n2473 4.5005
R30780 VSS.n2598 VSS.n2473 4.5005
R30781 VSS.n2601 VSS.n2473 4.5005
R30782 VSS.n2603 VSS.n2473 4.5005
R30783 VSS.n2604 VSS.n2473 4.5005
R30784 VSS.n2606 VSS.n2473 4.5005
R30785 VSS.n2609 VSS.n2473 4.5005
R30786 VSS.n2611 VSS.n2473 4.5005
R30787 VSS.n2612 VSS.n2473 4.5005
R30788 VSS.n2614 VSS.n2473 4.5005
R30789 VSS.n2617 VSS.n2473 4.5005
R30790 VSS.n2619 VSS.n2473 4.5005
R30791 VSS.n2620 VSS.n2473 4.5005
R30792 VSS.n2622 VSS.n2473 4.5005
R30793 VSS.n2625 VSS.n2473 4.5005
R30794 VSS.n2627 VSS.n2473 4.5005
R30795 VSS.n2628 VSS.n2473 4.5005
R30796 VSS.n2630 VSS.n2473 4.5005
R30797 VSS.n2633 VSS.n2473 4.5005
R30798 VSS.n2635 VSS.n2473 4.5005
R30799 VSS.n2636 VSS.n2473 4.5005
R30800 VSS.n2638 VSS.n2473 4.5005
R30801 VSS.n2640 VSS.n2473 4.5005
R30802 VSS.n2642 VSS.n2473 4.5005
R30803 VSS.n2643 VSS.n2473 4.5005
R30804 VSS.n2645 VSS.n2473 4.5005
R30805 VSS.n2648 VSS.n2473 4.5005
R30806 VSS.n2650 VSS.n2473 4.5005
R30807 VSS.n2651 VSS.n2473 4.5005
R30808 VSS.n2653 VSS.n2473 4.5005
R30809 VSS.n2656 VSS.n2473 4.5005
R30810 VSS.n2658 VSS.n2473 4.5005
R30811 VSS.n2659 VSS.n2473 4.5005
R30812 VSS.n2661 VSS.n2473 4.5005
R30813 VSS.n2664 VSS.n2473 4.5005
R30814 VSS.n2666 VSS.n2473 4.5005
R30815 VSS.n2667 VSS.n2473 4.5005
R30816 VSS.n2669 VSS.n2473 4.5005
R30817 VSS.n2672 VSS.n2473 4.5005
R30818 VSS.n2674 VSS.n2473 4.5005
R30819 VSS.n2675 VSS.n2473 4.5005
R30820 VSS.n2677 VSS.n2473 4.5005
R30821 VSS.n2680 VSS.n2473 4.5005
R30822 VSS.n2682 VSS.n2473 4.5005
R30823 VSS.n2683 VSS.n2473 4.5005
R30824 VSS.n2685 VSS.n2473 4.5005
R30825 VSS.n2688 VSS.n2473 4.5005
R30826 VSS.n2690 VSS.n2473 4.5005
R30827 VSS.n2691 VSS.n2473 4.5005
R30828 VSS.n2693 VSS.n2473 4.5005
R30829 VSS.n2696 VSS.n2473 4.5005
R30830 VSS.n2698 VSS.n2473 4.5005
R30831 VSS.n2699 VSS.n2473 4.5005
R30832 VSS.n2701 VSS.n2473 4.5005
R30833 VSS.n2704 VSS.n2473 4.5005
R30834 VSS.n2706 VSS.n2473 4.5005
R30835 VSS.n2707 VSS.n2473 4.5005
R30836 VSS.n2709 VSS.n2473 4.5005
R30837 VSS.n2712 VSS.n2473 4.5005
R30838 VSS.n2714 VSS.n2473 4.5005
R30839 VSS.n2715 VSS.n2473 4.5005
R30840 VSS.n2717 VSS.n2473 4.5005
R30841 VSS.n2720 VSS.n2473 4.5005
R30842 VSS.n2722 VSS.n2473 4.5005
R30843 VSS.n2723 VSS.n2473 4.5005
R30844 VSS.n2725 VSS.n2473 4.5005
R30845 VSS.n2793 VSS.n2473 4.5005
R30846 VSS.n2859 VSS.n2473 4.5005
R30847 VSS.n3051 VSS.n2358 4.5005
R30848 VSS.n2358 VSS.n2351 4.5005
R30849 VSS.n2483 VSS.n2358 4.5005
R30850 VSS.n2484 VSS.n2358 4.5005
R30851 VSS.n2486 VSS.n2358 4.5005
R30852 VSS.n2489 VSS.n2358 4.5005
R30853 VSS.n2491 VSS.n2358 4.5005
R30854 VSS.n2492 VSS.n2358 4.5005
R30855 VSS.n2494 VSS.n2358 4.5005
R30856 VSS.n2497 VSS.n2358 4.5005
R30857 VSS.n2499 VSS.n2358 4.5005
R30858 VSS.n2500 VSS.n2358 4.5005
R30859 VSS.n2502 VSS.n2358 4.5005
R30860 VSS.n2505 VSS.n2358 4.5005
R30861 VSS.n2507 VSS.n2358 4.5005
R30862 VSS.n2508 VSS.n2358 4.5005
R30863 VSS.n2510 VSS.n2358 4.5005
R30864 VSS.n2513 VSS.n2358 4.5005
R30865 VSS.n2515 VSS.n2358 4.5005
R30866 VSS.n2516 VSS.n2358 4.5005
R30867 VSS.n2518 VSS.n2358 4.5005
R30868 VSS.n2521 VSS.n2358 4.5005
R30869 VSS.n2523 VSS.n2358 4.5005
R30870 VSS.n2524 VSS.n2358 4.5005
R30871 VSS.n2526 VSS.n2358 4.5005
R30872 VSS.n2529 VSS.n2358 4.5005
R30873 VSS.n2531 VSS.n2358 4.5005
R30874 VSS.n2532 VSS.n2358 4.5005
R30875 VSS.n2534 VSS.n2358 4.5005
R30876 VSS.n2537 VSS.n2358 4.5005
R30877 VSS.n2539 VSS.n2358 4.5005
R30878 VSS.n2540 VSS.n2358 4.5005
R30879 VSS.n2542 VSS.n2358 4.5005
R30880 VSS.n2545 VSS.n2358 4.5005
R30881 VSS.n2547 VSS.n2358 4.5005
R30882 VSS.n2548 VSS.n2358 4.5005
R30883 VSS.n2550 VSS.n2358 4.5005
R30884 VSS.n2553 VSS.n2358 4.5005
R30885 VSS.n2555 VSS.n2358 4.5005
R30886 VSS.n2556 VSS.n2358 4.5005
R30887 VSS.n2558 VSS.n2358 4.5005
R30888 VSS.n2561 VSS.n2358 4.5005
R30889 VSS.n2563 VSS.n2358 4.5005
R30890 VSS.n2564 VSS.n2358 4.5005
R30891 VSS.n2566 VSS.n2358 4.5005
R30892 VSS.n2569 VSS.n2358 4.5005
R30893 VSS.n2571 VSS.n2358 4.5005
R30894 VSS.n2572 VSS.n2358 4.5005
R30895 VSS.n2574 VSS.n2358 4.5005
R30896 VSS.n2577 VSS.n2358 4.5005
R30897 VSS.n2579 VSS.n2358 4.5005
R30898 VSS.n2580 VSS.n2358 4.5005
R30899 VSS.n2582 VSS.n2358 4.5005
R30900 VSS.n2585 VSS.n2358 4.5005
R30901 VSS.n2587 VSS.n2358 4.5005
R30902 VSS.n2588 VSS.n2358 4.5005
R30903 VSS.n2590 VSS.n2358 4.5005
R30904 VSS.n2593 VSS.n2358 4.5005
R30905 VSS.n2595 VSS.n2358 4.5005
R30906 VSS.n2596 VSS.n2358 4.5005
R30907 VSS.n2598 VSS.n2358 4.5005
R30908 VSS.n2601 VSS.n2358 4.5005
R30909 VSS.n2603 VSS.n2358 4.5005
R30910 VSS.n2604 VSS.n2358 4.5005
R30911 VSS.n2606 VSS.n2358 4.5005
R30912 VSS.n2609 VSS.n2358 4.5005
R30913 VSS.n2611 VSS.n2358 4.5005
R30914 VSS.n2612 VSS.n2358 4.5005
R30915 VSS.n2614 VSS.n2358 4.5005
R30916 VSS.n2617 VSS.n2358 4.5005
R30917 VSS.n2619 VSS.n2358 4.5005
R30918 VSS.n2620 VSS.n2358 4.5005
R30919 VSS.n2622 VSS.n2358 4.5005
R30920 VSS.n2625 VSS.n2358 4.5005
R30921 VSS.n2627 VSS.n2358 4.5005
R30922 VSS.n2628 VSS.n2358 4.5005
R30923 VSS.n2630 VSS.n2358 4.5005
R30924 VSS.n2633 VSS.n2358 4.5005
R30925 VSS.n2635 VSS.n2358 4.5005
R30926 VSS.n2636 VSS.n2358 4.5005
R30927 VSS.n2638 VSS.n2358 4.5005
R30928 VSS.n2640 VSS.n2358 4.5005
R30929 VSS.n2642 VSS.n2358 4.5005
R30930 VSS.n2643 VSS.n2358 4.5005
R30931 VSS.n2645 VSS.n2358 4.5005
R30932 VSS.n2648 VSS.n2358 4.5005
R30933 VSS.n2650 VSS.n2358 4.5005
R30934 VSS.n2651 VSS.n2358 4.5005
R30935 VSS.n2653 VSS.n2358 4.5005
R30936 VSS.n2656 VSS.n2358 4.5005
R30937 VSS.n2658 VSS.n2358 4.5005
R30938 VSS.n2659 VSS.n2358 4.5005
R30939 VSS.n2661 VSS.n2358 4.5005
R30940 VSS.n2664 VSS.n2358 4.5005
R30941 VSS.n2666 VSS.n2358 4.5005
R30942 VSS.n2667 VSS.n2358 4.5005
R30943 VSS.n2669 VSS.n2358 4.5005
R30944 VSS.n2672 VSS.n2358 4.5005
R30945 VSS.n2674 VSS.n2358 4.5005
R30946 VSS.n2675 VSS.n2358 4.5005
R30947 VSS.n2677 VSS.n2358 4.5005
R30948 VSS.n2680 VSS.n2358 4.5005
R30949 VSS.n2682 VSS.n2358 4.5005
R30950 VSS.n2683 VSS.n2358 4.5005
R30951 VSS.n2685 VSS.n2358 4.5005
R30952 VSS.n2688 VSS.n2358 4.5005
R30953 VSS.n2690 VSS.n2358 4.5005
R30954 VSS.n2691 VSS.n2358 4.5005
R30955 VSS.n2693 VSS.n2358 4.5005
R30956 VSS.n2696 VSS.n2358 4.5005
R30957 VSS.n2698 VSS.n2358 4.5005
R30958 VSS.n2699 VSS.n2358 4.5005
R30959 VSS.n2701 VSS.n2358 4.5005
R30960 VSS.n2704 VSS.n2358 4.5005
R30961 VSS.n2706 VSS.n2358 4.5005
R30962 VSS.n2707 VSS.n2358 4.5005
R30963 VSS.n2709 VSS.n2358 4.5005
R30964 VSS.n2712 VSS.n2358 4.5005
R30965 VSS.n2714 VSS.n2358 4.5005
R30966 VSS.n2715 VSS.n2358 4.5005
R30967 VSS.n2717 VSS.n2358 4.5005
R30968 VSS.n2720 VSS.n2358 4.5005
R30969 VSS.n2722 VSS.n2358 4.5005
R30970 VSS.n2723 VSS.n2358 4.5005
R30971 VSS.n2725 VSS.n2358 4.5005
R30972 VSS.n2793 VSS.n2358 4.5005
R30973 VSS.n2859 VSS.n2358 4.5005
R30974 VSS.n3051 VSS.n2474 4.5005
R30975 VSS.n2474 VSS.n2351 4.5005
R30976 VSS.n2483 VSS.n2474 4.5005
R30977 VSS.n2484 VSS.n2474 4.5005
R30978 VSS.n2486 VSS.n2474 4.5005
R30979 VSS.n2489 VSS.n2474 4.5005
R30980 VSS.n2491 VSS.n2474 4.5005
R30981 VSS.n2492 VSS.n2474 4.5005
R30982 VSS.n2494 VSS.n2474 4.5005
R30983 VSS.n2497 VSS.n2474 4.5005
R30984 VSS.n2499 VSS.n2474 4.5005
R30985 VSS.n2500 VSS.n2474 4.5005
R30986 VSS.n2502 VSS.n2474 4.5005
R30987 VSS.n2505 VSS.n2474 4.5005
R30988 VSS.n2507 VSS.n2474 4.5005
R30989 VSS.n2508 VSS.n2474 4.5005
R30990 VSS.n2510 VSS.n2474 4.5005
R30991 VSS.n2513 VSS.n2474 4.5005
R30992 VSS.n2515 VSS.n2474 4.5005
R30993 VSS.n2516 VSS.n2474 4.5005
R30994 VSS.n2518 VSS.n2474 4.5005
R30995 VSS.n2521 VSS.n2474 4.5005
R30996 VSS.n2523 VSS.n2474 4.5005
R30997 VSS.n2524 VSS.n2474 4.5005
R30998 VSS.n2526 VSS.n2474 4.5005
R30999 VSS.n2529 VSS.n2474 4.5005
R31000 VSS.n2531 VSS.n2474 4.5005
R31001 VSS.n2532 VSS.n2474 4.5005
R31002 VSS.n2534 VSS.n2474 4.5005
R31003 VSS.n2537 VSS.n2474 4.5005
R31004 VSS.n2539 VSS.n2474 4.5005
R31005 VSS.n2540 VSS.n2474 4.5005
R31006 VSS.n2542 VSS.n2474 4.5005
R31007 VSS.n2545 VSS.n2474 4.5005
R31008 VSS.n2547 VSS.n2474 4.5005
R31009 VSS.n2548 VSS.n2474 4.5005
R31010 VSS.n2550 VSS.n2474 4.5005
R31011 VSS.n2553 VSS.n2474 4.5005
R31012 VSS.n2555 VSS.n2474 4.5005
R31013 VSS.n2556 VSS.n2474 4.5005
R31014 VSS.n2558 VSS.n2474 4.5005
R31015 VSS.n2561 VSS.n2474 4.5005
R31016 VSS.n2563 VSS.n2474 4.5005
R31017 VSS.n2564 VSS.n2474 4.5005
R31018 VSS.n2566 VSS.n2474 4.5005
R31019 VSS.n2569 VSS.n2474 4.5005
R31020 VSS.n2571 VSS.n2474 4.5005
R31021 VSS.n2572 VSS.n2474 4.5005
R31022 VSS.n2574 VSS.n2474 4.5005
R31023 VSS.n2577 VSS.n2474 4.5005
R31024 VSS.n2579 VSS.n2474 4.5005
R31025 VSS.n2580 VSS.n2474 4.5005
R31026 VSS.n2582 VSS.n2474 4.5005
R31027 VSS.n2585 VSS.n2474 4.5005
R31028 VSS.n2587 VSS.n2474 4.5005
R31029 VSS.n2588 VSS.n2474 4.5005
R31030 VSS.n2590 VSS.n2474 4.5005
R31031 VSS.n2593 VSS.n2474 4.5005
R31032 VSS.n2595 VSS.n2474 4.5005
R31033 VSS.n2596 VSS.n2474 4.5005
R31034 VSS.n2598 VSS.n2474 4.5005
R31035 VSS.n2601 VSS.n2474 4.5005
R31036 VSS.n2603 VSS.n2474 4.5005
R31037 VSS.n2604 VSS.n2474 4.5005
R31038 VSS.n2606 VSS.n2474 4.5005
R31039 VSS.n2609 VSS.n2474 4.5005
R31040 VSS.n2611 VSS.n2474 4.5005
R31041 VSS.n2612 VSS.n2474 4.5005
R31042 VSS.n2614 VSS.n2474 4.5005
R31043 VSS.n2617 VSS.n2474 4.5005
R31044 VSS.n2619 VSS.n2474 4.5005
R31045 VSS.n2620 VSS.n2474 4.5005
R31046 VSS.n2622 VSS.n2474 4.5005
R31047 VSS.n2625 VSS.n2474 4.5005
R31048 VSS.n2627 VSS.n2474 4.5005
R31049 VSS.n2628 VSS.n2474 4.5005
R31050 VSS.n2630 VSS.n2474 4.5005
R31051 VSS.n2633 VSS.n2474 4.5005
R31052 VSS.n2635 VSS.n2474 4.5005
R31053 VSS.n2636 VSS.n2474 4.5005
R31054 VSS.n2638 VSS.n2474 4.5005
R31055 VSS.n2640 VSS.n2474 4.5005
R31056 VSS.n2642 VSS.n2474 4.5005
R31057 VSS.n2643 VSS.n2474 4.5005
R31058 VSS.n2645 VSS.n2474 4.5005
R31059 VSS.n2648 VSS.n2474 4.5005
R31060 VSS.n2650 VSS.n2474 4.5005
R31061 VSS.n2651 VSS.n2474 4.5005
R31062 VSS.n2653 VSS.n2474 4.5005
R31063 VSS.n2656 VSS.n2474 4.5005
R31064 VSS.n2658 VSS.n2474 4.5005
R31065 VSS.n2659 VSS.n2474 4.5005
R31066 VSS.n2661 VSS.n2474 4.5005
R31067 VSS.n2664 VSS.n2474 4.5005
R31068 VSS.n2666 VSS.n2474 4.5005
R31069 VSS.n2667 VSS.n2474 4.5005
R31070 VSS.n2669 VSS.n2474 4.5005
R31071 VSS.n2672 VSS.n2474 4.5005
R31072 VSS.n2674 VSS.n2474 4.5005
R31073 VSS.n2675 VSS.n2474 4.5005
R31074 VSS.n2677 VSS.n2474 4.5005
R31075 VSS.n2680 VSS.n2474 4.5005
R31076 VSS.n2682 VSS.n2474 4.5005
R31077 VSS.n2683 VSS.n2474 4.5005
R31078 VSS.n2685 VSS.n2474 4.5005
R31079 VSS.n2688 VSS.n2474 4.5005
R31080 VSS.n2690 VSS.n2474 4.5005
R31081 VSS.n2691 VSS.n2474 4.5005
R31082 VSS.n2693 VSS.n2474 4.5005
R31083 VSS.n2696 VSS.n2474 4.5005
R31084 VSS.n2698 VSS.n2474 4.5005
R31085 VSS.n2699 VSS.n2474 4.5005
R31086 VSS.n2701 VSS.n2474 4.5005
R31087 VSS.n2704 VSS.n2474 4.5005
R31088 VSS.n2706 VSS.n2474 4.5005
R31089 VSS.n2707 VSS.n2474 4.5005
R31090 VSS.n2709 VSS.n2474 4.5005
R31091 VSS.n2712 VSS.n2474 4.5005
R31092 VSS.n2714 VSS.n2474 4.5005
R31093 VSS.n2715 VSS.n2474 4.5005
R31094 VSS.n2717 VSS.n2474 4.5005
R31095 VSS.n2720 VSS.n2474 4.5005
R31096 VSS.n2722 VSS.n2474 4.5005
R31097 VSS.n2723 VSS.n2474 4.5005
R31098 VSS.n2725 VSS.n2474 4.5005
R31099 VSS.n2793 VSS.n2474 4.5005
R31100 VSS.n2859 VSS.n2474 4.5005
R31101 VSS.n3051 VSS.n2357 4.5005
R31102 VSS.n2357 VSS.n2351 4.5005
R31103 VSS.n2483 VSS.n2357 4.5005
R31104 VSS.n2484 VSS.n2357 4.5005
R31105 VSS.n2486 VSS.n2357 4.5005
R31106 VSS.n2489 VSS.n2357 4.5005
R31107 VSS.n2491 VSS.n2357 4.5005
R31108 VSS.n2492 VSS.n2357 4.5005
R31109 VSS.n2494 VSS.n2357 4.5005
R31110 VSS.n2497 VSS.n2357 4.5005
R31111 VSS.n2499 VSS.n2357 4.5005
R31112 VSS.n2500 VSS.n2357 4.5005
R31113 VSS.n2502 VSS.n2357 4.5005
R31114 VSS.n2505 VSS.n2357 4.5005
R31115 VSS.n2507 VSS.n2357 4.5005
R31116 VSS.n2508 VSS.n2357 4.5005
R31117 VSS.n2510 VSS.n2357 4.5005
R31118 VSS.n2513 VSS.n2357 4.5005
R31119 VSS.n2515 VSS.n2357 4.5005
R31120 VSS.n2516 VSS.n2357 4.5005
R31121 VSS.n2518 VSS.n2357 4.5005
R31122 VSS.n2521 VSS.n2357 4.5005
R31123 VSS.n2523 VSS.n2357 4.5005
R31124 VSS.n2524 VSS.n2357 4.5005
R31125 VSS.n2526 VSS.n2357 4.5005
R31126 VSS.n2529 VSS.n2357 4.5005
R31127 VSS.n2531 VSS.n2357 4.5005
R31128 VSS.n2532 VSS.n2357 4.5005
R31129 VSS.n2534 VSS.n2357 4.5005
R31130 VSS.n2537 VSS.n2357 4.5005
R31131 VSS.n2539 VSS.n2357 4.5005
R31132 VSS.n2540 VSS.n2357 4.5005
R31133 VSS.n2542 VSS.n2357 4.5005
R31134 VSS.n2545 VSS.n2357 4.5005
R31135 VSS.n2547 VSS.n2357 4.5005
R31136 VSS.n2548 VSS.n2357 4.5005
R31137 VSS.n2550 VSS.n2357 4.5005
R31138 VSS.n2553 VSS.n2357 4.5005
R31139 VSS.n2555 VSS.n2357 4.5005
R31140 VSS.n2556 VSS.n2357 4.5005
R31141 VSS.n2558 VSS.n2357 4.5005
R31142 VSS.n2561 VSS.n2357 4.5005
R31143 VSS.n2563 VSS.n2357 4.5005
R31144 VSS.n2564 VSS.n2357 4.5005
R31145 VSS.n2566 VSS.n2357 4.5005
R31146 VSS.n2569 VSS.n2357 4.5005
R31147 VSS.n2571 VSS.n2357 4.5005
R31148 VSS.n2572 VSS.n2357 4.5005
R31149 VSS.n2574 VSS.n2357 4.5005
R31150 VSS.n2577 VSS.n2357 4.5005
R31151 VSS.n2579 VSS.n2357 4.5005
R31152 VSS.n2580 VSS.n2357 4.5005
R31153 VSS.n2582 VSS.n2357 4.5005
R31154 VSS.n2585 VSS.n2357 4.5005
R31155 VSS.n2587 VSS.n2357 4.5005
R31156 VSS.n2588 VSS.n2357 4.5005
R31157 VSS.n2590 VSS.n2357 4.5005
R31158 VSS.n2593 VSS.n2357 4.5005
R31159 VSS.n2595 VSS.n2357 4.5005
R31160 VSS.n2596 VSS.n2357 4.5005
R31161 VSS.n2598 VSS.n2357 4.5005
R31162 VSS.n2601 VSS.n2357 4.5005
R31163 VSS.n2603 VSS.n2357 4.5005
R31164 VSS.n2604 VSS.n2357 4.5005
R31165 VSS.n2606 VSS.n2357 4.5005
R31166 VSS.n2609 VSS.n2357 4.5005
R31167 VSS.n2611 VSS.n2357 4.5005
R31168 VSS.n2612 VSS.n2357 4.5005
R31169 VSS.n2614 VSS.n2357 4.5005
R31170 VSS.n2617 VSS.n2357 4.5005
R31171 VSS.n2619 VSS.n2357 4.5005
R31172 VSS.n2620 VSS.n2357 4.5005
R31173 VSS.n2622 VSS.n2357 4.5005
R31174 VSS.n2625 VSS.n2357 4.5005
R31175 VSS.n2627 VSS.n2357 4.5005
R31176 VSS.n2628 VSS.n2357 4.5005
R31177 VSS.n2630 VSS.n2357 4.5005
R31178 VSS.n2633 VSS.n2357 4.5005
R31179 VSS.n2635 VSS.n2357 4.5005
R31180 VSS.n2636 VSS.n2357 4.5005
R31181 VSS.n2638 VSS.n2357 4.5005
R31182 VSS.n2640 VSS.n2357 4.5005
R31183 VSS.n2642 VSS.n2357 4.5005
R31184 VSS.n2643 VSS.n2357 4.5005
R31185 VSS.n2645 VSS.n2357 4.5005
R31186 VSS.n2648 VSS.n2357 4.5005
R31187 VSS.n2650 VSS.n2357 4.5005
R31188 VSS.n2651 VSS.n2357 4.5005
R31189 VSS.n2653 VSS.n2357 4.5005
R31190 VSS.n2656 VSS.n2357 4.5005
R31191 VSS.n2658 VSS.n2357 4.5005
R31192 VSS.n2659 VSS.n2357 4.5005
R31193 VSS.n2661 VSS.n2357 4.5005
R31194 VSS.n2664 VSS.n2357 4.5005
R31195 VSS.n2666 VSS.n2357 4.5005
R31196 VSS.n2667 VSS.n2357 4.5005
R31197 VSS.n2669 VSS.n2357 4.5005
R31198 VSS.n2672 VSS.n2357 4.5005
R31199 VSS.n2674 VSS.n2357 4.5005
R31200 VSS.n2675 VSS.n2357 4.5005
R31201 VSS.n2677 VSS.n2357 4.5005
R31202 VSS.n2680 VSS.n2357 4.5005
R31203 VSS.n2682 VSS.n2357 4.5005
R31204 VSS.n2683 VSS.n2357 4.5005
R31205 VSS.n2685 VSS.n2357 4.5005
R31206 VSS.n2688 VSS.n2357 4.5005
R31207 VSS.n2690 VSS.n2357 4.5005
R31208 VSS.n2691 VSS.n2357 4.5005
R31209 VSS.n2693 VSS.n2357 4.5005
R31210 VSS.n2696 VSS.n2357 4.5005
R31211 VSS.n2698 VSS.n2357 4.5005
R31212 VSS.n2699 VSS.n2357 4.5005
R31213 VSS.n2701 VSS.n2357 4.5005
R31214 VSS.n2704 VSS.n2357 4.5005
R31215 VSS.n2706 VSS.n2357 4.5005
R31216 VSS.n2707 VSS.n2357 4.5005
R31217 VSS.n2709 VSS.n2357 4.5005
R31218 VSS.n2712 VSS.n2357 4.5005
R31219 VSS.n2714 VSS.n2357 4.5005
R31220 VSS.n2715 VSS.n2357 4.5005
R31221 VSS.n2717 VSS.n2357 4.5005
R31222 VSS.n2720 VSS.n2357 4.5005
R31223 VSS.n2722 VSS.n2357 4.5005
R31224 VSS.n2723 VSS.n2357 4.5005
R31225 VSS.n2725 VSS.n2357 4.5005
R31226 VSS.n2793 VSS.n2357 4.5005
R31227 VSS.n2859 VSS.n2357 4.5005
R31228 VSS.n3051 VSS.n2475 4.5005
R31229 VSS.n2475 VSS.n2351 4.5005
R31230 VSS.n2483 VSS.n2475 4.5005
R31231 VSS.n2484 VSS.n2475 4.5005
R31232 VSS.n2486 VSS.n2475 4.5005
R31233 VSS.n2489 VSS.n2475 4.5005
R31234 VSS.n2491 VSS.n2475 4.5005
R31235 VSS.n2492 VSS.n2475 4.5005
R31236 VSS.n2494 VSS.n2475 4.5005
R31237 VSS.n2497 VSS.n2475 4.5005
R31238 VSS.n2499 VSS.n2475 4.5005
R31239 VSS.n2500 VSS.n2475 4.5005
R31240 VSS.n2502 VSS.n2475 4.5005
R31241 VSS.n2505 VSS.n2475 4.5005
R31242 VSS.n2507 VSS.n2475 4.5005
R31243 VSS.n2508 VSS.n2475 4.5005
R31244 VSS.n2510 VSS.n2475 4.5005
R31245 VSS.n2513 VSS.n2475 4.5005
R31246 VSS.n2515 VSS.n2475 4.5005
R31247 VSS.n2516 VSS.n2475 4.5005
R31248 VSS.n2518 VSS.n2475 4.5005
R31249 VSS.n2521 VSS.n2475 4.5005
R31250 VSS.n2523 VSS.n2475 4.5005
R31251 VSS.n2524 VSS.n2475 4.5005
R31252 VSS.n2526 VSS.n2475 4.5005
R31253 VSS.n2529 VSS.n2475 4.5005
R31254 VSS.n2531 VSS.n2475 4.5005
R31255 VSS.n2532 VSS.n2475 4.5005
R31256 VSS.n2534 VSS.n2475 4.5005
R31257 VSS.n2537 VSS.n2475 4.5005
R31258 VSS.n2539 VSS.n2475 4.5005
R31259 VSS.n2540 VSS.n2475 4.5005
R31260 VSS.n2542 VSS.n2475 4.5005
R31261 VSS.n2545 VSS.n2475 4.5005
R31262 VSS.n2547 VSS.n2475 4.5005
R31263 VSS.n2548 VSS.n2475 4.5005
R31264 VSS.n2550 VSS.n2475 4.5005
R31265 VSS.n2553 VSS.n2475 4.5005
R31266 VSS.n2555 VSS.n2475 4.5005
R31267 VSS.n2556 VSS.n2475 4.5005
R31268 VSS.n2558 VSS.n2475 4.5005
R31269 VSS.n2561 VSS.n2475 4.5005
R31270 VSS.n2563 VSS.n2475 4.5005
R31271 VSS.n2564 VSS.n2475 4.5005
R31272 VSS.n2566 VSS.n2475 4.5005
R31273 VSS.n2569 VSS.n2475 4.5005
R31274 VSS.n2571 VSS.n2475 4.5005
R31275 VSS.n2572 VSS.n2475 4.5005
R31276 VSS.n2574 VSS.n2475 4.5005
R31277 VSS.n2577 VSS.n2475 4.5005
R31278 VSS.n2579 VSS.n2475 4.5005
R31279 VSS.n2580 VSS.n2475 4.5005
R31280 VSS.n2582 VSS.n2475 4.5005
R31281 VSS.n2585 VSS.n2475 4.5005
R31282 VSS.n2587 VSS.n2475 4.5005
R31283 VSS.n2588 VSS.n2475 4.5005
R31284 VSS.n2590 VSS.n2475 4.5005
R31285 VSS.n2593 VSS.n2475 4.5005
R31286 VSS.n2595 VSS.n2475 4.5005
R31287 VSS.n2596 VSS.n2475 4.5005
R31288 VSS.n2598 VSS.n2475 4.5005
R31289 VSS.n2601 VSS.n2475 4.5005
R31290 VSS.n2603 VSS.n2475 4.5005
R31291 VSS.n2604 VSS.n2475 4.5005
R31292 VSS.n2606 VSS.n2475 4.5005
R31293 VSS.n2609 VSS.n2475 4.5005
R31294 VSS.n2611 VSS.n2475 4.5005
R31295 VSS.n2612 VSS.n2475 4.5005
R31296 VSS.n2614 VSS.n2475 4.5005
R31297 VSS.n2617 VSS.n2475 4.5005
R31298 VSS.n2619 VSS.n2475 4.5005
R31299 VSS.n2620 VSS.n2475 4.5005
R31300 VSS.n2622 VSS.n2475 4.5005
R31301 VSS.n2625 VSS.n2475 4.5005
R31302 VSS.n2627 VSS.n2475 4.5005
R31303 VSS.n2628 VSS.n2475 4.5005
R31304 VSS.n2630 VSS.n2475 4.5005
R31305 VSS.n2633 VSS.n2475 4.5005
R31306 VSS.n2635 VSS.n2475 4.5005
R31307 VSS.n2636 VSS.n2475 4.5005
R31308 VSS.n2638 VSS.n2475 4.5005
R31309 VSS.n2640 VSS.n2475 4.5005
R31310 VSS.n2642 VSS.n2475 4.5005
R31311 VSS.n2643 VSS.n2475 4.5005
R31312 VSS.n2645 VSS.n2475 4.5005
R31313 VSS.n2648 VSS.n2475 4.5005
R31314 VSS.n2650 VSS.n2475 4.5005
R31315 VSS.n2651 VSS.n2475 4.5005
R31316 VSS.n2653 VSS.n2475 4.5005
R31317 VSS.n2656 VSS.n2475 4.5005
R31318 VSS.n2658 VSS.n2475 4.5005
R31319 VSS.n2659 VSS.n2475 4.5005
R31320 VSS.n2661 VSS.n2475 4.5005
R31321 VSS.n2664 VSS.n2475 4.5005
R31322 VSS.n2666 VSS.n2475 4.5005
R31323 VSS.n2667 VSS.n2475 4.5005
R31324 VSS.n2669 VSS.n2475 4.5005
R31325 VSS.n2672 VSS.n2475 4.5005
R31326 VSS.n2674 VSS.n2475 4.5005
R31327 VSS.n2675 VSS.n2475 4.5005
R31328 VSS.n2677 VSS.n2475 4.5005
R31329 VSS.n2680 VSS.n2475 4.5005
R31330 VSS.n2682 VSS.n2475 4.5005
R31331 VSS.n2683 VSS.n2475 4.5005
R31332 VSS.n2685 VSS.n2475 4.5005
R31333 VSS.n2688 VSS.n2475 4.5005
R31334 VSS.n2690 VSS.n2475 4.5005
R31335 VSS.n2691 VSS.n2475 4.5005
R31336 VSS.n2693 VSS.n2475 4.5005
R31337 VSS.n2696 VSS.n2475 4.5005
R31338 VSS.n2698 VSS.n2475 4.5005
R31339 VSS.n2699 VSS.n2475 4.5005
R31340 VSS.n2701 VSS.n2475 4.5005
R31341 VSS.n2704 VSS.n2475 4.5005
R31342 VSS.n2706 VSS.n2475 4.5005
R31343 VSS.n2707 VSS.n2475 4.5005
R31344 VSS.n2709 VSS.n2475 4.5005
R31345 VSS.n2712 VSS.n2475 4.5005
R31346 VSS.n2714 VSS.n2475 4.5005
R31347 VSS.n2715 VSS.n2475 4.5005
R31348 VSS.n2717 VSS.n2475 4.5005
R31349 VSS.n2720 VSS.n2475 4.5005
R31350 VSS.n2722 VSS.n2475 4.5005
R31351 VSS.n2723 VSS.n2475 4.5005
R31352 VSS.n2725 VSS.n2475 4.5005
R31353 VSS.n2793 VSS.n2475 4.5005
R31354 VSS.n2859 VSS.n2475 4.5005
R31355 VSS.n3051 VSS.n2356 4.5005
R31356 VSS.n2356 VSS.n2351 4.5005
R31357 VSS.n2483 VSS.n2356 4.5005
R31358 VSS.n2484 VSS.n2356 4.5005
R31359 VSS.n2486 VSS.n2356 4.5005
R31360 VSS.n2489 VSS.n2356 4.5005
R31361 VSS.n2491 VSS.n2356 4.5005
R31362 VSS.n2492 VSS.n2356 4.5005
R31363 VSS.n2494 VSS.n2356 4.5005
R31364 VSS.n2497 VSS.n2356 4.5005
R31365 VSS.n2499 VSS.n2356 4.5005
R31366 VSS.n2500 VSS.n2356 4.5005
R31367 VSS.n2502 VSS.n2356 4.5005
R31368 VSS.n2505 VSS.n2356 4.5005
R31369 VSS.n2507 VSS.n2356 4.5005
R31370 VSS.n2508 VSS.n2356 4.5005
R31371 VSS.n2510 VSS.n2356 4.5005
R31372 VSS.n2513 VSS.n2356 4.5005
R31373 VSS.n2515 VSS.n2356 4.5005
R31374 VSS.n2516 VSS.n2356 4.5005
R31375 VSS.n2518 VSS.n2356 4.5005
R31376 VSS.n2521 VSS.n2356 4.5005
R31377 VSS.n2523 VSS.n2356 4.5005
R31378 VSS.n2524 VSS.n2356 4.5005
R31379 VSS.n2526 VSS.n2356 4.5005
R31380 VSS.n2529 VSS.n2356 4.5005
R31381 VSS.n2531 VSS.n2356 4.5005
R31382 VSS.n2532 VSS.n2356 4.5005
R31383 VSS.n2534 VSS.n2356 4.5005
R31384 VSS.n2537 VSS.n2356 4.5005
R31385 VSS.n2539 VSS.n2356 4.5005
R31386 VSS.n2540 VSS.n2356 4.5005
R31387 VSS.n2542 VSS.n2356 4.5005
R31388 VSS.n2545 VSS.n2356 4.5005
R31389 VSS.n2547 VSS.n2356 4.5005
R31390 VSS.n2548 VSS.n2356 4.5005
R31391 VSS.n2550 VSS.n2356 4.5005
R31392 VSS.n2553 VSS.n2356 4.5005
R31393 VSS.n2555 VSS.n2356 4.5005
R31394 VSS.n2556 VSS.n2356 4.5005
R31395 VSS.n2558 VSS.n2356 4.5005
R31396 VSS.n2561 VSS.n2356 4.5005
R31397 VSS.n2563 VSS.n2356 4.5005
R31398 VSS.n2564 VSS.n2356 4.5005
R31399 VSS.n2566 VSS.n2356 4.5005
R31400 VSS.n2569 VSS.n2356 4.5005
R31401 VSS.n2571 VSS.n2356 4.5005
R31402 VSS.n2572 VSS.n2356 4.5005
R31403 VSS.n2574 VSS.n2356 4.5005
R31404 VSS.n2577 VSS.n2356 4.5005
R31405 VSS.n2579 VSS.n2356 4.5005
R31406 VSS.n2580 VSS.n2356 4.5005
R31407 VSS.n2582 VSS.n2356 4.5005
R31408 VSS.n2585 VSS.n2356 4.5005
R31409 VSS.n2587 VSS.n2356 4.5005
R31410 VSS.n2588 VSS.n2356 4.5005
R31411 VSS.n2590 VSS.n2356 4.5005
R31412 VSS.n2593 VSS.n2356 4.5005
R31413 VSS.n2595 VSS.n2356 4.5005
R31414 VSS.n2596 VSS.n2356 4.5005
R31415 VSS.n2598 VSS.n2356 4.5005
R31416 VSS.n2601 VSS.n2356 4.5005
R31417 VSS.n2603 VSS.n2356 4.5005
R31418 VSS.n2604 VSS.n2356 4.5005
R31419 VSS.n2606 VSS.n2356 4.5005
R31420 VSS.n2609 VSS.n2356 4.5005
R31421 VSS.n2611 VSS.n2356 4.5005
R31422 VSS.n2612 VSS.n2356 4.5005
R31423 VSS.n2614 VSS.n2356 4.5005
R31424 VSS.n2617 VSS.n2356 4.5005
R31425 VSS.n2619 VSS.n2356 4.5005
R31426 VSS.n2620 VSS.n2356 4.5005
R31427 VSS.n2622 VSS.n2356 4.5005
R31428 VSS.n2625 VSS.n2356 4.5005
R31429 VSS.n2627 VSS.n2356 4.5005
R31430 VSS.n2628 VSS.n2356 4.5005
R31431 VSS.n2630 VSS.n2356 4.5005
R31432 VSS.n2633 VSS.n2356 4.5005
R31433 VSS.n2635 VSS.n2356 4.5005
R31434 VSS.n2636 VSS.n2356 4.5005
R31435 VSS.n2638 VSS.n2356 4.5005
R31436 VSS.n2640 VSS.n2356 4.5005
R31437 VSS.n2642 VSS.n2356 4.5005
R31438 VSS.n2643 VSS.n2356 4.5005
R31439 VSS.n2645 VSS.n2356 4.5005
R31440 VSS.n2648 VSS.n2356 4.5005
R31441 VSS.n2650 VSS.n2356 4.5005
R31442 VSS.n2651 VSS.n2356 4.5005
R31443 VSS.n2653 VSS.n2356 4.5005
R31444 VSS.n2656 VSS.n2356 4.5005
R31445 VSS.n2658 VSS.n2356 4.5005
R31446 VSS.n2659 VSS.n2356 4.5005
R31447 VSS.n2661 VSS.n2356 4.5005
R31448 VSS.n2664 VSS.n2356 4.5005
R31449 VSS.n2666 VSS.n2356 4.5005
R31450 VSS.n2667 VSS.n2356 4.5005
R31451 VSS.n2669 VSS.n2356 4.5005
R31452 VSS.n2672 VSS.n2356 4.5005
R31453 VSS.n2674 VSS.n2356 4.5005
R31454 VSS.n2675 VSS.n2356 4.5005
R31455 VSS.n2677 VSS.n2356 4.5005
R31456 VSS.n2680 VSS.n2356 4.5005
R31457 VSS.n2682 VSS.n2356 4.5005
R31458 VSS.n2683 VSS.n2356 4.5005
R31459 VSS.n2685 VSS.n2356 4.5005
R31460 VSS.n2688 VSS.n2356 4.5005
R31461 VSS.n2690 VSS.n2356 4.5005
R31462 VSS.n2691 VSS.n2356 4.5005
R31463 VSS.n2693 VSS.n2356 4.5005
R31464 VSS.n2696 VSS.n2356 4.5005
R31465 VSS.n2698 VSS.n2356 4.5005
R31466 VSS.n2699 VSS.n2356 4.5005
R31467 VSS.n2701 VSS.n2356 4.5005
R31468 VSS.n2704 VSS.n2356 4.5005
R31469 VSS.n2706 VSS.n2356 4.5005
R31470 VSS.n2707 VSS.n2356 4.5005
R31471 VSS.n2709 VSS.n2356 4.5005
R31472 VSS.n2712 VSS.n2356 4.5005
R31473 VSS.n2714 VSS.n2356 4.5005
R31474 VSS.n2715 VSS.n2356 4.5005
R31475 VSS.n2717 VSS.n2356 4.5005
R31476 VSS.n2720 VSS.n2356 4.5005
R31477 VSS.n2722 VSS.n2356 4.5005
R31478 VSS.n2723 VSS.n2356 4.5005
R31479 VSS.n2725 VSS.n2356 4.5005
R31480 VSS.n2793 VSS.n2356 4.5005
R31481 VSS.n2859 VSS.n2356 4.5005
R31482 VSS.n3051 VSS.n2476 4.5005
R31483 VSS.n2476 VSS.n2351 4.5005
R31484 VSS.n2483 VSS.n2476 4.5005
R31485 VSS.n2484 VSS.n2476 4.5005
R31486 VSS.n2486 VSS.n2476 4.5005
R31487 VSS.n2489 VSS.n2476 4.5005
R31488 VSS.n2491 VSS.n2476 4.5005
R31489 VSS.n2492 VSS.n2476 4.5005
R31490 VSS.n2494 VSS.n2476 4.5005
R31491 VSS.n2497 VSS.n2476 4.5005
R31492 VSS.n2499 VSS.n2476 4.5005
R31493 VSS.n2500 VSS.n2476 4.5005
R31494 VSS.n2502 VSS.n2476 4.5005
R31495 VSS.n2505 VSS.n2476 4.5005
R31496 VSS.n2507 VSS.n2476 4.5005
R31497 VSS.n2508 VSS.n2476 4.5005
R31498 VSS.n2510 VSS.n2476 4.5005
R31499 VSS.n2513 VSS.n2476 4.5005
R31500 VSS.n2515 VSS.n2476 4.5005
R31501 VSS.n2516 VSS.n2476 4.5005
R31502 VSS.n2518 VSS.n2476 4.5005
R31503 VSS.n2521 VSS.n2476 4.5005
R31504 VSS.n2523 VSS.n2476 4.5005
R31505 VSS.n2524 VSS.n2476 4.5005
R31506 VSS.n2526 VSS.n2476 4.5005
R31507 VSS.n2529 VSS.n2476 4.5005
R31508 VSS.n2531 VSS.n2476 4.5005
R31509 VSS.n2532 VSS.n2476 4.5005
R31510 VSS.n2534 VSS.n2476 4.5005
R31511 VSS.n2537 VSS.n2476 4.5005
R31512 VSS.n2539 VSS.n2476 4.5005
R31513 VSS.n2540 VSS.n2476 4.5005
R31514 VSS.n2542 VSS.n2476 4.5005
R31515 VSS.n2545 VSS.n2476 4.5005
R31516 VSS.n2547 VSS.n2476 4.5005
R31517 VSS.n2548 VSS.n2476 4.5005
R31518 VSS.n2550 VSS.n2476 4.5005
R31519 VSS.n2553 VSS.n2476 4.5005
R31520 VSS.n2555 VSS.n2476 4.5005
R31521 VSS.n2556 VSS.n2476 4.5005
R31522 VSS.n2558 VSS.n2476 4.5005
R31523 VSS.n2561 VSS.n2476 4.5005
R31524 VSS.n2563 VSS.n2476 4.5005
R31525 VSS.n2564 VSS.n2476 4.5005
R31526 VSS.n2566 VSS.n2476 4.5005
R31527 VSS.n2569 VSS.n2476 4.5005
R31528 VSS.n2571 VSS.n2476 4.5005
R31529 VSS.n2572 VSS.n2476 4.5005
R31530 VSS.n2574 VSS.n2476 4.5005
R31531 VSS.n2577 VSS.n2476 4.5005
R31532 VSS.n2579 VSS.n2476 4.5005
R31533 VSS.n2580 VSS.n2476 4.5005
R31534 VSS.n2582 VSS.n2476 4.5005
R31535 VSS.n2585 VSS.n2476 4.5005
R31536 VSS.n2587 VSS.n2476 4.5005
R31537 VSS.n2588 VSS.n2476 4.5005
R31538 VSS.n2590 VSS.n2476 4.5005
R31539 VSS.n2593 VSS.n2476 4.5005
R31540 VSS.n2595 VSS.n2476 4.5005
R31541 VSS.n2596 VSS.n2476 4.5005
R31542 VSS.n2598 VSS.n2476 4.5005
R31543 VSS.n2601 VSS.n2476 4.5005
R31544 VSS.n2603 VSS.n2476 4.5005
R31545 VSS.n2604 VSS.n2476 4.5005
R31546 VSS.n2606 VSS.n2476 4.5005
R31547 VSS.n2609 VSS.n2476 4.5005
R31548 VSS.n2611 VSS.n2476 4.5005
R31549 VSS.n2612 VSS.n2476 4.5005
R31550 VSS.n2614 VSS.n2476 4.5005
R31551 VSS.n2617 VSS.n2476 4.5005
R31552 VSS.n2619 VSS.n2476 4.5005
R31553 VSS.n2620 VSS.n2476 4.5005
R31554 VSS.n2622 VSS.n2476 4.5005
R31555 VSS.n2625 VSS.n2476 4.5005
R31556 VSS.n2627 VSS.n2476 4.5005
R31557 VSS.n2628 VSS.n2476 4.5005
R31558 VSS.n2630 VSS.n2476 4.5005
R31559 VSS.n2633 VSS.n2476 4.5005
R31560 VSS.n2635 VSS.n2476 4.5005
R31561 VSS.n2636 VSS.n2476 4.5005
R31562 VSS.n2638 VSS.n2476 4.5005
R31563 VSS.n2640 VSS.n2476 4.5005
R31564 VSS.n2642 VSS.n2476 4.5005
R31565 VSS.n2643 VSS.n2476 4.5005
R31566 VSS.n2645 VSS.n2476 4.5005
R31567 VSS.n2648 VSS.n2476 4.5005
R31568 VSS.n2650 VSS.n2476 4.5005
R31569 VSS.n2651 VSS.n2476 4.5005
R31570 VSS.n2653 VSS.n2476 4.5005
R31571 VSS.n2656 VSS.n2476 4.5005
R31572 VSS.n2658 VSS.n2476 4.5005
R31573 VSS.n2659 VSS.n2476 4.5005
R31574 VSS.n2661 VSS.n2476 4.5005
R31575 VSS.n2664 VSS.n2476 4.5005
R31576 VSS.n2666 VSS.n2476 4.5005
R31577 VSS.n2667 VSS.n2476 4.5005
R31578 VSS.n2669 VSS.n2476 4.5005
R31579 VSS.n2672 VSS.n2476 4.5005
R31580 VSS.n2674 VSS.n2476 4.5005
R31581 VSS.n2675 VSS.n2476 4.5005
R31582 VSS.n2677 VSS.n2476 4.5005
R31583 VSS.n2680 VSS.n2476 4.5005
R31584 VSS.n2682 VSS.n2476 4.5005
R31585 VSS.n2683 VSS.n2476 4.5005
R31586 VSS.n2685 VSS.n2476 4.5005
R31587 VSS.n2688 VSS.n2476 4.5005
R31588 VSS.n2690 VSS.n2476 4.5005
R31589 VSS.n2691 VSS.n2476 4.5005
R31590 VSS.n2693 VSS.n2476 4.5005
R31591 VSS.n2696 VSS.n2476 4.5005
R31592 VSS.n2698 VSS.n2476 4.5005
R31593 VSS.n2699 VSS.n2476 4.5005
R31594 VSS.n2701 VSS.n2476 4.5005
R31595 VSS.n2704 VSS.n2476 4.5005
R31596 VSS.n2706 VSS.n2476 4.5005
R31597 VSS.n2707 VSS.n2476 4.5005
R31598 VSS.n2709 VSS.n2476 4.5005
R31599 VSS.n2712 VSS.n2476 4.5005
R31600 VSS.n2714 VSS.n2476 4.5005
R31601 VSS.n2715 VSS.n2476 4.5005
R31602 VSS.n2717 VSS.n2476 4.5005
R31603 VSS.n2720 VSS.n2476 4.5005
R31604 VSS.n2722 VSS.n2476 4.5005
R31605 VSS.n2723 VSS.n2476 4.5005
R31606 VSS.n2725 VSS.n2476 4.5005
R31607 VSS.n2793 VSS.n2476 4.5005
R31608 VSS.n2859 VSS.n2476 4.5005
R31609 VSS.n3051 VSS.n2355 4.5005
R31610 VSS.n2355 VSS.n2351 4.5005
R31611 VSS.n2483 VSS.n2355 4.5005
R31612 VSS.n2484 VSS.n2355 4.5005
R31613 VSS.n2486 VSS.n2355 4.5005
R31614 VSS.n2489 VSS.n2355 4.5005
R31615 VSS.n2491 VSS.n2355 4.5005
R31616 VSS.n2492 VSS.n2355 4.5005
R31617 VSS.n2494 VSS.n2355 4.5005
R31618 VSS.n2497 VSS.n2355 4.5005
R31619 VSS.n2499 VSS.n2355 4.5005
R31620 VSS.n2500 VSS.n2355 4.5005
R31621 VSS.n2502 VSS.n2355 4.5005
R31622 VSS.n2505 VSS.n2355 4.5005
R31623 VSS.n2507 VSS.n2355 4.5005
R31624 VSS.n2508 VSS.n2355 4.5005
R31625 VSS.n2510 VSS.n2355 4.5005
R31626 VSS.n2513 VSS.n2355 4.5005
R31627 VSS.n2515 VSS.n2355 4.5005
R31628 VSS.n2516 VSS.n2355 4.5005
R31629 VSS.n2518 VSS.n2355 4.5005
R31630 VSS.n2521 VSS.n2355 4.5005
R31631 VSS.n2523 VSS.n2355 4.5005
R31632 VSS.n2524 VSS.n2355 4.5005
R31633 VSS.n2526 VSS.n2355 4.5005
R31634 VSS.n2529 VSS.n2355 4.5005
R31635 VSS.n2531 VSS.n2355 4.5005
R31636 VSS.n2532 VSS.n2355 4.5005
R31637 VSS.n2534 VSS.n2355 4.5005
R31638 VSS.n2537 VSS.n2355 4.5005
R31639 VSS.n2539 VSS.n2355 4.5005
R31640 VSS.n2540 VSS.n2355 4.5005
R31641 VSS.n2542 VSS.n2355 4.5005
R31642 VSS.n2545 VSS.n2355 4.5005
R31643 VSS.n2547 VSS.n2355 4.5005
R31644 VSS.n2548 VSS.n2355 4.5005
R31645 VSS.n2550 VSS.n2355 4.5005
R31646 VSS.n2553 VSS.n2355 4.5005
R31647 VSS.n2555 VSS.n2355 4.5005
R31648 VSS.n2556 VSS.n2355 4.5005
R31649 VSS.n2558 VSS.n2355 4.5005
R31650 VSS.n2561 VSS.n2355 4.5005
R31651 VSS.n2563 VSS.n2355 4.5005
R31652 VSS.n2564 VSS.n2355 4.5005
R31653 VSS.n2566 VSS.n2355 4.5005
R31654 VSS.n2569 VSS.n2355 4.5005
R31655 VSS.n2571 VSS.n2355 4.5005
R31656 VSS.n2572 VSS.n2355 4.5005
R31657 VSS.n2574 VSS.n2355 4.5005
R31658 VSS.n2577 VSS.n2355 4.5005
R31659 VSS.n2579 VSS.n2355 4.5005
R31660 VSS.n2580 VSS.n2355 4.5005
R31661 VSS.n2582 VSS.n2355 4.5005
R31662 VSS.n2585 VSS.n2355 4.5005
R31663 VSS.n2587 VSS.n2355 4.5005
R31664 VSS.n2588 VSS.n2355 4.5005
R31665 VSS.n2590 VSS.n2355 4.5005
R31666 VSS.n2593 VSS.n2355 4.5005
R31667 VSS.n2595 VSS.n2355 4.5005
R31668 VSS.n2596 VSS.n2355 4.5005
R31669 VSS.n2598 VSS.n2355 4.5005
R31670 VSS.n2601 VSS.n2355 4.5005
R31671 VSS.n2603 VSS.n2355 4.5005
R31672 VSS.n2604 VSS.n2355 4.5005
R31673 VSS.n2606 VSS.n2355 4.5005
R31674 VSS.n2609 VSS.n2355 4.5005
R31675 VSS.n2611 VSS.n2355 4.5005
R31676 VSS.n2612 VSS.n2355 4.5005
R31677 VSS.n2614 VSS.n2355 4.5005
R31678 VSS.n2617 VSS.n2355 4.5005
R31679 VSS.n2619 VSS.n2355 4.5005
R31680 VSS.n2620 VSS.n2355 4.5005
R31681 VSS.n2622 VSS.n2355 4.5005
R31682 VSS.n2625 VSS.n2355 4.5005
R31683 VSS.n2627 VSS.n2355 4.5005
R31684 VSS.n2628 VSS.n2355 4.5005
R31685 VSS.n2630 VSS.n2355 4.5005
R31686 VSS.n2633 VSS.n2355 4.5005
R31687 VSS.n2635 VSS.n2355 4.5005
R31688 VSS.n2636 VSS.n2355 4.5005
R31689 VSS.n2638 VSS.n2355 4.5005
R31690 VSS.n2640 VSS.n2355 4.5005
R31691 VSS.n2642 VSS.n2355 4.5005
R31692 VSS.n2643 VSS.n2355 4.5005
R31693 VSS.n2645 VSS.n2355 4.5005
R31694 VSS.n2648 VSS.n2355 4.5005
R31695 VSS.n2650 VSS.n2355 4.5005
R31696 VSS.n2651 VSS.n2355 4.5005
R31697 VSS.n2653 VSS.n2355 4.5005
R31698 VSS.n2656 VSS.n2355 4.5005
R31699 VSS.n2658 VSS.n2355 4.5005
R31700 VSS.n2659 VSS.n2355 4.5005
R31701 VSS.n2661 VSS.n2355 4.5005
R31702 VSS.n2664 VSS.n2355 4.5005
R31703 VSS.n2666 VSS.n2355 4.5005
R31704 VSS.n2667 VSS.n2355 4.5005
R31705 VSS.n2669 VSS.n2355 4.5005
R31706 VSS.n2672 VSS.n2355 4.5005
R31707 VSS.n2674 VSS.n2355 4.5005
R31708 VSS.n2675 VSS.n2355 4.5005
R31709 VSS.n2677 VSS.n2355 4.5005
R31710 VSS.n2680 VSS.n2355 4.5005
R31711 VSS.n2682 VSS.n2355 4.5005
R31712 VSS.n2683 VSS.n2355 4.5005
R31713 VSS.n2685 VSS.n2355 4.5005
R31714 VSS.n2688 VSS.n2355 4.5005
R31715 VSS.n2690 VSS.n2355 4.5005
R31716 VSS.n2691 VSS.n2355 4.5005
R31717 VSS.n2693 VSS.n2355 4.5005
R31718 VSS.n2696 VSS.n2355 4.5005
R31719 VSS.n2698 VSS.n2355 4.5005
R31720 VSS.n2699 VSS.n2355 4.5005
R31721 VSS.n2701 VSS.n2355 4.5005
R31722 VSS.n2704 VSS.n2355 4.5005
R31723 VSS.n2706 VSS.n2355 4.5005
R31724 VSS.n2707 VSS.n2355 4.5005
R31725 VSS.n2709 VSS.n2355 4.5005
R31726 VSS.n2712 VSS.n2355 4.5005
R31727 VSS.n2714 VSS.n2355 4.5005
R31728 VSS.n2715 VSS.n2355 4.5005
R31729 VSS.n2717 VSS.n2355 4.5005
R31730 VSS.n2720 VSS.n2355 4.5005
R31731 VSS.n2722 VSS.n2355 4.5005
R31732 VSS.n2723 VSS.n2355 4.5005
R31733 VSS.n2725 VSS.n2355 4.5005
R31734 VSS.n2793 VSS.n2355 4.5005
R31735 VSS.n2859 VSS.n2355 4.5005
R31736 VSS.n3051 VSS.n2477 4.5005
R31737 VSS.n2477 VSS.n2351 4.5005
R31738 VSS.n2483 VSS.n2477 4.5005
R31739 VSS.n2484 VSS.n2477 4.5005
R31740 VSS.n2486 VSS.n2477 4.5005
R31741 VSS.n2489 VSS.n2477 4.5005
R31742 VSS.n2491 VSS.n2477 4.5005
R31743 VSS.n2492 VSS.n2477 4.5005
R31744 VSS.n2494 VSS.n2477 4.5005
R31745 VSS.n2497 VSS.n2477 4.5005
R31746 VSS.n2499 VSS.n2477 4.5005
R31747 VSS.n2500 VSS.n2477 4.5005
R31748 VSS.n2502 VSS.n2477 4.5005
R31749 VSS.n2505 VSS.n2477 4.5005
R31750 VSS.n2507 VSS.n2477 4.5005
R31751 VSS.n2508 VSS.n2477 4.5005
R31752 VSS.n2510 VSS.n2477 4.5005
R31753 VSS.n2513 VSS.n2477 4.5005
R31754 VSS.n2515 VSS.n2477 4.5005
R31755 VSS.n2516 VSS.n2477 4.5005
R31756 VSS.n2518 VSS.n2477 4.5005
R31757 VSS.n2521 VSS.n2477 4.5005
R31758 VSS.n2523 VSS.n2477 4.5005
R31759 VSS.n2524 VSS.n2477 4.5005
R31760 VSS.n2526 VSS.n2477 4.5005
R31761 VSS.n2529 VSS.n2477 4.5005
R31762 VSS.n2531 VSS.n2477 4.5005
R31763 VSS.n2532 VSS.n2477 4.5005
R31764 VSS.n2534 VSS.n2477 4.5005
R31765 VSS.n2537 VSS.n2477 4.5005
R31766 VSS.n2539 VSS.n2477 4.5005
R31767 VSS.n2540 VSS.n2477 4.5005
R31768 VSS.n2542 VSS.n2477 4.5005
R31769 VSS.n2545 VSS.n2477 4.5005
R31770 VSS.n2547 VSS.n2477 4.5005
R31771 VSS.n2548 VSS.n2477 4.5005
R31772 VSS.n2550 VSS.n2477 4.5005
R31773 VSS.n2553 VSS.n2477 4.5005
R31774 VSS.n2555 VSS.n2477 4.5005
R31775 VSS.n2556 VSS.n2477 4.5005
R31776 VSS.n2558 VSS.n2477 4.5005
R31777 VSS.n2561 VSS.n2477 4.5005
R31778 VSS.n2563 VSS.n2477 4.5005
R31779 VSS.n2564 VSS.n2477 4.5005
R31780 VSS.n2566 VSS.n2477 4.5005
R31781 VSS.n2569 VSS.n2477 4.5005
R31782 VSS.n2571 VSS.n2477 4.5005
R31783 VSS.n2572 VSS.n2477 4.5005
R31784 VSS.n2574 VSS.n2477 4.5005
R31785 VSS.n2577 VSS.n2477 4.5005
R31786 VSS.n2579 VSS.n2477 4.5005
R31787 VSS.n2580 VSS.n2477 4.5005
R31788 VSS.n2582 VSS.n2477 4.5005
R31789 VSS.n2585 VSS.n2477 4.5005
R31790 VSS.n2587 VSS.n2477 4.5005
R31791 VSS.n2588 VSS.n2477 4.5005
R31792 VSS.n2590 VSS.n2477 4.5005
R31793 VSS.n2593 VSS.n2477 4.5005
R31794 VSS.n2595 VSS.n2477 4.5005
R31795 VSS.n2596 VSS.n2477 4.5005
R31796 VSS.n2598 VSS.n2477 4.5005
R31797 VSS.n2601 VSS.n2477 4.5005
R31798 VSS.n2603 VSS.n2477 4.5005
R31799 VSS.n2604 VSS.n2477 4.5005
R31800 VSS.n2606 VSS.n2477 4.5005
R31801 VSS.n2609 VSS.n2477 4.5005
R31802 VSS.n2611 VSS.n2477 4.5005
R31803 VSS.n2612 VSS.n2477 4.5005
R31804 VSS.n2614 VSS.n2477 4.5005
R31805 VSS.n2617 VSS.n2477 4.5005
R31806 VSS.n2619 VSS.n2477 4.5005
R31807 VSS.n2620 VSS.n2477 4.5005
R31808 VSS.n2622 VSS.n2477 4.5005
R31809 VSS.n2625 VSS.n2477 4.5005
R31810 VSS.n2627 VSS.n2477 4.5005
R31811 VSS.n2628 VSS.n2477 4.5005
R31812 VSS.n2630 VSS.n2477 4.5005
R31813 VSS.n2633 VSS.n2477 4.5005
R31814 VSS.n2635 VSS.n2477 4.5005
R31815 VSS.n2636 VSS.n2477 4.5005
R31816 VSS.n2638 VSS.n2477 4.5005
R31817 VSS.n2640 VSS.n2477 4.5005
R31818 VSS.n2642 VSS.n2477 4.5005
R31819 VSS.n2643 VSS.n2477 4.5005
R31820 VSS.n2645 VSS.n2477 4.5005
R31821 VSS.n2648 VSS.n2477 4.5005
R31822 VSS.n2650 VSS.n2477 4.5005
R31823 VSS.n2651 VSS.n2477 4.5005
R31824 VSS.n2653 VSS.n2477 4.5005
R31825 VSS.n2656 VSS.n2477 4.5005
R31826 VSS.n2658 VSS.n2477 4.5005
R31827 VSS.n2659 VSS.n2477 4.5005
R31828 VSS.n2661 VSS.n2477 4.5005
R31829 VSS.n2664 VSS.n2477 4.5005
R31830 VSS.n2666 VSS.n2477 4.5005
R31831 VSS.n2667 VSS.n2477 4.5005
R31832 VSS.n2669 VSS.n2477 4.5005
R31833 VSS.n2672 VSS.n2477 4.5005
R31834 VSS.n2674 VSS.n2477 4.5005
R31835 VSS.n2675 VSS.n2477 4.5005
R31836 VSS.n2677 VSS.n2477 4.5005
R31837 VSS.n2680 VSS.n2477 4.5005
R31838 VSS.n2682 VSS.n2477 4.5005
R31839 VSS.n2683 VSS.n2477 4.5005
R31840 VSS.n2685 VSS.n2477 4.5005
R31841 VSS.n2688 VSS.n2477 4.5005
R31842 VSS.n2690 VSS.n2477 4.5005
R31843 VSS.n2691 VSS.n2477 4.5005
R31844 VSS.n2693 VSS.n2477 4.5005
R31845 VSS.n2696 VSS.n2477 4.5005
R31846 VSS.n2698 VSS.n2477 4.5005
R31847 VSS.n2699 VSS.n2477 4.5005
R31848 VSS.n2701 VSS.n2477 4.5005
R31849 VSS.n2704 VSS.n2477 4.5005
R31850 VSS.n2706 VSS.n2477 4.5005
R31851 VSS.n2707 VSS.n2477 4.5005
R31852 VSS.n2709 VSS.n2477 4.5005
R31853 VSS.n2712 VSS.n2477 4.5005
R31854 VSS.n2714 VSS.n2477 4.5005
R31855 VSS.n2715 VSS.n2477 4.5005
R31856 VSS.n2717 VSS.n2477 4.5005
R31857 VSS.n2720 VSS.n2477 4.5005
R31858 VSS.n2722 VSS.n2477 4.5005
R31859 VSS.n2723 VSS.n2477 4.5005
R31860 VSS.n2725 VSS.n2477 4.5005
R31861 VSS.n2793 VSS.n2477 4.5005
R31862 VSS.n2859 VSS.n2477 4.5005
R31863 VSS.n3051 VSS.n2354 4.5005
R31864 VSS.n2354 VSS.n2351 4.5005
R31865 VSS.n2483 VSS.n2354 4.5005
R31866 VSS.n2484 VSS.n2354 4.5005
R31867 VSS.n2486 VSS.n2354 4.5005
R31868 VSS.n2489 VSS.n2354 4.5005
R31869 VSS.n2491 VSS.n2354 4.5005
R31870 VSS.n2492 VSS.n2354 4.5005
R31871 VSS.n2494 VSS.n2354 4.5005
R31872 VSS.n2497 VSS.n2354 4.5005
R31873 VSS.n2499 VSS.n2354 4.5005
R31874 VSS.n2500 VSS.n2354 4.5005
R31875 VSS.n2502 VSS.n2354 4.5005
R31876 VSS.n2505 VSS.n2354 4.5005
R31877 VSS.n2507 VSS.n2354 4.5005
R31878 VSS.n2508 VSS.n2354 4.5005
R31879 VSS.n2510 VSS.n2354 4.5005
R31880 VSS.n2513 VSS.n2354 4.5005
R31881 VSS.n2515 VSS.n2354 4.5005
R31882 VSS.n2516 VSS.n2354 4.5005
R31883 VSS.n2518 VSS.n2354 4.5005
R31884 VSS.n2521 VSS.n2354 4.5005
R31885 VSS.n2523 VSS.n2354 4.5005
R31886 VSS.n2524 VSS.n2354 4.5005
R31887 VSS.n2526 VSS.n2354 4.5005
R31888 VSS.n2529 VSS.n2354 4.5005
R31889 VSS.n2531 VSS.n2354 4.5005
R31890 VSS.n2532 VSS.n2354 4.5005
R31891 VSS.n2534 VSS.n2354 4.5005
R31892 VSS.n2537 VSS.n2354 4.5005
R31893 VSS.n2539 VSS.n2354 4.5005
R31894 VSS.n2540 VSS.n2354 4.5005
R31895 VSS.n2542 VSS.n2354 4.5005
R31896 VSS.n2545 VSS.n2354 4.5005
R31897 VSS.n2547 VSS.n2354 4.5005
R31898 VSS.n2548 VSS.n2354 4.5005
R31899 VSS.n2550 VSS.n2354 4.5005
R31900 VSS.n2553 VSS.n2354 4.5005
R31901 VSS.n2555 VSS.n2354 4.5005
R31902 VSS.n2556 VSS.n2354 4.5005
R31903 VSS.n2558 VSS.n2354 4.5005
R31904 VSS.n2561 VSS.n2354 4.5005
R31905 VSS.n2563 VSS.n2354 4.5005
R31906 VSS.n2564 VSS.n2354 4.5005
R31907 VSS.n2566 VSS.n2354 4.5005
R31908 VSS.n2569 VSS.n2354 4.5005
R31909 VSS.n2571 VSS.n2354 4.5005
R31910 VSS.n2572 VSS.n2354 4.5005
R31911 VSS.n2574 VSS.n2354 4.5005
R31912 VSS.n2577 VSS.n2354 4.5005
R31913 VSS.n2579 VSS.n2354 4.5005
R31914 VSS.n2580 VSS.n2354 4.5005
R31915 VSS.n2582 VSS.n2354 4.5005
R31916 VSS.n2585 VSS.n2354 4.5005
R31917 VSS.n2587 VSS.n2354 4.5005
R31918 VSS.n2588 VSS.n2354 4.5005
R31919 VSS.n2590 VSS.n2354 4.5005
R31920 VSS.n2593 VSS.n2354 4.5005
R31921 VSS.n2595 VSS.n2354 4.5005
R31922 VSS.n2596 VSS.n2354 4.5005
R31923 VSS.n2598 VSS.n2354 4.5005
R31924 VSS.n2601 VSS.n2354 4.5005
R31925 VSS.n2603 VSS.n2354 4.5005
R31926 VSS.n2604 VSS.n2354 4.5005
R31927 VSS.n2606 VSS.n2354 4.5005
R31928 VSS.n2609 VSS.n2354 4.5005
R31929 VSS.n2611 VSS.n2354 4.5005
R31930 VSS.n2612 VSS.n2354 4.5005
R31931 VSS.n2614 VSS.n2354 4.5005
R31932 VSS.n2617 VSS.n2354 4.5005
R31933 VSS.n2619 VSS.n2354 4.5005
R31934 VSS.n2620 VSS.n2354 4.5005
R31935 VSS.n2622 VSS.n2354 4.5005
R31936 VSS.n2625 VSS.n2354 4.5005
R31937 VSS.n2627 VSS.n2354 4.5005
R31938 VSS.n2628 VSS.n2354 4.5005
R31939 VSS.n2630 VSS.n2354 4.5005
R31940 VSS.n2633 VSS.n2354 4.5005
R31941 VSS.n2635 VSS.n2354 4.5005
R31942 VSS.n2636 VSS.n2354 4.5005
R31943 VSS.n2638 VSS.n2354 4.5005
R31944 VSS.n2640 VSS.n2354 4.5005
R31945 VSS.n2642 VSS.n2354 4.5005
R31946 VSS.n2643 VSS.n2354 4.5005
R31947 VSS.n2645 VSS.n2354 4.5005
R31948 VSS.n2648 VSS.n2354 4.5005
R31949 VSS.n2650 VSS.n2354 4.5005
R31950 VSS.n2651 VSS.n2354 4.5005
R31951 VSS.n2653 VSS.n2354 4.5005
R31952 VSS.n2656 VSS.n2354 4.5005
R31953 VSS.n2658 VSS.n2354 4.5005
R31954 VSS.n2659 VSS.n2354 4.5005
R31955 VSS.n2661 VSS.n2354 4.5005
R31956 VSS.n2664 VSS.n2354 4.5005
R31957 VSS.n2666 VSS.n2354 4.5005
R31958 VSS.n2667 VSS.n2354 4.5005
R31959 VSS.n2669 VSS.n2354 4.5005
R31960 VSS.n2672 VSS.n2354 4.5005
R31961 VSS.n2674 VSS.n2354 4.5005
R31962 VSS.n2675 VSS.n2354 4.5005
R31963 VSS.n2677 VSS.n2354 4.5005
R31964 VSS.n2680 VSS.n2354 4.5005
R31965 VSS.n2682 VSS.n2354 4.5005
R31966 VSS.n2683 VSS.n2354 4.5005
R31967 VSS.n2685 VSS.n2354 4.5005
R31968 VSS.n2688 VSS.n2354 4.5005
R31969 VSS.n2690 VSS.n2354 4.5005
R31970 VSS.n2691 VSS.n2354 4.5005
R31971 VSS.n2693 VSS.n2354 4.5005
R31972 VSS.n2696 VSS.n2354 4.5005
R31973 VSS.n2698 VSS.n2354 4.5005
R31974 VSS.n2699 VSS.n2354 4.5005
R31975 VSS.n2701 VSS.n2354 4.5005
R31976 VSS.n2704 VSS.n2354 4.5005
R31977 VSS.n2706 VSS.n2354 4.5005
R31978 VSS.n2707 VSS.n2354 4.5005
R31979 VSS.n2709 VSS.n2354 4.5005
R31980 VSS.n2712 VSS.n2354 4.5005
R31981 VSS.n2714 VSS.n2354 4.5005
R31982 VSS.n2715 VSS.n2354 4.5005
R31983 VSS.n2717 VSS.n2354 4.5005
R31984 VSS.n2720 VSS.n2354 4.5005
R31985 VSS.n2722 VSS.n2354 4.5005
R31986 VSS.n2723 VSS.n2354 4.5005
R31987 VSS.n2725 VSS.n2354 4.5005
R31988 VSS.n2793 VSS.n2354 4.5005
R31989 VSS.n2859 VSS.n2354 4.5005
R31990 VSS.n3051 VSS.n2478 4.5005
R31991 VSS.n2478 VSS.n2351 4.5005
R31992 VSS.n2483 VSS.n2478 4.5005
R31993 VSS.n2484 VSS.n2478 4.5005
R31994 VSS.n2486 VSS.n2478 4.5005
R31995 VSS.n2489 VSS.n2478 4.5005
R31996 VSS.n2491 VSS.n2478 4.5005
R31997 VSS.n2492 VSS.n2478 4.5005
R31998 VSS.n2494 VSS.n2478 4.5005
R31999 VSS.n2497 VSS.n2478 4.5005
R32000 VSS.n2499 VSS.n2478 4.5005
R32001 VSS.n2500 VSS.n2478 4.5005
R32002 VSS.n2502 VSS.n2478 4.5005
R32003 VSS.n2505 VSS.n2478 4.5005
R32004 VSS.n2507 VSS.n2478 4.5005
R32005 VSS.n2508 VSS.n2478 4.5005
R32006 VSS.n2510 VSS.n2478 4.5005
R32007 VSS.n2513 VSS.n2478 4.5005
R32008 VSS.n2515 VSS.n2478 4.5005
R32009 VSS.n2516 VSS.n2478 4.5005
R32010 VSS.n2518 VSS.n2478 4.5005
R32011 VSS.n2521 VSS.n2478 4.5005
R32012 VSS.n2523 VSS.n2478 4.5005
R32013 VSS.n2524 VSS.n2478 4.5005
R32014 VSS.n2526 VSS.n2478 4.5005
R32015 VSS.n2529 VSS.n2478 4.5005
R32016 VSS.n2531 VSS.n2478 4.5005
R32017 VSS.n2532 VSS.n2478 4.5005
R32018 VSS.n2534 VSS.n2478 4.5005
R32019 VSS.n2537 VSS.n2478 4.5005
R32020 VSS.n2539 VSS.n2478 4.5005
R32021 VSS.n2540 VSS.n2478 4.5005
R32022 VSS.n2542 VSS.n2478 4.5005
R32023 VSS.n2545 VSS.n2478 4.5005
R32024 VSS.n2547 VSS.n2478 4.5005
R32025 VSS.n2548 VSS.n2478 4.5005
R32026 VSS.n2550 VSS.n2478 4.5005
R32027 VSS.n2553 VSS.n2478 4.5005
R32028 VSS.n2555 VSS.n2478 4.5005
R32029 VSS.n2556 VSS.n2478 4.5005
R32030 VSS.n2558 VSS.n2478 4.5005
R32031 VSS.n2561 VSS.n2478 4.5005
R32032 VSS.n2563 VSS.n2478 4.5005
R32033 VSS.n2564 VSS.n2478 4.5005
R32034 VSS.n2566 VSS.n2478 4.5005
R32035 VSS.n2569 VSS.n2478 4.5005
R32036 VSS.n2571 VSS.n2478 4.5005
R32037 VSS.n2572 VSS.n2478 4.5005
R32038 VSS.n2574 VSS.n2478 4.5005
R32039 VSS.n2577 VSS.n2478 4.5005
R32040 VSS.n2579 VSS.n2478 4.5005
R32041 VSS.n2580 VSS.n2478 4.5005
R32042 VSS.n2582 VSS.n2478 4.5005
R32043 VSS.n2585 VSS.n2478 4.5005
R32044 VSS.n2587 VSS.n2478 4.5005
R32045 VSS.n2588 VSS.n2478 4.5005
R32046 VSS.n2590 VSS.n2478 4.5005
R32047 VSS.n2593 VSS.n2478 4.5005
R32048 VSS.n2595 VSS.n2478 4.5005
R32049 VSS.n2596 VSS.n2478 4.5005
R32050 VSS.n2598 VSS.n2478 4.5005
R32051 VSS.n2601 VSS.n2478 4.5005
R32052 VSS.n2603 VSS.n2478 4.5005
R32053 VSS.n2604 VSS.n2478 4.5005
R32054 VSS.n2606 VSS.n2478 4.5005
R32055 VSS.n2609 VSS.n2478 4.5005
R32056 VSS.n2611 VSS.n2478 4.5005
R32057 VSS.n2612 VSS.n2478 4.5005
R32058 VSS.n2614 VSS.n2478 4.5005
R32059 VSS.n2617 VSS.n2478 4.5005
R32060 VSS.n2619 VSS.n2478 4.5005
R32061 VSS.n2620 VSS.n2478 4.5005
R32062 VSS.n2622 VSS.n2478 4.5005
R32063 VSS.n2625 VSS.n2478 4.5005
R32064 VSS.n2627 VSS.n2478 4.5005
R32065 VSS.n2628 VSS.n2478 4.5005
R32066 VSS.n2630 VSS.n2478 4.5005
R32067 VSS.n2633 VSS.n2478 4.5005
R32068 VSS.n2635 VSS.n2478 4.5005
R32069 VSS.n2636 VSS.n2478 4.5005
R32070 VSS.n2638 VSS.n2478 4.5005
R32071 VSS.n2640 VSS.n2478 4.5005
R32072 VSS.n2642 VSS.n2478 4.5005
R32073 VSS.n2643 VSS.n2478 4.5005
R32074 VSS.n2645 VSS.n2478 4.5005
R32075 VSS.n2648 VSS.n2478 4.5005
R32076 VSS.n2650 VSS.n2478 4.5005
R32077 VSS.n2651 VSS.n2478 4.5005
R32078 VSS.n2653 VSS.n2478 4.5005
R32079 VSS.n2656 VSS.n2478 4.5005
R32080 VSS.n2658 VSS.n2478 4.5005
R32081 VSS.n2659 VSS.n2478 4.5005
R32082 VSS.n2661 VSS.n2478 4.5005
R32083 VSS.n2664 VSS.n2478 4.5005
R32084 VSS.n2666 VSS.n2478 4.5005
R32085 VSS.n2667 VSS.n2478 4.5005
R32086 VSS.n2669 VSS.n2478 4.5005
R32087 VSS.n2672 VSS.n2478 4.5005
R32088 VSS.n2674 VSS.n2478 4.5005
R32089 VSS.n2675 VSS.n2478 4.5005
R32090 VSS.n2677 VSS.n2478 4.5005
R32091 VSS.n2680 VSS.n2478 4.5005
R32092 VSS.n2682 VSS.n2478 4.5005
R32093 VSS.n2683 VSS.n2478 4.5005
R32094 VSS.n2685 VSS.n2478 4.5005
R32095 VSS.n2688 VSS.n2478 4.5005
R32096 VSS.n2690 VSS.n2478 4.5005
R32097 VSS.n2691 VSS.n2478 4.5005
R32098 VSS.n2693 VSS.n2478 4.5005
R32099 VSS.n2696 VSS.n2478 4.5005
R32100 VSS.n2698 VSS.n2478 4.5005
R32101 VSS.n2699 VSS.n2478 4.5005
R32102 VSS.n2701 VSS.n2478 4.5005
R32103 VSS.n2704 VSS.n2478 4.5005
R32104 VSS.n2706 VSS.n2478 4.5005
R32105 VSS.n2707 VSS.n2478 4.5005
R32106 VSS.n2709 VSS.n2478 4.5005
R32107 VSS.n2712 VSS.n2478 4.5005
R32108 VSS.n2714 VSS.n2478 4.5005
R32109 VSS.n2715 VSS.n2478 4.5005
R32110 VSS.n2717 VSS.n2478 4.5005
R32111 VSS.n2720 VSS.n2478 4.5005
R32112 VSS.n2722 VSS.n2478 4.5005
R32113 VSS.n2723 VSS.n2478 4.5005
R32114 VSS.n2725 VSS.n2478 4.5005
R32115 VSS.n2793 VSS.n2478 4.5005
R32116 VSS.n2859 VSS.n2478 4.5005
R32117 VSS.n3051 VSS.n2353 4.5005
R32118 VSS.n2353 VSS.n2351 4.5005
R32119 VSS.n2483 VSS.n2353 4.5005
R32120 VSS.n2484 VSS.n2353 4.5005
R32121 VSS.n2486 VSS.n2353 4.5005
R32122 VSS.n2489 VSS.n2353 4.5005
R32123 VSS.n2491 VSS.n2353 4.5005
R32124 VSS.n2492 VSS.n2353 4.5005
R32125 VSS.n2494 VSS.n2353 4.5005
R32126 VSS.n2497 VSS.n2353 4.5005
R32127 VSS.n2499 VSS.n2353 4.5005
R32128 VSS.n2500 VSS.n2353 4.5005
R32129 VSS.n2502 VSS.n2353 4.5005
R32130 VSS.n2505 VSS.n2353 4.5005
R32131 VSS.n2507 VSS.n2353 4.5005
R32132 VSS.n2508 VSS.n2353 4.5005
R32133 VSS.n2510 VSS.n2353 4.5005
R32134 VSS.n2513 VSS.n2353 4.5005
R32135 VSS.n2515 VSS.n2353 4.5005
R32136 VSS.n2516 VSS.n2353 4.5005
R32137 VSS.n2518 VSS.n2353 4.5005
R32138 VSS.n2521 VSS.n2353 4.5005
R32139 VSS.n2523 VSS.n2353 4.5005
R32140 VSS.n2524 VSS.n2353 4.5005
R32141 VSS.n2526 VSS.n2353 4.5005
R32142 VSS.n2529 VSS.n2353 4.5005
R32143 VSS.n2531 VSS.n2353 4.5005
R32144 VSS.n2532 VSS.n2353 4.5005
R32145 VSS.n2534 VSS.n2353 4.5005
R32146 VSS.n2537 VSS.n2353 4.5005
R32147 VSS.n2539 VSS.n2353 4.5005
R32148 VSS.n2540 VSS.n2353 4.5005
R32149 VSS.n2542 VSS.n2353 4.5005
R32150 VSS.n2545 VSS.n2353 4.5005
R32151 VSS.n2547 VSS.n2353 4.5005
R32152 VSS.n2548 VSS.n2353 4.5005
R32153 VSS.n2550 VSS.n2353 4.5005
R32154 VSS.n2553 VSS.n2353 4.5005
R32155 VSS.n2555 VSS.n2353 4.5005
R32156 VSS.n2556 VSS.n2353 4.5005
R32157 VSS.n2558 VSS.n2353 4.5005
R32158 VSS.n2561 VSS.n2353 4.5005
R32159 VSS.n2563 VSS.n2353 4.5005
R32160 VSS.n2564 VSS.n2353 4.5005
R32161 VSS.n2566 VSS.n2353 4.5005
R32162 VSS.n2569 VSS.n2353 4.5005
R32163 VSS.n2571 VSS.n2353 4.5005
R32164 VSS.n2572 VSS.n2353 4.5005
R32165 VSS.n2574 VSS.n2353 4.5005
R32166 VSS.n2577 VSS.n2353 4.5005
R32167 VSS.n2579 VSS.n2353 4.5005
R32168 VSS.n2580 VSS.n2353 4.5005
R32169 VSS.n2582 VSS.n2353 4.5005
R32170 VSS.n2585 VSS.n2353 4.5005
R32171 VSS.n2587 VSS.n2353 4.5005
R32172 VSS.n2588 VSS.n2353 4.5005
R32173 VSS.n2590 VSS.n2353 4.5005
R32174 VSS.n2593 VSS.n2353 4.5005
R32175 VSS.n2595 VSS.n2353 4.5005
R32176 VSS.n2596 VSS.n2353 4.5005
R32177 VSS.n2598 VSS.n2353 4.5005
R32178 VSS.n2601 VSS.n2353 4.5005
R32179 VSS.n2603 VSS.n2353 4.5005
R32180 VSS.n2604 VSS.n2353 4.5005
R32181 VSS.n2606 VSS.n2353 4.5005
R32182 VSS.n2609 VSS.n2353 4.5005
R32183 VSS.n2611 VSS.n2353 4.5005
R32184 VSS.n2612 VSS.n2353 4.5005
R32185 VSS.n2614 VSS.n2353 4.5005
R32186 VSS.n2617 VSS.n2353 4.5005
R32187 VSS.n2619 VSS.n2353 4.5005
R32188 VSS.n2620 VSS.n2353 4.5005
R32189 VSS.n2622 VSS.n2353 4.5005
R32190 VSS.n2625 VSS.n2353 4.5005
R32191 VSS.n2627 VSS.n2353 4.5005
R32192 VSS.n2628 VSS.n2353 4.5005
R32193 VSS.n2630 VSS.n2353 4.5005
R32194 VSS.n2633 VSS.n2353 4.5005
R32195 VSS.n2635 VSS.n2353 4.5005
R32196 VSS.n2636 VSS.n2353 4.5005
R32197 VSS.n2638 VSS.n2353 4.5005
R32198 VSS.n2640 VSS.n2353 4.5005
R32199 VSS.n2642 VSS.n2353 4.5005
R32200 VSS.n2643 VSS.n2353 4.5005
R32201 VSS.n2645 VSS.n2353 4.5005
R32202 VSS.n2648 VSS.n2353 4.5005
R32203 VSS.n2650 VSS.n2353 4.5005
R32204 VSS.n2651 VSS.n2353 4.5005
R32205 VSS.n2653 VSS.n2353 4.5005
R32206 VSS.n2656 VSS.n2353 4.5005
R32207 VSS.n2658 VSS.n2353 4.5005
R32208 VSS.n2659 VSS.n2353 4.5005
R32209 VSS.n2661 VSS.n2353 4.5005
R32210 VSS.n2664 VSS.n2353 4.5005
R32211 VSS.n2666 VSS.n2353 4.5005
R32212 VSS.n2667 VSS.n2353 4.5005
R32213 VSS.n2669 VSS.n2353 4.5005
R32214 VSS.n2672 VSS.n2353 4.5005
R32215 VSS.n2674 VSS.n2353 4.5005
R32216 VSS.n2675 VSS.n2353 4.5005
R32217 VSS.n2677 VSS.n2353 4.5005
R32218 VSS.n2680 VSS.n2353 4.5005
R32219 VSS.n2682 VSS.n2353 4.5005
R32220 VSS.n2683 VSS.n2353 4.5005
R32221 VSS.n2685 VSS.n2353 4.5005
R32222 VSS.n2688 VSS.n2353 4.5005
R32223 VSS.n2690 VSS.n2353 4.5005
R32224 VSS.n2691 VSS.n2353 4.5005
R32225 VSS.n2693 VSS.n2353 4.5005
R32226 VSS.n2696 VSS.n2353 4.5005
R32227 VSS.n2698 VSS.n2353 4.5005
R32228 VSS.n2699 VSS.n2353 4.5005
R32229 VSS.n2701 VSS.n2353 4.5005
R32230 VSS.n2704 VSS.n2353 4.5005
R32231 VSS.n2706 VSS.n2353 4.5005
R32232 VSS.n2707 VSS.n2353 4.5005
R32233 VSS.n2709 VSS.n2353 4.5005
R32234 VSS.n2712 VSS.n2353 4.5005
R32235 VSS.n2714 VSS.n2353 4.5005
R32236 VSS.n2715 VSS.n2353 4.5005
R32237 VSS.n2717 VSS.n2353 4.5005
R32238 VSS.n2720 VSS.n2353 4.5005
R32239 VSS.n2722 VSS.n2353 4.5005
R32240 VSS.n2723 VSS.n2353 4.5005
R32241 VSS.n2725 VSS.n2353 4.5005
R32242 VSS.n2793 VSS.n2353 4.5005
R32243 VSS.n2859 VSS.n2353 4.5005
R32244 VSS.n3051 VSS.n2479 4.5005
R32245 VSS.n2479 VSS.n2351 4.5005
R32246 VSS.n2483 VSS.n2479 4.5005
R32247 VSS.n2484 VSS.n2479 4.5005
R32248 VSS.n2486 VSS.n2479 4.5005
R32249 VSS.n2489 VSS.n2479 4.5005
R32250 VSS.n2491 VSS.n2479 4.5005
R32251 VSS.n2492 VSS.n2479 4.5005
R32252 VSS.n2494 VSS.n2479 4.5005
R32253 VSS.n2497 VSS.n2479 4.5005
R32254 VSS.n2499 VSS.n2479 4.5005
R32255 VSS.n2500 VSS.n2479 4.5005
R32256 VSS.n2502 VSS.n2479 4.5005
R32257 VSS.n2505 VSS.n2479 4.5005
R32258 VSS.n2507 VSS.n2479 4.5005
R32259 VSS.n2508 VSS.n2479 4.5005
R32260 VSS.n2510 VSS.n2479 4.5005
R32261 VSS.n2513 VSS.n2479 4.5005
R32262 VSS.n2515 VSS.n2479 4.5005
R32263 VSS.n2516 VSS.n2479 4.5005
R32264 VSS.n2518 VSS.n2479 4.5005
R32265 VSS.n2521 VSS.n2479 4.5005
R32266 VSS.n2523 VSS.n2479 4.5005
R32267 VSS.n2524 VSS.n2479 4.5005
R32268 VSS.n2526 VSS.n2479 4.5005
R32269 VSS.n2529 VSS.n2479 4.5005
R32270 VSS.n2531 VSS.n2479 4.5005
R32271 VSS.n2532 VSS.n2479 4.5005
R32272 VSS.n2534 VSS.n2479 4.5005
R32273 VSS.n2537 VSS.n2479 4.5005
R32274 VSS.n2539 VSS.n2479 4.5005
R32275 VSS.n2540 VSS.n2479 4.5005
R32276 VSS.n2542 VSS.n2479 4.5005
R32277 VSS.n2545 VSS.n2479 4.5005
R32278 VSS.n2547 VSS.n2479 4.5005
R32279 VSS.n2548 VSS.n2479 4.5005
R32280 VSS.n2550 VSS.n2479 4.5005
R32281 VSS.n2553 VSS.n2479 4.5005
R32282 VSS.n2555 VSS.n2479 4.5005
R32283 VSS.n2556 VSS.n2479 4.5005
R32284 VSS.n2558 VSS.n2479 4.5005
R32285 VSS.n2561 VSS.n2479 4.5005
R32286 VSS.n2563 VSS.n2479 4.5005
R32287 VSS.n2564 VSS.n2479 4.5005
R32288 VSS.n2566 VSS.n2479 4.5005
R32289 VSS.n2569 VSS.n2479 4.5005
R32290 VSS.n2571 VSS.n2479 4.5005
R32291 VSS.n2572 VSS.n2479 4.5005
R32292 VSS.n2574 VSS.n2479 4.5005
R32293 VSS.n2577 VSS.n2479 4.5005
R32294 VSS.n2579 VSS.n2479 4.5005
R32295 VSS.n2580 VSS.n2479 4.5005
R32296 VSS.n2582 VSS.n2479 4.5005
R32297 VSS.n2585 VSS.n2479 4.5005
R32298 VSS.n2587 VSS.n2479 4.5005
R32299 VSS.n2588 VSS.n2479 4.5005
R32300 VSS.n2590 VSS.n2479 4.5005
R32301 VSS.n2593 VSS.n2479 4.5005
R32302 VSS.n2595 VSS.n2479 4.5005
R32303 VSS.n2596 VSS.n2479 4.5005
R32304 VSS.n2598 VSS.n2479 4.5005
R32305 VSS.n2601 VSS.n2479 4.5005
R32306 VSS.n2603 VSS.n2479 4.5005
R32307 VSS.n2604 VSS.n2479 4.5005
R32308 VSS.n2606 VSS.n2479 4.5005
R32309 VSS.n2609 VSS.n2479 4.5005
R32310 VSS.n2611 VSS.n2479 4.5005
R32311 VSS.n2612 VSS.n2479 4.5005
R32312 VSS.n2614 VSS.n2479 4.5005
R32313 VSS.n2617 VSS.n2479 4.5005
R32314 VSS.n2619 VSS.n2479 4.5005
R32315 VSS.n2620 VSS.n2479 4.5005
R32316 VSS.n2622 VSS.n2479 4.5005
R32317 VSS.n2625 VSS.n2479 4.5005
R32318 VSS.n2627 VSS.n2479 4.5005
R32319 VSS.n2628 VSS.n2479 4.5005
R32320 VSS.n2630 VSS.n2479 4.5005
R32321 VSS.n2633 VSS.n2479 4.5005
R32322 VSS.n2635 VSS.n2479 4.5005
R32323 VSS.n2636 VSS.n2479 4.5005
R32324 VSS.n2638 VSS.n2479 4.5005
R32325 VSS.n2640 VSS.n2479 4.5005
R32326 VSS.n2642 VSS.n2479 4.5005
R32327 VSS.n2643 VSS.n2479 4.5005
R32328 VSS.n2645 VSS.n2479 4.5005
R32329 VSS.n2648 VSS.n2479 4.5005
R32330 VSS.n2650 VSS.n2479 4.5005
R32331 VSS.n2651 VSS.n2479 4.5005
R32332 VSS.n2653 VSS.n2479 4.5005
R32333 VSS.n2656 VSS.n2479 4.5005
R32334 VSS.n2658 VSS.n2479 4.5005
R32335 VSS.n2659 VSS.n2479 4.5005
R32336 VSS.n2661 VSS.n2479 4.5005
R32337 VSS.n2664 VSS.n2479 4.5005
R32338 VSS.n2666 VSS.n2479 4.5005
R32339 VSS.n2667 VSS.n2479 4.5005
R32340 VSS.n2669 VSS.n2479 4.5005
R32341 VSS.n2672 VSS.n2479 4.5005
R32342 VSS.n2674 VSS.n2479 4.5005
R32343 VSS.n2675 VSS.n2479 4.5005
R32344 VSS.n2677 VSS.n2479 4.5005
R32345 VSS.n2680 VSS.n2479 4.5005
R32346 VSS.n2682 VSS.n2479 4.5005
R32347 VSS.n2683 VSS.n2479 4.5005
R32348 VSS.n2685 VSS.n2479 4.5005
R32349 VSS.n2688 VSS.n2479 4.5005
R32350 VSS.n2690 VSS.n2479 4.5005
R32351 VSS.n2691 VSS.n2479 4.5005
R32352 VSS.n2693 VSS.n2479 4.5005
R32353 VSS.n2696 VSS.n2479 4.5005
R32354 VSS.n2698 VSS.n2479 4.5005
R32355 VSS.n2699 VSS.n2479 4.5005
R32356 VSS.n2701 VSS.n2479 4.5005
R32357 VSS.n2704 VSS.n2479 4.5005
R32358 VSS.n2706 VSS.n2479 4.5005
R32359 VSS.n2707 VSS.n2479 4.5005
R32360 VSS.n2709 VSS.n2479 4.5005
R32361 VSS.n2712 VSS.n2479 4.5005
R32362 VSS.n2714 VSS.n2479 4.5005
R32363 VSS.n2715 VSS.n2479 4.5005
R32364 VSS.n2717 VSS.n2479 4.5005
R32365 VSS.n2720 VSS.n2479 4.5005
R32366 VSS.n2722 VSS.n2479 4.5005
R32367 VSS.n2723 VSS.n2479 4.5005
R32368 VSS.n2725 VSS.n2479 4.5005
R32369 VSS.n2793 VSS.n2479 4.5005
R32370 VSS.n2859 VSS.n2479 4.5005
R32371 VSS.n3051 VSS.n2352 4.5005
R32372 VSS.n2352 VSS.n2351 4.5005
R32373 VSS.n2483 VSS.n2352 4.5005
R32374 VSS.n2484 VSS.n2352 4.5005
R32375 VSS.n2486 VSS.n2352 4.5005
R32376 VSS.n2489 VSS.n2352 4.5005
R32377 VSS.n2491 VSS.n2352 4.5005
R32378 VSS.n2492 VSS.n2352 4.5005
R32379 VSS.n2494 VSS.n2352 4.5005
R32380 VSS.n2497 VSS.n2352 4.5005
R32381 VSS.n2499 VSS.n2352 4.5005
R32382 VSS.n2500 VSS.n2352 4.5005
R32383 VSS.n2502 VSS.n2352 4.5005
R32384 VSS.n2505 VSS.n2352 4.5005
R32385 VSS.n2507 VSS.n2352 4.5005
R32386 VSS.n2508 VSS.n2352 4.5005
R32387 VSS.n2510 VSS.n2352 4.5005
R32388 VSS.n2513 VSS.n2352 4.5005
R32389 VSS.n2515 VSS.n2352 4.5005
R32390 VSS.n2516 VSS.n2352 4.5005
R32391 VSS.n2518 VSS.n2352 4.5005
R32392 VSS.n2521 VSS.n2352 4.5005
R32393 VSS.n2523 VSS.n2352 4.5005
R32394 VSS.n2524 VSS.n2352 4.5005
R32395 VSS.n2526 VSS.n2352 4.5005
R32396 VSS.n2529 VSS.n2352 4.5005
R32397 VSS.n2531 VSS.n2352 4.5005
R32398 VSS.n2532 VSS.n2352 4.5005
R32399 VSS.n2534 VSS.n2352 4.5005
R32400 VSS.n2537 VSS.n2352 4.5005
R32401 VSS.n2539 VSS.n2352 4.5005
R32402 VSS.n2540 VSS.n2352 4.5005
R32403 VSS.n2542 VSS.n2352 4.5005
R32404 VSS.n2545 VSS.n2352 4.5005
R32405 VSS.n2547 VSS.n2352 4.5005
R32406 VSS.n2548 VSS.n2352 4.5005
R32407 VSS.n2550 VSS.n2352 4.5005
R32408 VSS.n2553 VSS.n2352 4.5005
R32409 VSS.n2555 VSS.n2352 4.5005
R32410 VSS.n2556 VSS.n2352 4.5005
R32411 VSS.n2558 VSS.n2352 4.5005
R32412 VSS.n2561 VSS.n2352 4.5005
R32413 VSS.n2563 VSS.n2352 4.5005
R32414 VSS.n2564 VSS.n2352 4.5005
R32415 VSS.n2566 VSS.n2352 4.5005
R32416 VSS.n2569 VSS.n2352 4.5005
R32417 VSS.n2571 VSS.n2352 4.5005
R32418 VSS.n2572 VSS.n2352 4.5005
R32419 VSS.n2574 VSS.n2352 4.5005
R32420 VSS.n2577 VSS.n2352 4.5005
R32421 VSS.n2579 VSS.n2352 4.5005
R32422 VSS.n2580 VSS.n2352 4.5005
R32423 VSS.n2582 VSS.n2352 4.5005
R32424 VSS.n2585 VSS.n2352 4.5005
R32425 VSS.n2587 VSS.n2352 4.5005
R32426 VSS.n2588 VSS.n2352 4.5005
R32427 VSS.n2590 VSS.n2352 4.5005
R32428 VSS.n2593 VSS.n2352 4.5005
R32429 VSS.n2595 VSS.n2352 4.5005
R32430 VSS.n2596 VSS.n2352 4.5005
R32431 VSS.n2598 VSS.n2352 4.5005
R32432 VSS.n2601 VSS.n2352 4.5005
R32433 VSS.n2603 VSS.n2352 4.5005
R32434 VSS.n2604 VSS.n2352 4.5005
R32435 VSS.n2606 VSS.n2352 4.5005
R32436 VSS.n2609 VSS.n2352 4.5005
R32437 VSS.n2611 VSS.n2352 4.5005
R32438 VSS.n2612 VSS.n2352 4.5005
R32439 VSS.n2614 VSS.n2352 4.5005
R32440 VSS.n2617 VSS.n2352 4.5005
R32441 VSS.n2619 VSS.n2352 4.5005
R32442 VSS.n2620 VSS.n2352 4.5005
R32443 VSS.n2622 VSS.n2352 4.5005
R32444 VSS.n2625 VSS.n2352 4.5005
R32445 VSS.n2627 VSS.n2352 4.5005
R32446 VSS.n2628 VSS.n2352 4.5005
R32447 VSS.n2630 VSS.n2352 4.5005
R32448 VSS.n2633 VSS.n2352 4.5005
R32449 VSS.n2635 VSS.n2352 4.5005
R32450 VSS.n2636 VSS.n2352 4.5005
R32451 VSS.n2638 VSS.n2352 4.5005
R32452 VSS.n2640 VSS.n2352 4.5005
R32453 VSS.n2642 VSS.n2352 4.5005
R32454 VSS.n2643 VSS.n2352 4.5005
R32455 VSS.n2645 VSS.n2352 4.5005
R32456 VSS.n2648 VSS.n2352 4.5005
R32457 VSS.n2650 VSS.n2352 4.5005
R32458 VSS.n2651 VSS.n2352 4.5005
R32459 VSS.n2653 VSS.n2352 4.5005
R32460 VSS.n2656 VSS.n2352 4.5005
R32461 VSS.n2658 VSS.n2352 4.5005
R32462 VSS.n2659 VSS.n2352 4.5005
R32463 VSS.n2661 VSS.n2352 4.5005
R32464 VSS.n2664 VSS.n2352 4.5005
R32465 VSS.n2666 VSS.n2352 4.5005
R32466 VSS.n2667 VSS.n2352 4.5005
R32467 VSS.n2669 VSS.n2352 4.5005
R32468 VSS.n2672 VSS.n2352 4.5005
R32469 VSS.n2674 VSS.n2352 4.5005
R32470 VSS.n2675 VSS.n2352 4.5005
R32471 VSS.n2677 VSS.n2352 4.5005
R32472 VSS.n2680 VSS.n2352 4.5005
R32473 VSS.n2682 VSS.n2352 4.5005
R32474 VSS.n2683 VSS.n2352 4.5005
R32475 VSS.n2685 VSS.n2352 4.5005
R32476 VSS.n2688 VSS.n2352 4.5005
R32477 VSS.n2690 VSS.n2352 4.5005
R32478 VSS.n2691 VSS.n2352 4.5005
R32479 VSS.n2693 VSS.n2352 4.5005
R32480 VSS.n2696 VSS.n2352 4.5005
R32481 VSS.n2698 VSS.n2352 4.5005
R32482 VSS.n2699 VSS.n2352 4.5005
R32483 VSS.n2701 VSS.n2352 4.5005
R32484 VSS.n2704 VSS.n2352 4.5005
R32485 VSS.n2706 VSS.n2352 4.5005
R32486 VSS.n2707 VSS.n2352 4.5005
R32487 VSS.n2709 VSS.n2352 4.5005
R32488 VSS.n2712 VSS.n2352 4.5005
R32489 VSS.n2714 VSS.n2352 4.5005
R32490 VSS.n2715 VSS.n2352 4.5005
R32491 VSS.n2717 VSS.n2352 4.5005
R32492 VSS.n2720 VSS.n2352 4.5005
R32493 VSS.n2722 VSS.n2352 4.5005
R32494 VSS.n2723 VSS.n2352 4.5005
R32495 VSS.n2725 VSS.n2352 4.5005
R32496 VSS.n2791 VSS.n2352 4.5005
R32497 VSS.n2793 VSS.n2352 4.5005
R32498 VSS.n2859 VSS.n2352 4.5005
R32499 VSS.t42 VSS.n3795 4.02533
R32500 VSS.n3794 VSS.n3793 3.52045
R32501 VSS.n2243 VSS.n2242 3.43927
R32502 VSS.n1699 VSS.n1030 3.34639
R32503 VSS.n3402 VSS.n3401 3.34378
R32504 VSS.n4180 VSS.n4160 3.28169
R32505 VSS.t10 VSS.n3560 3.27652
R32506 VSS.n2242 VSS.n2241 3.25134
R32507 VSS.n3214 VSS.n3213 2.96825
R32508 VSS.n3209 VSS.n3206 2.79275
R32509 VSS.n3054 VSS.n3053 2.77277
R32510 VSS.n4148 VSS.n4147 2.6005
R32511 VSS.n4147 VSS.n4146 2.6005
R32512 VSS.n3855 VSS.n3854 2.6005
R32513 VSS.n675 VSS.n606 2.6005
R32514 VSS.n606 VSS.n457 2.6005
R32515 VSS.n706 VSS.n604 2.6005
R32516 VSS.n3421 VSS.n3420 2.6005
R32517 VSS.n3422 VSS.n3421 2.6005
R32518 VSS.n3506 VSS.n3505 2.6005
R32519 VSS.n1753 VSS.n1752 2.6005
R32520 VSS.n2184 VSS.n2183 2.6005
R32521 VSS.n2185 VSS.n2184 2.6005
R32522 VSS.n2100 VSS.n2099 2.6005
R32523 VSS.n1917 VSS.n1656 2.6005
R32524 VSS.n2185 VSS.n1656 2.6005
R32525 VSS.n2005 VSS.n2004 2.6005
R32526 VSS.n2005 VSS.n1620 2.6005
R32527 VSS.n4503 VSS.n4188 2.59835
R32528 VSS.n2099 VSS.n2098 2.45036
R32529 VSS.n3507 VSS.n3506 2.45036
R32530 VSS.n1754 VSS.n1753 2.45036
R32531 VSS.n3854 VSS.n709 2.45036
R32532 VSS.n3802 VSS.n706 2.45036
R32533 VSS.n4179 VSS.n4178 2.438
R32534 VSS.n4503 VSS.n4415 2.25083
R32535 VSS.n4503 VSS.n446 2.25083
R32536 VSS.n4503 VSS.n445 2.25083
R32537 VSS.n4503 VSS.n444 2.25083
R32538 VSS.n4503 VSS.n443 2.25083
R32539 VSS.n4503 VSS.n442 2.25083
R32540 VSS.n4503 VSS.n441 2.25083
R32541 VSS.n4503 VSS.n440 2.25083
R32542 VSS.n4503 VSS.n439 2.25083
R32543 VSS.n4503 VSS.n438 2.25083
R32544 VSS.n4503 VSS.n437 2.25083
R32545 VSS.n4503 VSS.n436 2.25083
R32546 VSS.n4503 VSS.n435 2.25083
R32547 VSS.n4503 VSS.n434 2.25083
R32548 VSS.n4503 VSS.n433 2.25083
R32549 VSS.n4503 VSS.n432 2.25083
R32550 VSS.n4503 VSS.n431 2.25083
R32551 VSS.n4503 VSS.n430 2.25083
R32552 VSS.n4503 VSS.n429 2.25083
R32553 VSS.n4503 VSS.n428 2.25083
R32554 VSS.n4503 VSS.n427 2.25083
R32555 VSS.n4503 VSS.n426 2.25083
R32556 VSS.n4503 VSS.n425 2.25083
R32557 VSS.n4503 VSS.n424 2.25083
R32558 VSS.n4503 VSS.n423 2.25083
R32559 VSS.n4503 VSS.n422 2.25083
R32560 VSS.n4503 VSS.n421 2.25083
R32561 VSS.n4503 VSS.n420 2.25083
R32562 VSS.n4503 VSS.n419 2.25083
R32563 VSS.n4503 VSS.n418 2.25083
R32564 VSS.n4503 VSS.n417 2.25083
R32565 VSS.n4503 VSS.n416 2.25083
R32566 VSS.n4503 VSS.n415 2.25083
R32567 VSS.n4503 VSS.n414 2.25083
R32568 VSS.n4503 VSS.n413 2.25083
R32569 VSS.n4503 VSS.n412 2.25083
R32570 VSS.n4503 VSS.n411 2.25083
R32571 VSS.n4503 VSS.n410 2.25083
R32572 VSS.n4503 VSS.n409 2.25083
R32573 VSS.n4503 VSS.n408 2.25083
R32574 VSS.n4503 VSS.n407 2.25083
R32575 VSS.n4503 VSS.n4 2.25083
R32576 VSS.n4503 VSS.n406 2.25083
R32577 VSS.n4503 VSS.n405 2.25083
R32578 VSS.n4503 VSS.n404 2.25083
R32579 VSS.n4503 VSS.n403 2.25083
R32580 VSS.n4503 VSS.n402 2.25083
R32581 VSS.n4503 VSS.n401 2.25083
R32582 VSS.n4503 VSS.n400 2.25083
R32583 VSS.n4503 VSS.n399 2.25083
R32584 VSS.n4503 VSS.n398 2.25083
R32585 VSS.n4503 VSS.n397 2.25083
R32586 VSS.n4503 VSS.n396 2.25083
R32587 VSS.n4503 VSS.n395 2.25083
R32588 VSS.n4503 VSS.n394 2.25083
R32589 VSS.n4503 VSS.n393 2.25083
R32590 VSS.n4503 VSS.n392 2.25083
R32591 VSS.n4503 VSS.n391 2.25083
R32592 VSS.n4503 VSS.n390 2.25083
R32593 VSS.n4503 VSS.n389 2.25083
R32594 VSS.n4503 VSS.n388 2.25083
R32595 VSS.n4503 VSS.n387 2.25083
R32596 VSS.n4503 VSS.n386 2.25083
R32597 VSS.n385 VSS.n321 2.25083
R32598 VSS.n383 VSS.n382 2.25083
R32599 VSS.n383 VSS.n381 2.25083
R32600 VSS.n383 VSS.n380 2.25083
R32601 VSS.n383 VSS.n379 2.25083
R32602 VSS.n383 VSS.n378 2.25083
R32603 VSS.n383 VSS.n377 2.25083
R32604 VSS.n383 VSS.n376 2.25083
R32605 VSS.n383 VSS.n375 2.25083
R32606 VSS.n383 VSS.n374 2.25083
R32607 VSS.n383 VSS.n373 2.25083
R32608 VSS.n383 VSS.n372 2.25083
R32609 VSS.n383 VSS.n371 2.25083
R32610 VSS.n383 VSS.n370 2.25083
R32611 VSS.n383 VSS.n369 2.25083
R32612 VSS.n383 VSS.n368 2.25083
R32613 VSS.n383 VSS.n367 2.25083
R32614 VSS.n383 VSS.n366 2.25083
R32615 VSS.n383 VSS.n365 2.25083
R32616 VSS.n383 VSS.n364 2.25083
R32617 VSS.n383 VSS.n363 2.25083
R32618 VSS.n383 VSS.n362 2.25083
R32619 VSS.n383 VSS.n361 2.25083
R32620 VSS.n383 VSS.n360 2.25083
R32621 VSS.n383 VSS.n359 2.25083
R32622 VSS.n383 VSS.n358 2.25083
R32623 VSS.n383 VSS.n357 2.25083
R32624 VSS.n383 VSS.n356 2.25083
R32625 VSS.n383 VSS.n355 2.25083
R32626 VSS.n383 VSS.n354 2.25083
R32627 VSS.n383 VSS.n353 2.25083
R32628 VSS.n383 VSS.n352 2.25083
R32629 VSS.n383 VSS.n351 2.25083
R32630 VSS.n383 VSS.n350 2.25083
R32631 VSS.n383 VSS.n349 2.25083
R32632 VSS.n383 VSS.n348 2.25083
R32633 VSS.n383 VSS.n347 2.25083
R32634 VSS.n383 VSS.n346 2.25083
R32635 VSS.n383 VSS.n345 2.25083
R32636 VSS.n383 VSS.n344 2.25083
R32637 VSS.n383 VSS.n343 2.25083
R32638 VSS.n383 VSS.n342 2.25083
R32639 VSS.n383 VSS.n68 2.25083
R32640 VSS.n383 VSS.n341 2.25083
R32641 VSS.n383 VSS.n340 2.25083
R32642 VSS.n383 VSS.n339 2.25083
R32643 VSS.n383 VSS.n338 2.25083
R32644 VSS.n383 VSS.n337 2.25083
R32645 VSS.n383 VSS.n336 2.25083
R32646 VSS.n383 VSS.n335 2.25083
R32647 VSS.n383 VSS.n334 2.25083
R32648 VSS.n383 VSS.n333 2.25083
R32649 VSS.n383 VSS.n332 2.25083
R32650 VSS.n383 VSS.n331 2.25083
R32651 VSS.n383 VSS.n330 2.25083
R32652 VSS.n383 VSS.n329 2.25083
R32653 VSS.n383 VSS.n328 2.25083
R32654 VSS.n383 VSS.n327 2.25083
R32655 VSS.n383 VSS.n326 2.25083
R32656 VSS.n383 VSS.n325 2.25083
R32657 VSS.n383 VSS.n324 2.25083
R32658 VSS.n383 VSS.n323 2.25083
R32659 VSS.n383 VSS.n322 2.25083
R32660 VSS.n4416 VSS.n383 2.25083
R32661 VSS.n4414 VSS.n4251 2.25083
R32662 VSS.n321 VSS.n258 2.25083
R32663 VSS.n4414 VSS.n4250 2.25083
R32664 VSS.n321 VSS.n259 2.25083
R32665 VSS.n4414 VSS.n4249 2.25083
R32666 VSS.n321 VSS.n260 2.25083
R32667 VSS.n4414 VSS.n4248 2.25083
R32668 VSS.n321 VSS.n261 2.25083
R32669 VSS.n4414 VSS.n4247 2.25083
R32670 VSS.n321 VSS.n262 2.25083
R32671 VSS.n4414 VSS.n4246 2.25083
R32672 VSS.n321 VSS.n263 2.25083
R32673 VSS.n4414 VSS.n4245 2.25083
R32674 VSS.n321 VSS.n264 2.25083
R32675 VSS.n4414 VSS.n4244 2.25083
R32676 VSS.n321 VSS.n265 2.25083
R32677 VSS.n4414 VSS.n4243 2.25083
R32678 VSS.n321 VSS.n266 2.25083
R32679 VSS.n4414 VSS.n4242 2.25083
R32680 VSS.n321 VSS.n267 2.25083
R32681 VSS.n4414 VSS.n4241 2.25083
R32682 VSS.n321 VSS.n268 2.25083
R32683 VSS.n4414 VSS.n4240 2.25083
R32684 VSS.n321 VSS.n269 2.25083
R32685 VSS.n4414 VSS.n4239 2.25083
R32686 VSS.n321 VSS.n270 2.25083
R32687 VSS.n4414 VSS.n4238 2.25083
R32688 VSS.n321 VSS.n271 2.25083
R32689 VSS.n4414 VSS.n4237 2.25083
R32690 VSS.n321 VSS.n272 2.25083
R32691 VSS.n4414 VSS.n4236 2.25083
R32692 VSS.n321 VSS.n273 2.25083
R32693 VSS.n4414 VSS.n4235 2.25083
R32694 VSS.n321 VSS.n274 2.25083
R32695 VSS.n4414 VSS.n4234 2.25083
R32696 VSS.n321 VSS.n275 2.25083
R32697 VSS.n4414 VSS.n4233 2.25083
R32698 VSS.n321 VSS.n276 2.25083
R32699 VSS.n4414 VSS.n4232 2.25083
R32700 VSS.n321 VSS.n277 2.25083
R32701 VSS.n4414 VSS.n4231 2.25083
R32702 VSS.n321 VSS.n278 2.25083
R32703 VSS.n4414 VSS.n4230 2.25083
R32704 VSS.n321 VSS.n279 2.25083
R32705 VSS.n4414 VSS.n4229 2.25083
R32706 VSS.n321 VSS.n280 2.25083
R32707 VSS.n4414 VSS.n4228 2.25083
R32708 VSS.n321 VSS.n281 2.25083
R32709 VSS.n4414 VSS.n4227 2.25083
R32710 VSS.n321 VSS.n282 2.25083
R32711 VSS.n4414 VSS.n4226 2.25083
R32712 VSS.n321 VSS.n283 2.25083
R32713 VSS.n4414 VSS.n4225 2.25083
R32714 VSS.n321 VSS.n284 2.25083
R32715 VSS.n4414 VSS.n4224 2.25083
R32716 VSS.n321 VSS.n285 2.25083
R32717 VSS.n4414 VSS.n4223 2.25083
R32718 VSS.n321 VSS.n286 2.25083
R32719 VSS.n4414 VSS.n4222 2.25083
R32720 VSS.n321 VSS.n287 2.25083
R32721 VSS.n4414 VSS.n4221 2.25083
R32722 VSS.n321 VSS.n288 2.25083
R32723 VSS.n4414 VSS.n4220 2.25083
R32724 VSS.n321 VSS.n289 2.25083
R32725 VSS.n4414 VSS.n4219 2.25083
R32726 VSS.n321 VSS.n290 2.25083
R32727 VSS.n4414 VSS.n4218 2.25083
R32728 VSS.n321 VSS.n291 2.25083
R32729 VSS.n4414 VSS.n4217 2.25083
R32730 VSS.n321 VSS.n292 2.25083
R32731 VSS.n4414 VSS.n4216 2.25083
R32732 VSS.n321 VSS.n293 2.25083
R32733 VSS.n4414 VSS.n4215 2.25083
R32734 VSS.n321 VSS.n294 2.25083
R32735 VSS.n4414 VSS.n4214 2.25083
R32736 VSS.n321 VSS.n295 2.25083
R32737 VSS.n4414 VSS.n4213 2.25083
R32738 VSS.n321 VSS.n296 2.25083
R32739 VSS.n4414 VSS.n4212 2.25083
R32740 VSS.n321 VSS.n297 2.25083
R32741 VSS.n4414 VSS.n4211 2.25083
R32742 VSS.n321 VSS.n298 2.25083
R32743 VSS.n4414 VSS.n4210 2.25083
R32744 VSS.n321 VSS.n299 2.25083
R32745 VSS.n4414 VSS.n4209 2.25083
R32746 VSS.n321 VSS.n300 2.25083
R32747 VSS.n4414 VSS.n4208 2.25083
R32748 VSS.n321 VSS.n301 2.25083
R32749 VSS.n4414 VSS.n4207 2.25083
R32750 VSS.n321 VSS.n302 2.25083
R32751 VSS.n4414 VSS.n4206 2.25083
R32752 VSS.n321 VSS.n303 2.25083
R32753 VSS.n4414 VSS.n4205 2.25083
R32754 VSS.n321 VSS.n304 2.25083
R32755 VSS.n4414 VSS.n4204 2.25083
R32756 VSS.n321 VSS.n305 2.25083
R32757 VSS.n4414 VSS.n4203 2.25083
R32758 VSS.n321 VSS.n306 2.25083
R32759 VSS.n4414 VSS.n4202 2.25083
R32760 VSS.n321 VSS.n307 2.25083
R32761 VSS.n4414 VSS.n4201 2.25083
R32762 VSS.n321 VSS.n308 2.25083
R32763 VSS.n4414 VSS.n4200 2.25083
R32764 VSS.n321 VSS.n309 2.25083
R32765 VSS.n4414 VSS.n4199 2.25083
R32766 VSS.n321 VSS.n310 2.25083
R32767 VSS.n4414 VSS.n4198 2.25083
R32768 VSS.n321 VSS.n311 2.25083
R32769 VSS.n4414 VSS.n4197 2.25083
R32770 VSS.n321 VSS.n312 2.25083
R32771 VSS.n4414 VSS.n4196 2.25083
R32772 VSS.n321 VSS.n313 2.25083
R32773 VSS.n4414 VSS.n4195 2.25083
R32774 VSS.n321 VSS.n314 2.25083
R32775 VSS.n4414 VSS.n4194 2.25083
R32776 VSS.n321 VSS.n315 2.25083
R32777 VSS.n4414 VSS.n4193 2.25083
R32778 VSS.n321 VSS.n316 2.25083
R32779 VSS.n4414 VSS.n4192 2.25083
R32780 VSS.n321 VSS.n317 2.25083
R32781 VSS.n4414 VSS.n4191 2.25083
R32782 VSS.n321 VSS.n318 2.25083
R32783 VSS.n4414 VSS.n4190 2.25083
R32784 VSS.n321 VSS.n319 2.25083
R32785 VSS.n4414 VSS.n4189 2.25083
R32786 VSS.n321 VSS.n320 2.25083
R32787 VSS.n4414 VSS.n194 2.25083
R32788 VSS.n4505 VSS.n257 2.25083
R32789 VSS.n3053 VSS.n3052 2.25083
R32790 VSS.n3053 VSS.n2350 2.25083
R32791 VSS.n3053 VSS.n2349 2.25083
R32792 VSS.n3053 VSS.n2348 2.25083
R32793 VSS.n3053 VSS.n2347 2.25083
R32794 VSS.n3053 VSS.n2346 2.25083
R32795 VSS.n3053 VSS.n2345 2.25083
R32796 VSS.n3053 VSS.n2344 2.25083
R32797 VSS.n3053 VSS.n2343 2.25083
R32798 VSS.n3053 VSS.n2342 2.25083
R32799 VSS.n3053 VSS.n2341 2.25083
R32800 VSS.n3053 VSS.n2340 2.25083
R32801 VSS.n3053 VSS.n2339 2.25083
R32802 VSS.n3053 VSS.n2338 2.25083
R32803 VSS.n3053 VSS.n2337 2.25083
R32804 VSS.n3053 VSS.n2336 2.25083
R32805 VSS.n3053 VSS.n2335 2.25083
R32806 VSS.n3053 VSS.n2334 2.25083
R32807 VSS.n3053 VSS.n2333 2.25083
R32808 VSS.n3053 VSS.n2332 2.25083
R32809 VSS.n3053 VSS.n2331 2.25083
R32810 VSS.n3053 VSS.n2330 2.25083
R32811 VSS.n3053 VSS.n2329 2.25083
R32812 VSS.n3053 VSS.n2328 2.25083
R32813 VSS.n3053 VSS.n2327 2.25083
R32814 VSS.n3053 VSS.n2326 2.25083
R32815 VSS.n3053 VSS.n2325 2.25083
R32816 VSS.n3053 VSS.n2324 2.25083
R32817 VSS.n3053 VSS.n2323 2.25083
R32818 VSS.n3053 VSS.n2322 2.25083
R32819 VSS.n3053 VSS.n2321 2.25083
R32820 VSS.n3053 VSS.n2320 2.25083
R32821 VSS.n3053 VSS.n2319 2.25083
R32822 VSS.n3053 VSS.n2318 2.25083
R32823 VSS.n3053 VSS.n2317 2.25083
R32824 VSS.n3053 VSS.n2316 2.25083
R32825 VSS.n3053 VSS.n2315 2.25083
R32826 VSS.n3053 VSS.n2314 2.25083
R32827 VSS.n3053 VSS.n2313 2.25083
R32828 VSS.n3053 VSS.n2312 2.25083
R32829 VSS.n3053 VSS.n2311 2.25083
R32830 VSS.n3053 VSS.n2310 2.25083
R32831 VSS.n3053 VSS.n2309 2.25083
R32832 VSS.n3053 VSS.n2308 2.25083
R32833 VSS.n3053 VSS.n2307 2.25083
R32834 VSS.n3053 VSS.n2306 2.25083
R32835 VSS.n3053 VSS.n2305 2.25083
R32836 VSS.n3053 VSS.n2304 2.25083
R32837 VSS.n3053 VSS.n2303 2.25083
R32838 VSS.n3053 VSS.n2302 2.25083
R32839 VSS.n3053 VSS.n2301 2.25083
R32840 VSS.n3053 VSS.n2300 2.25083
R32841 VSS.n3053 VSS.n2299 2.25083
R32842 VSS.n3053 VSS.n2298 2.25083
R32843 VSS.n3053 VSS.n2297 2.25083
R32844 VSS.n3053 VSS.n2296 2.25083
R32845 VSS.n3053 VSS.n2295 2.25083
R32846 VSS.n3053 VSS.n2294 2.25083
R32847 VSS.n3053 VSS.n2293 2.25083
R32848 VSS.n3053 VSS.n2292 2.25083
R32849 VSS.n3053 VSS.n2291 2.25083
R32850 VSS.n3053 VSS.n2290 2.25083
R32851 VSS.n3053 VSS.n2289 2.25083
R32852 VSS.n3053 VSS.n2288 2.25083
R32853 VSS.n2859 VSS.n2287 2.25083
R32854 VSS.n2482 VSS.n2416 2.25083
R32855 VSS.n2485 VSS.n2416 2.25083
R32856 VSS.n2490 VSS.n2416 2.25083
R32857 VSS.n2493 VSS.n2416 2.25083
R32858 VSS.n2498 VSS.n2416 2.25083
R32859 VSS.n2501 VSS.n2416 2.25083
R32860 VSS.n2506 VSS.n2416 2.25083
R32861 VSS.n2509 VSS.n2416 2.25083
R32862 VSS.n2514 VSS.n2416 2.25083
R32863 VSS.n2517 VSS.n2416 2.25083
R32864 VSS.n2522 VSS.n2416 2.25083
R32865 VSS.n2525 VSS.n2416 2.25083
R32866 VSS.n2530 VSS.n2416 2.25083
R32867 VSS.n2533 VSS.n2416 2.25083
R32868 VSS.n2538 VSS.n2416 2.25083
R32869 VSS.n2541 VSS.n2416 2.25083
R32870 VSS.n2546 VSS.n2416 2.25083
R32871 VSS.n2549 VSS.n2416 2.25083
R32872 VSS.n2554 VSS.n2416 2.25083
R32873 VSS.n2557 VSS.n2416 2.25083
R32874 VSS.n2562 VSS.n2416 2.25083
R32875 VSS.n2565 VSS.n2416 2.25083
R32876 VSS.n2570 VSS.n2416 2.25083
R32877 VSS.n2573 VSS.n2416 2.25083
R32878 VSS.n2578 VSS.n2416 2.25083
R32879 VSS.n2581 VSS.n2416 2.25083
R32880 VSS.n2586 VSS.n2416 2.25083
R32881 VSS.n2589 VSS.n2416 2.25083
R32882 VSS.n2594 VSS.n2416 2.25083
R32883 VSS.n2597 VSS.n2416 2.25083
R32884 VSS.n2602 VSS.n2416 2.25083
R32885 VSS.n2605 VSS.n2416 2.25083
R32886 VSS.n2610 VSS.n2416 2.25083
R32887 VSS.n2613 VSS.n2416 2.25083
R32888 VSS.n2618 VSS.n2416 2.25083
R32889 VSS.n2621 VSS.n2416 2.25083
R32890 VSS.n2626 VSS.n2416 2.25083
R32891 VSS.n2629 VSS.n2416 2.25083
R32892 VSS.n2634 VSS.n2416 2.25083
R32893 VSS.n2637 VSS.n2416 2.25083
R32894 VSS.n2641 VSS.n2416 2.25083
R32895 VSS.n2644 VSS.n2416 2.25083
R32896 VSS.n2649 VSS.n2416 2.25083
R32897 VSS.n2652 VSS.n2416 2.25083
R32898 VSS.n2657 VSS.n2416 2.25083
R32899 VSS.n2660 VSS.n2416 2.25083
R32900 VSS.n2665 VSS.n2416 2.25083
R32901 VSS.n2668 VSS.n2416 2.25083
R32902 VSS.n2673 VSS.n2416 2.25083
R32903 VSS.n2676 VSS.n2416 2.25083
R32904 VSS.n2681 VSS.n2416 2.25083
R32905 VSS.n2684 VSS.n2416 2.25083
R32906 VSS.n2689 VSS.n2416 2.25083
R32907 VSS.n2692 VSS.n2416 2.25083
R32908 VSS.n2697 VSS.n2416 2.25083
R32909 VSS.n2700 VSS.n2416 2.25083
R32910 VSS.n2705 VSS.n2416 2.25083
R32911 VSS.n2708 VSS.n2416 2.25083
R32912 VSS.n2713 VSS.n2416 2.25083
R32913 VSS.n2716 VSS.n2416 2.25083
R32914 VSS.n2721 VSS.n2416 2.25083
R32915 VSS.n2724 VSS.n2416 2.25083
R32916 VSS.n2792 VSS.n2416 2.25083
R32917 VSS.n2858 VSS.n2794 2.25083
R32918 VSS.n2791 VSS.n2790 2.25083
R32919 VSS.n2858 VSS.n2795 2.25083
R32920 VSS.n2791 VSS.n2789 2.25083
R32921 VSS.n2858 VSS.n2796 2.25083
R32922 VSS.n2791 VSS.n2788 2.25083
R32923 VSS.n2858 VSS.n2797 2.25083
R32924 VSS.n2791 VSS.n2787 2.25083
R32925 VSS.n2858 VSS.n2798 2.25083
R32926 VSS.n2791 VSS.n2786 2.25083
R32927 VSS.n2858 VSS.n2799 2.25083
R32928 VSS.n2791 VSS.n2785 2.25083
R32929 VSS.n2858 VSS.n2800 2.25083
R32930 VSS.n2791 VSS.n2784 2.25083
R32931 VSS.n2858 VSS.n2801 2.25083
R32932 VSS.n2791 VSS.n2783 2.25083
R32933 VSS.n2858 VSS.n2802 2.25083
R32934 VSS.n2791 VSS.n2782 2.25083
R32935 VSS.n2858 VSS.n2803 2.25083
R32936 VSS.n2791 VSS.n2781 2.25083
R32937 VSS.n2858 VSS.n2804 2.25083
R32938 VSS.n2791 VSS.n2780 2.25083
R32939 VSS.n2858 VSS.n2805 2.25083
R32940 VSS.n2791 VSS.n2779 2.25083
R32941 VSS.n2858 VSS.n2806 2.25083
R32942 VSS.n2791 VSS.n2778 2.25083
R32943 VSS.n2858 VSS.n2807 2.25083
R32944 VSS.n2791 VSS.n2777 2.25083
R32945 VSS.n2858 VSS.n2808 2.25083
R32946 VSS.n2791 VSS.n2776 2.25083
R32947 VSS.n2858 VSS.n2809 2.25083
R32948 VSS.n2791 VSS.n2775 2.25083
R32949 VSS.n2858 VSS.n2810 2.25083
R32950 VSS.n2791 VSS.n2774 2.25083
R32951 VSS.n2858 VSS.n2811 2.25083
R32952 VSS.n2791 VSS.n2773 2.25083
R32953 VSS.n2858 VSS.n2812 2.25083
R32954 VSS.n2791 VSS.n2772 2.25083
R32955 VSS.n2858 VSS.n2813 2.25083
R32956 VSS.n2791 VSS.n2771 2.25083
R32957 VSS.n2858 VSS.n2814 2.25083
R32958 VSS.n2791 VSS.n2770 2.25083
R32959 VSS.n2858 VSS.n2815 2.25083
R32960 VSS.n2791 VSS.n2769 2.25083
R32961 VSS.n2858 VSS.n2816 2.25083
R32962 VSS.n2791 VSS.n2768 2.25083
R32963 VSS.n2858 VSS.n2817 2.25083
R32964 VSS.n2791 VSS.n2767 2.25083
R32965 VSS.n2858 VSS.n2818 2.25083
R32966 VSS.n2791 VSS.n2766 2.25083
R32967 VSS.n2858 VSS.n2819 2.25083
R32968 VSS.n2791 VSS.n2765 2.25083
R32969 VSS.n2858 VSS.n2820 2.25083
R32970 VSS.n2791 VSS.n2764 2.25083
R32971 VSS.n2858 VSS.n2821 2.25083
R32972 VSS.n2791 VSS.n2763 2.25083
R32973 VSS.n2858 VSS.n2822 2.25083
R32974 VSS.n2791 VSS.n2762 2.25083
R32975 VSS.n2858 VSS.n2823 2.25083
R32976 VSS.n2791 VSS.n2761 2.25083
R32977 VSS.n2858 VSS.n2824 2.25083
R32978 VSS.n2791 VSS.n2760 2.25083
R32979 VSS.n2858 VSS.n2825 2.25083
R32980 VSS.n2791 VSS.n2759 2.25083
R32981 VSS.n2858 VSS.n2826 2.25083
R32982 VSS.n2791 VSS.n2758 2.25083
R32983 VSS.n2858 VSS.n2827 2.25083
R32984 VSS.n2791 VSS.n2757 2.25083
R32985 VSS.n2858 VSS.n2828 2.25083
R32986 VSS.n2791 VSS.n2756 2.25083
R32987 VSS.n2858 VSS.n2829 2.25083
R32988 VSS.n2791 VSS.n2755 2.25083
R32989 VSS.n2858 VSS.n2830 2.25083
R32990 VSS.n2791 VSS.n2754 2.25083
R32991 VSS.n2858 VSS.n2831 2.25083
R32992 VSS.n2791 VSS.n2753 2.25083
R32993 VSS.n2858 VSS.n2832 2.25083
R32994 VSS.n2791 VSS.n2752 2.25083
R32995 VSS.n2858 VSS.n2833 2.25083
R32996 VSS.n2791 VSS.n2751 2.25083
R32997 VSS.n2858 VSS.n2834 2.25083
R32998 VSS.n2791 VSS.n2750 2.25083
R32999 VSS.n2858 VSS.n2835 2.25083
R33000 VSS.n2791 VSS.n2749 2.25083
R33001 VSS.n2858 VSS.n2836 2.25083
R33002 VSS.n2791 VSS.n2748 2.25083
R33003 VSS.n2858 VSS.n2837 2.25083
R33004 VSS.n2791 VSS.n2747 2.25083
R33005 VSS.n2858 VSS.n2838 2.25083
R33006 VSS.n2791 VSS.n2746 2.25083
R33007 VSS.n2858 VSS.n2839 2.25083
R33008 VSS.n2791 VSS.n2745 2.25083
R33009 VSS.n2858 VSS.n2840 2.25083
R33010 VSS.n2791 VSS.n2744 2.25083
R33011 VSS.n2858 VSS.n2841 2.25083
R33012 VSS.n2791 VSS.n2743 2.25083
R33013 VSS.n2858 VSS.n2842 2.25083
R33014 VSS.n2791 VSS.n2742 2.25083
R33015 VSS.n2858 VSS.n2843 2.25083
R33016 VSS.n2791 VSS.n2741 2.25083
R33017 VSS.n2858 VSS.n2844 2.25083
R33018 VSS.n2791 VSS.n2740 2.25083
R33019 VSS.n2858 VSS.n2845 2.25083
R33020 VSS.n2791 VSS.n2739 2.25083
R33021 VSS.n2858 VSS.n2846 2.25083
R33022 VSS.n2791 VSS.n2738 2.25083
R33023 VSS.n2858 VSS.n2847 2.25083
R33024 VSS.n2791 VSS.n2737 2.25083
R33025 VSS.n2858 VSS.n2848 2.25083
R33026 VSS.n2791 VSS.n2736 2.25083
R33027 VSS.n2858 VSS.n2849 2.25083
R33028 VSS.n2791 VSS.n2735 2.25083
R33029 VSS.n2858 VSS.n2850 2.25083
R33030 VSS.n2791 VSS.n2734 2.25083
R33031 VSS.n2858 VSS.n2851 2.25083
R33032 VSS.n2791 VSS.n2733 2.25083
R33033 VSS.n2858 VSS.n2852 2.25083
R33034 VSS.n2791 VSS.n2732 2.25083
R33035 VSS.n2858 VSS.n2853 2.25083
R33036 VSS.n2791 VSS.n2731 2.25083
R33037 VSS.n2858 VSS.n2854 2.25083
R33038 VSS.n2791 VSS.n2730 2.25083
R33039 VSS.n2858 VSS.n2855 2.25083
R33040 VSS.n2791 VSS.n2729 2.25083
R33041 VSS.n2858 VSS.n2856 2.25083
R33042 VSS.n2791 VSS.n2728 2.25083
R33043 VSS.n2858 VSS.n2857 2.25083
R33044 VSS.n4159 VSS.t48 2.24691
R33045 VSS.n3800 VSS.n3799 1.69274
R33046 VSS.n2108 VSS.n2107 1.63353
R33047 VSS.n3510 VSS.n771 1.63234
R33048 VSS.n2244 VSS.n2243 1.53355
R33049 VSS.n3798 VSS.n3797 1.3005
R33050 VSS.n3797 VSS.n3796 1.3005
R33051 VSS.n3800 VSS.n3558 1.21968
R33052 VSS.n3508 VSS.n774 1.19711
R33053 VSS.n3511 VSS.n3510 1.14563
R33054 VSS.n2107 VSS.n1659 0.983395
R33055 VSS.n4146 VSS.t44 0.936506
R33056 VSS.n2109 VSS.n2108 0.80221
R33057 VSS.n3799 VSS.n3798 0.785632
R33058 VSS.n3505 VSS.n771 0.664842
R33059 VSS.n3401 VSS.n3400 0.643325
R33060 VSS.n3798 VSS.n469 0.580763
R33061 VSS.n3386 VSS.n1030 0.57992
R33062 VSS.n4125 VSS.n470 0.578278
R33063 VSS.n713 VSS.n710 0.578278
R33064 VSS.n3799 VSS.n3559 0.578278
R33065 VSS.n3795 VSS.n3559 0.578278
R33066 VSS.n617 VSS.n616 0.578278
R33067 VSS.n3831 VSS.n3803 0.578278
R33068 VSS.n944 VSS.n894 0.578278
R33069 VSS.n773 VSS.n771 0.578278
R33070 VSS.n1738 VSS.n1703 0.578278
R33071 VSS.n1799 VSS.n1652 0.578278
R33072 VSS.n2097 VSS.n2096 0.578278
R33073 VSS.n1867 VSS.n1866 0.578278
R33074 VSS.n2128 VSS.n2127 0.578278
R33075 VSS.n1866 VSS.n1655 0.574928
R33076 VSS.n2127 VSS.n2126 0.574928
R33077 VSS.n4145 VSS.n470 0.574927
R33078 VSS.n616 VSS.n615 0.574927
R33079 VSS.n3423 VSS.n894 0.574927
R33080 VSS.n2186 VSS.n1652 0.574927
R33081 VSS.n3875 VSS.n3874 0.568921
R33082 VSS.t9 VSS.t28 0.562104
R33083 VSS.t3 VSS.t10 0.562104
R33084 VSS.t0 VSS.t26 0.562104
R33085 VSS.t6 VSS.t40 0.562104
R33086 VSS.n4027 VSS.n708 0.562104
R33087 VSS.n4161 VSS.t11 0.5465
R33088 VSS.n4161 VSS.t27 0.5465
R33089 VSS.n4163 VSS.t21 0.5465
R33090 VSS.n4163 VSS.t29 0.5465
R33091 VSS.n4165 VSS.t37 0.5465
R33092 VSS.n4165 VSS.t43 0.5465
R33093 VSS.n4167 VSS.t31 0.5465
R33094 VSS.n4167 VSS.t17 0.5465
R33095 VSS.n4169 VSS.t45 0.5465
R33096 VSS.n4169 VSS.t23 0.5465
R33097 VSS.n4171 VSS.t19 0.5465
R33098 VSS.n4171 VSS.t39 0.5465
R33099 VSS.n4173 VSS.t25 0.5465
R33100 VSS.n4173 VSS.t33 0.5465
R33101 VSS.n4175 VSS.t35 0.5465
R33102 VSS.n4175 VSS.t47 0.5465
R33103 VSS.n4177 VSS.t15 0.5465
R33104 VSS.n4177 VSS.t49 0.5465
R33105 VSS.n710 VSS.n709 0.545303
R33106 VSS.n3803 VSS.n3802 0.545303
R33107 VSS.n3507 VSS.n773 0.545303
R33108 VSS.n1754 VSS.n1703 0.545303
R33109 VSS.n2098 VSS.n2097 0.545303
R33110 VSS.n3404 VSS.n3403 0.473227
R33111 VSS.n3405 VSS.n3404 0.473227
R33112 VSS.n3407 VSS.n3406 0.473227
R33113 VSS.n3406 VSS.n3405 0.473227
R33114 VSS.n3187 VSS.n1405 0.459182
R33115 VSS.n4030 VSS.n4029 0.433833
R33116 VSS.n4029 VSS.n4028 0.433833
R33117 VSS.n1759 VSS.n1758 0.433833
R33118 VSS.n1758 VSS.n775 0.433833
R33119 VSS.n1701 VSS.n1700 0.433833
R33120 VSS.n1701 VSS.n775 0.433833
R33121 VSS.n2108 VSS.n1619 0.433833
R33122 VSS.n2239 VSS.n1619 0.433833
R33123 VSS.n1939 VSS.n1621 0.433833
R33124 VSS.n2239 VSS.n1621 0.433833
R33125 VSS.n2238 VSS.n2237 0.433833
R33126 VSS.n2239 VSS.n2238 0.433833
R33127 VSS.n3205 VSS.n1376 0.411087
R33128 VSS.n1820 VSS.n1687 0.38975
R33129 VSS.n1822 VSS.n1821 0.38975
R33130 VSS.n1823 VSS.n1683 0.38975
R33131 VSS.n1825 VSS.n1824 0.38975
R33132 VSS.n1724 VSS.n1685 0.38975
R33133 VSS.n1725 VSS.n1723 0.38975
R33134 VSS.n1727 VSS.n1726 0.38975
R33135 VSS.n1714 VSS.n1713 0.38975
R33136 VSS.n1736 VSS.n1735 0.38975
R33137 VSS.n1737 VSS.n1712 0.38975
R33138 VSS.n1740 VSS.n1739 0.38975
R33139 VSS.n1705 VSS.n1704 0.38975
R33140 VSS.n1751 VSS.n1750 0.38975
R33141 VSS.n3491 VSS.n801 0.374
R33142 VSS.n3492 VSS.n799 0.374
R33143 VSS.n3493 VSS.n797 0.374
R33144 VSS.n3494 VSS.n795 0.374
R33145 VSS.n3495 VSS.n793 0.374
R33146 VSS.n3496 VSS.n791 0.374
R33147 VSS.n3497 VSS.n789 0.374
R33148 VSS.n3498 VSS.n787 0.374
R33149 VSS.n3499 VSS.n785 0.374
R33150 VSS.n3500 VSS.n783 0.374
R33151 VSS.n3501 VSS.n778 0.374
R33152 VSS.n3503 VSS.n3502 0.374
R33153 VSS.n3417 VSS.n901 0.374
R33154 VSS.n3416 VSS.n902 0.374
R33155 VSS.n3415 VSS.n903 0.374
R33156 VSS.n3413 VSS.n904 0.374
R33157 VSS.n3412 VSS.n905 0.374
R33158 VSS.n3411 VSS.n906 0.374
R33159 VSS.n3410 VSS.n907 0.374
R33160 VSS.n3409 VSS.n908 0.374
R33161 VSS.n3408 VSS.n909 0.374
R33162 VSS.n1014 VSS.n910 0.374
R33163 VSS.n1013 VSS.n1012 0.374
R33164 VSS.n3418 VSS.n900 0.362917
R33165 VSS.n3780 VSS.n3778 0.361
R33166 VSS.n1379 VSS.n1376 0.3605
R33167 VSS.n1381 VSS.n1379 0.3605
R33168 VSS.n1383 VSS.n1381 0.3605
R33169 VSS.n1385 VSS.n1383 0.3605
R33170 VSS.n1387 VSS.n1385 0.3605
R33171 VSS.n1389 VSS.n1387 0.3605
R33172 VSS.n1391 VSS.n1389 0.3605
R33173 VSS.n1395 VSS.n1393 0.3605
R33174 VSS.n1397 VSS.n1395 0.3605
R33175 VSS.n1399 VSS.n1397 0.3605
R33176 VSS.n1401 VSS.n1399 0.3605
R33177 VSS.n1403 VSS.n1401 0.3605
R33178 VSS.n1405 VSS.n1403 0.3605
R33179 VSS.n4033 VSS.n594 0.35825
R33180 VSS.n4032 VSS.n592 0.35825
R33181 VSS.n4031 VSS.n590 0.35825
R33182 VSS.n605 VSS.n588 0.35825
R33183 VSS.n689 VSS.n586 0.35825
R33184 VSS.n690 VSS.n584 0.35825
R33185 VSS.n691 VSS.n582 0.35825
R33186 VSS.n692 VSS.n580 0.35825
R33187 VSS.n693 VSS.n578 0.35825
R33188 VSS.n694 VSS.n576 0.35825
R33189 VSS.n695 VSS.n574 0.35825
R33190 VSS.n696 VSS.n572 0.35825
R33191 VSS.n697 VSS.n570 0.35825
R33192 VSS.n698 VSS.n568 0.35825
R33193 VSS.n699 VSS.n566 0.35825
R33194 VSS.n700 VSS.n564 0.35825
R33195 VSS.n701 VSS.n562 0.35825
R33196 VSS.n702 VSS.n560 0.35825
R33197 VSS.n688 VSS.n558 0.35825
R33198 VSS.n687 VSS.n556 0.35825
R33199 VSS.n686 VSS.n554 0.35825
R33200 VSS.n685 VSS.n552 0.35825
R33201 VSS.n684 VSS.n550 0.35825
R33202 VSS.n683 VSS.n548 0.35825
R33203 VSS.n682 VSS.n546 0.35825
R33204 VSS.n681 VSS.n544 0.35825
R33205 VSS.n680 VSS.n542 0.35825
R33206 VSS.n679 VSS.n540 0.35825
R33207 VSS.n678 VSS.n538 0.35825
R33208 VSS.n677 VSS.n536 0.35825
R33209 VSS.n1760 VSS.n768 0.35375
R33210 VSS.n676 VSS.n607 0.34925
R33211 VSS.n674 VSS.n673 0.34925
R33212 VSS.n672 VSS.n608 0.34925
R33213 VSS.n618 VSS.n610 0.34925
R33214 VSS.n660 VSS.n659 0.34925
R33215 VSS.n658 VSS.n614 0.34925
R33216 VSS.n657 VSS.n619 0.34925
R33217 VSS.n656 VSS.n655 0.34925
R33218 VSS.n654 VSS.n620 0.34925
R33219 VSS.n628 VSS.n622 0.34925
R33220 VSS.n645 VSS.n644 0.34925
R33221 VSS.n643 VSS.n626 0.34925
R33222 VSS.n642 VSS.n634 0.34925
R33223 VSS.n641 VSS.n501 0.347
R33224 VSS.n640 VSS.n499 0.347
R33225 VSS.n639 VSS.n497 0.347
R33226 VSS.n638 VSS.n495 0.347
R33227 VSS.n637 VSS.n493 0.347
R33228 VSS.n636 VSS.n491 0.347
R33229 VSS.n635 VSS.n489 0.347
R33230 VSS.n487 VSS.n460 0.347
R33231 VSS.n4156 VSS.n461 0.347
R33232 VSS.n4155 VSS.n462 0.347
R33233 VSS.n4154 VSS.n463 0.347
R33234 VSS.n4153 VSS.n464 0.347
R33235 VSS.n4152 VSS.n4151 0.347
R33236 VSS.n4150 VSS.n465 0.347
R33237 VSS.n3644 VSS.n3622 0.345779
R33238 VSS.n2240 VSS.n1433 0.334713
R33239 VSS.n3996 VSS.n3898 0.33125
R33240 VSS.n3995 VSS.n3899 0.33125
R33241 VSS.n3994 VSS.n3900 0.33125
R33242 VSS.n3993 VSS.n3901 0.33125
R33243 VSS.n3992 VSS.n3902 0.33125
R33244 VSS.n3991 VSS.n3903 0.33125
R33245 VSS.n4000 VSS.n3896 0.33125
R33246 VSS.n4001 VSS.n3894 0.33125
R33247 VSS.n4002 VSS.n3892 0.33125
R33248 VSS.n4003 VSS.n3890 0.33125
R33249 VSS.n4004 VSS.n3888 0.33125
R33250 VSS.n4005 VSS.n3886 0.33125
R33251 VSS.n4006 VSS.n3884 0.33125
R33252 VSS.n4007 VSS.n3878 0.33125
R33253 VSS.n3514 VSS.n769 0.33125
R33254 VSS.n780 VSS.n777 0.33125
R33255 VSS.n770 VSS.n765 0.33125
R33256 VSS.n3519 VSS.n764 0.33125
R33257 VSS.n3520 VSS.n763 0.33125
R33258 VSS.n3521 VSS.n762 0.33125
R33259 VSS.n3522 VSS.n761 0.33125
R33260 VSS.n3523 VSS.n760 0.33125
R33261 VSS.n3524 VSS.n759 0.33125
R33262 VSS.n3525 VSS.n758 0.33125
R33263 VSS.n3526 VSS.n757 0.33125
R33264 VSS.n3527 VSS.n756 0.33125
R33265 VSS.n3528 VSS.n755 0.33125
R33266 VSS.n1771 VSS.n1689 0.33125
R33267 VSS.n1770 VSS.n1690 0.33125
R33268 VSS.n1769 VSS.n1691 0.33125
R33269 VSS.n1768 VSS.n1692 0.33125
R33270 VSS.n1767 VSS.n1693 0.33125
R33271 VSS.n1766 VSS.n1694 0.33125
R33272 VSS.n1765 VSS.n1695 0.33125
R33273 VSS.n1764 VSS.n1696 0.33125
R33274 VSS.n1763 VSS.n1697 0.33125
R33275 VSS.n1762 VSS.n1761 0.33125
R33276 VSS.n3999 VSS.n3998 0.33125
R33277 VSS.n3187 VSS.n3186 0.328273
R33278 VSS.n1757 VSS.n1692 0.3255
R33279 VSS.n1757 VSS.n1756 0.3255
R33280 VSS.n1702 VSS.n795 0.3255
R33281 VSS.n1756 VSS.n1702 0.3255
R33282 VSS.n2107 VSS.n2106 0.3255
R33283 VSS.n2106 VSS.n1618 0.3255
R33284 VSS.n1926 VSS.n1925 0.3255
R33285 VSS.n1925 VSS.n1618 0.3255
R33286 VSS.n2197 VSS.n1622 0.3255
R33287 VSS.n1622 VSS.n1618 0.3255
R33288 VSS.n3990 VSS.n3989 0.3245
R33289 VSS.n3988 VSS.n3904 0.3245
R33290 VSS.n3908 VSS.n3907 0.3245
R33291 VSS.n474 VSS.n472 0.3245
R33292 VSS.n4142 VSS.n4141 0.3245
R33293 VSS.n4140 VSS.n473 0.3245
R33294 VSS.n4119 VSS.n476 0.3245
R33295 VSS.n4123 VSS.n4122 0.3245
R33296 VSS.n4124 VSS.n4118 0.3245
R33297 VSS.n4127 VSS.n4126 0.3245
R33298 VSS.n468 VSS.n467 0.3245
R33299 VSS.n4150 VSS.n4149 0.3245
R33300 VSS.n3529 VSS.n754 0.320764
R33301 VSS.n3644 VSS.n3643 0.319973
R33302 VSS.n3780 VSS.n3779 0.316
R33303 VSS.n1773 VSS.n1772 0.311
R33304 VSS.n893 VSS.n892 0.306382
R33305 VSS.n896 VSS.n893 0.306382
R33306 VSS.n3414 VSS.n897 0.306382
R33307 VSS.n897 VSS.n896 0.306382
R33308 VSS.n469 VSS.n465 0.294184
R33309 VSS.n1772 VSS.n1771 0.29325
R33310 VSS.n1182 VSS.n1181 0.292176
R33311 VSS.n3513 VSS.n3512 0.2885
R33312 VSS.n2211 VSS.n2193 0.287346
R33313 VSS.n2233 VSS.n1630 0.28625
R33314 VSS.n2234 VSS.n1625 0.28625
R33315 VSS.n2236 VSS.n2235 0.28625
R33316 VSS.n1627 VSS.n1624 0.28625
R33317 VSS.n2203 VSS.n2202 0.28625
R33318 VSS.n2204 VSS.n2201 0.28625
R33319 VSS.n2205 VSS.n2200 0.28625
R33320 VSS.n2206 VSS.n2199 0.28625
R33321 VSS.n2207 VSS.n2198 0.28625
R33322 VSS.n2208 VSS.n2196 0.28625
R33323 VSS.n2209 VSS.n2195 0.28625
R33324 VSS.n2210 VSS.n2194 0.28625
R33325 VSS.n2192 VSS.n2191 0.284711
R33326 VSS.n2191 VSS.n2190 0.284711
R33327 VSS.n2190 VSS.n2189 0.284711
R33328 VSS.n1794 VSS.n1651 0.284711
R33329 VSS.n1795 VSS.n1794 0.284711
R33330 VSS.n1796 VSS.n1795 0.284711
R33331 VSS.n1797 VSS.n1796 0.284711
R33332 VSS.n1800 VSS.n1797 0.284711
R33333 VSS.n1798 VSS.n1658 0.284711
R33334 VSS.n4144 VSS.n4143 0.274184
R33335 VSS.n4026 VSS.n4025 0.274184
R33336 VSS.n4027 VSS.n4026 0.274184
R33337 VSS.n627 VSS.n458 0.274184
R33338 VSS.n3852 VSS.n3851 0.274184
R33339 VSS.n3852 VSS.n708 0.274184
R33340 VSS.n3425 VSS.n3424 0.274184
R33341 VSS.n3510 VSS.n3509 0.274184
R33342 VSS.n3509 VSS.n3508 0.274184
R33343 VSS.n1698 VSS.n1686 0.274184
R33344 VSS.n1755 VSS.n1698 0.274184
R33345 VSS.n2188 VSS.n2187 0.274184
R33346 VSS.n2077 VSS.n1623 0.274184
R33347 VSS.n1623 VSS.n1620 0.274184
R33348 VSS.n1881 VSS.n1880 0.274184
R33349 VSS.n2125 VSS.n2124 0.274184
R33350 VSS.n1880 VSS.n1655 0.27286
R33351 VSS.n2126 VSS.n2125 0.27286
R33352 VSS.n2187 VSS.n2186 0.27286
R33353 VSS.n3424 VSS.n3423 0.27286
R33354 VSS.n615 VSS.n458 0.27286
R33355 VSS.n4145 VSS.n4144 0.27286
R33356 VSS.n664 VSS.n525 0.2705
R33357 VSS.n666 VSS.n664 0.2705
R33358 VSS.n666 VSS.n665 0.2705
R33359 VSS.n668 VSS.n524 0.2705
R33360 VSS.n668 VSS.n667 0.2705
R33361 VSS.n667 VSS.n607 0.2705
R33362 VSS.n669 VSS.n523 0.2705
R33363 VSS.n669 VSS.n609 0.2705
R33364 VSS.n673 VSS.n609 0.2705
R33365 VSS.n670 VSS.n522 0.2705
R33366 VSS.n671 VSS.n670 0.2705
R33367 VSS.n672 VSS.n671 0.2705
R33368 VSS.n663 VSS.n521 0.2705
R33369 VSS.n663 VSS.n611 0.2705
R33370 VSS.n611 VSS.n610 0.2705
R33371 VSS.n662 VSS.n520 0.2705
R33372 VSS.n662 VSS.n661 0.2705
R33373 VSS.n661 VSS.n660 0.2705
R33374 VSS.n612 VSS.n519 0.2705
R33375 VSS.n613 VSS.n612 0.2705
R33376 VSS.n614 VSS.n613 0.2705
R33377 VSS.n650 VSS.n518 0.2705
R33378 VSS.n650 VSS.n649 0.2705
R33379 VSS.n649 VSS.n619 0.2705
R33380 VSS.n651 VSS.n517 0.2705
R33381 VSS.n651 VSS.n621 0.2705
R33382 VSS.n655 VSS.n621 0.2705
R33383 VSS.n652 VSS.n516 0.2705
R33384 VSS.n653 VSS.n652 0.2705
R33385 VSS.n654 VSS.n653 0.2705
R33386 VSS.n648 VSS.n515 0.2705
R33387 VSS.n648 VSS.n623 0.2705
R33388 VSS.n623 VSS.n622 0.2705
R33389 VSS.n647 VSS.n514 0.2705
R33390 VSS.n647 VSS.n646 0.2705
R33391 VSS.n646 VSS.n645 0.2705
R33392 VSS.n624 VSS.n513 0.2705
R33393 VSS.n625 VSS.n624 0.2705
R33394 VSS.n626 VSS.n625 0.2705
R33395 VSS.n631 VSS.n511 0.2705
R33396 VSS.n631 VSS.n630 0.2705
R33397 VSS.n630 VSS.n629 0.2705
R33398 VSS.n632 VSS.n512 0.2705
R33399 VSS.n633 VSS.n632 0.2705
R33400 VSS.n634 VSS.n633 0.2705
R33401 VSS.n3918 VSS.n3914 0.2705
R33402 VSS.n3920 VSS.n3918 0.2705
R33403 VSS.n3920 VSS.n3905 0.2705
R33404 VSS.n3913 VSS.n3911 0.2705
R33405 VSS.n3911 VSS.n3906 0.2705
R33406 VSS.n3989 VSS.n3906 0.2705
R33407 VSS.n3986 VSS.n3985 0.2705
R33408 VSS.n3987 VSS.n3986 0.2705
R33409 VSS.n3988 VSS.n3987 0.2705
R33410 VSS.n3912 VSS.n3910 0.2705
R33411 VSS.n3910 VSS.n3909 0.2705
R33412 VSS.n3909 VSS.n3908 0.2705
R33413 VSS.n3981 VSS.n3980 0.2705
R33414 VSS.n3980 VSS.n3979 0.2705
R33415 VSS.n3979 VSS.n474 0.2705
R33416 VSS.n481 VSS.n479 0.2705
R33417 VSS.n479 VSS.n475 0.2705
R33418 VSS.n4141 VSS.n475 0.2705
R33419 VSS.n4138 VSS.n4137 0.2705
R33420 VSS.n4139 VSS.n4138 0.2705
R33421 VSS.n4140 VSS.n4139 0.2705
R33422 VSS.n480 VSS.n478 0.2705
R33423 VSS.n478 VSS.n477 0.2705
R33424 VSS.n477 VSS.n476 0.2705
R33425 VSS.n4120 VSS.n483 0.2705
R33426 VSS.n4121 VSS.n4120 0.2705
R33427 VSS.n4122 VSS.n4121 0.2705
R33428 VSS.n4116 VSS.n484 0.2705
R33429 VSS.n4117 VSS.n4116 0.2705
R33430 VSS.n4118 VSS.n4117 0.2705
R33431 VSS.n4130 VSS.n4129 0.2705
R33432 VSS.n4129 VSS.n4128 0.2705
R33433 VSS.n4128 VSS.n4127 0.2705
R33434 VSS.n4100 VSS.n4099 0.2705
R33435 VSS.n4101 VSS.n4100 0.2705
R33436 VSS.n4102 VSS.n4101 0.2705
R33437 VSS.n4103 VSS.n4102 0.2705
R33438 VSS.n4104 VSS.n4103 0.2705
R33439 VSS.n4105 VSS.n4104 0.2705
R33440 VSS.n4106 VSS.n4105 0.2705
R33441 VSS.n4107 VSS.n4106 0.2705
R33442 VSS.n4108 VSS.n4107 0.2705
R33443 VSS.n4109 VSS.n4108 0.2705
R33444 VSS.n4110 VSS.n4109 0.2705
R33445 VSS.n4111 VSS.n4110 0.2705
R33446 VSS.n4112 VSS.n4111 0.2705
R33447 VSS.n4113 VSS.n4112 0.2705
R33448 VSS.n4114 VSS.n4113 0.2705
R33449 VSS.n4115 VSS.n4114 0.2705
R33450 VSS.n4115 VSS.n466 0.2705
R33451 VSS.n467 VSS.n466 0.2705
R33452 VSS.n4098 VSS.n509 0.2705
R33453 VSS.n509 VSS.n507 0.2705
R33454 VSS.n507 VSS.n505 0.2705
R33455 VSS.n505 VSS.n503 0.2705
R33456 VSS.n503 VSS.n501 0.2705
R33457 VSS.n501 VSS.n499 0.2705
R33458 VSS.n499 VSS.n497 0.2705
R33459 VSS.n497 VSS.n495 0.2705
R33460 VSS.n495 VSS.n493 0.2705
R33461 VSS.n493 VSS.n491 0.2705
R33462 VSS.n491 VSS.n489 0.2705
R33463 VSS.n489 VSS.n487 0.2705
R33464 VSS.n487 VSS.n461 0.2705
R33465 VSS.n462 VSS.n461 0.2705
R33466 VSS.n463 VSS.n462 0.2705
R33467 VSS.n464 VSS.n463 0.2705
R33468 VSS.n4151 VSS.n464 0.2705
R33469 VSS.n4151 VSS.n4150 0.2705
R33470 VSS.n950 VSS.n877 0.2705
R33471 VSS.n951 VSS.n950 0.2705
R33472 VSS.n734 VSS.n732 0.2705
R33473 VSS.n735 VSS.n734 0.2705
R33474 VSS.n3430 VSS.n3429 0.2705
R33475 VSS.n3429 VSS.n3428 0.2705
R33476 VSS.n888 VSS.n887 0.2705
R33477 VSS.n889 VSS.n888 0.2705
R33478 VSS.n932 VSS.n886 0.2705
R33479 VSS.n933 VSS.n932 0.2705
R33480 VSS.n931 VSS.n885 0.2705
R33481 VSS.n934 VSS.n931 0.2705
R33482 VSS.n938 VSS.n884 0.2705
R33483 VSS.n938 VSS.n937 0.2705
R33484 VSS.n939 VSS.n883 0.2705
R33485 VSS.n939 VSS.n929 0.2705
R33486 VSS.n940 VSS.n882 0.2705
R33487 VSS.n941 VSS.n940 0.2705
R33488 VSS.n930 VSS.n881 0.2705
R33489 VSS.n930 VSS.n927 0.2705
R33490 VSS.n926 VSS.n880 0.2705
R33491 VSS.n946 VSS.n926 0.2705
R33492 VSS.n948 VSS.n879 0.2705
R33493 VSS.n948 VSS.n947 0.2705
R33494 VSS.n949 VSS.n878 0.2705
R33495 VSS.n949 VSS.n899 0.2705
R33496 VSS.n3534 VSS.n3533 0.2705
R33497 VSS.n3533 VSS.n3532 0.2705
R33498 VSS.n719 VSS.n718 0.2705
R33499 VSS.n720 VSS.n719 0.2705
R33500 VSS.n721 VSS.n720 0.2705
R33501 VSS.n722 VSS.n721 0.2705
R33502 VSS.n723 VSS.n722 0.2705
R33503 VSS.n724 VSS.n723 0.2705
R33504 VSS.n725 VSS.n724 0.2705
R33505 VSS.n726 VSS.n725 0.2705
R33506 VSS.n727 VSS.n726 0.2705
R33507 VSS.n728 VSS.n727 0.2705
R33508 VSS.n730 VSS.n728 0.2705
R33509 VSS.n731 VSS.n730 0.2705
R33510 VSS.n733 VSS.n731 0.2705
R33511 VSS.n3531 VSS.n733 0.2705
R33512 VSS.n745 VSS.n744 0.2705
R33513 VSS.n746 VSS.n745 0.2705
R33514 VSS.n747 VSS.n746 0.2705
R33515 VSS.n748 VSS.n747 0.2705
R33516 VSS.n749 VSS.n748 0.2705
R33517 VSS.n750 VSS.n749 0.2705
R33518 VSS.n751 VSS.n750 0.2705
R33519 VSS.n752 VSS.n751 0.2705
R33520 VSS.n753 VSS.n752 0.2705
R33521 VSS.n3530 VSS.n753 0.2705
R33522 VSS.n3529 VSS.n3528 0.2705
R33523 VSS.n3528 VSS.n3527 0.2705
R33524 VSS.n3527 VSS.n3526 0.2705
R33525 VSS.n3526 VSS.n3525 0.2705
R33526 VSS.n3525 VSS.n3524 0.2705
R33527 VSS.n3524 VSS.n3523 0.2705
R33528 VSS.n3523 VSS.n3522 0.2705
R33529 VSS.n3522 VSS.n3521 0.2705
R33530 VSS.n3521 VSS.n3520 0.2705
R33531 VSS.n3520 VSS.n3519 0.2705
R33532 VSS.n3519 VSS.n765 0.2705
R33533 VSS.n3513 VSS.n765 0.2705
R33534 VSS.n3514 VSS.n3513 0.2705
R33535 VSS.n767 VSS.n766 0.2705
R33536 VSS.n3515 VSS.n767 0.2705
R33537 VSS.n1763 VSS.n1762 0.2705
R33538 VSS.n1764 VSS.n1763 0.2705
R33539 VSS.n1765 VSS.n1764 0.2705
R33540 VSS.n1766 VSS.n1765 0.2705
R33541 VSS.n1767 VSS.n1766 0.2705
R33542 VSS.n1768 VSS.n1767 0.2705
R33543 VSS.n1769 VSS.n1768 0.2705
R33544 VSS.n1770 VSS.n1769 0.2705
R33545 VSS.n1771 VSS.n1770 0.2705
R33546 VSS.n1774 VSS.n1773 0.2705
R33547 VSS.n1775 VSS.n1774 0.2705
R33548 VSS.n1776 VSS.n1775 0.2705
R33549 VSS.n1777 VSS.n1776 0.2705
R33550 VSS.n1778 VSS.n1777 0.2705
R33551 VSS.n1779 VSS.n1778 0.2705
R33552 VSS.n1780 VSS.n1779 0.2705
R33553 VSS.n1781 VSS.n1780 0.2705
R33554 VSS.n1782 VSS.n1781 0.2705
R33555 VSS.n1858 VSS.n1854 0.2705
R33556 VSS.n1860 VSS.n1858 0.2705
R33557 VSS.n1862 VSS.n1860 0.2705
R33558 VSS.n1918 VSS.n1862 0.2705
R33559 VSS.n1897 VSS.n1853 0.2705
R33560 VSS.n1897 VSS.n1896 0.2705
R33561 VSS.n1896 VSS.n1865 0.2705
R33562 VSS.n1916 VSS.n1865 0.2705
R33563 VSS.n1898 VSS.n1852 0.2705
R33564 VSS.n1898 VSS.n1868 0.2705
R33565 VSS.n1914 VSS.n1868 0.2705
R33566 VSS.n1915 VSS.n1914 0.2705
R33567 VSS.n1899 VSS.n1851 0.2705
R33568 VSS.n1899 VSS.n1870 0.2705
R33569 VSS.n1913 VSS.n1870 0.2705
R33570 VSS.n1913 VSS.n1912 0.2705
R33571 VSS.n1900 VSS.n1850 0.2705
R33572 VSS.n1901 VSS.n1900 0.2705
R33573 VSS.n1901 VSS.n1869 0.2705
R33574 VSS.n1911 VSS.n1869 0.2705
R33575 VSS.n1903 VSS.n1849 0.2705
R33576 VSS.n1903 VSS.n1902 0.2705
R33577 VSS.n1902 VSS.n1871 0.2705
R33578 VSS.n1910 VSS.n1871 0.2705
R33579 VSS.n1904 VSS.n1848 0.2705
R33580 VSS.n1904 VSS.n1873 0.2705
R33581 VSS.n1908 VSS.n1873 0.2705
R33582 VSS.n1909 VSS.n1908 0.2705
R33583 VSS.n1905 VSS.n1847 0.2705
R33584 VSS.n1906 VSS.n1905 0.2705
R33585 VSS.n1907 VSS.n1906 0.2705
R33586 VSS.n1907 VSS.n1872 0.2705
R33587 VSS.n1895 VSS.n1846 0.2705
R33588 VSS.n1895 VSS.n1875 0.2705
R33589 VSS.n1875 VSS.n1874 0.2705
R33590 VSS.n1879 VSS.n1874 0.2705
R33591 VSS.n1894 VSS.n1845 0.2705
R33592 VSS.n1894 VSS.n1893 0.2705
R33593 VSS.n1893 VSS.n1892 0.2705
R33594 VSS.n1892 VSS.n1891 0.2705
R33595 VSS.n1876 VSS.n1844 0.2705
R33596 VSS.n1877 VSS.n1876 0.2705
R33597 VSS.n1878 VSS.n1877 0.2705
R33598 VSS.n1890 VSS.n1878 0.2705
R33599 VSS.n1885 VSS.n1843 0.2705
R33600 VSS.n1886 VSS.n1885 0.2705
R33601 VSS.n1887 VSS.n1886 0.2705
R33602 VSS.n1889 VSS.n1887 0.2705
R33603 VSS.n1884 VSS.n1842 0.2705
R33604 VSS.n1884 VSS.n1882 0.2705
R33605 VSS.n1882 VSS.n1660 0.2705
R33606 VSS.n1888 VSS.n1660 0.2705
R33607 VSS.n1883 VSS.n1841 0.2705
R33608 VSS.n1883 VSS.n1661 0.2705
R33609 VSS.n2181 VSS.n1661 0.2705
R33610 VSS.n1667 VSS.n1663 0.2705
R33611 VSS.n2179 VSS.n1663 0.2705
R33612 VSS.n2180 VSS.n2179 0.2705
R33613 VSS.n2177 VSS.n2176 0.2705
R33614 VSS.n2178 VSS.n2177 0.2705
R33615 VSS.n2178 VSS.n1662 0.2705
R33616 VSS.n1970 VSS.n1969 0.2705
R33617 VSS.n1971 VSS.n1970 0.2705
R33618 VSS.n1972 VSS.n1971 0.2705
R33619 VSS.n1973 VSS.n1972 0.2705
R33620 VSS.n1974 VSS.n1973 0.2705
R33621 VSS.n1975 VSS.n1974 0.2705
R33622 VSS.n1976 VSS.n1975 0.2705
R33623 VSS.n1977 VSS.n1976 0.2705
R33624 VSS.n1978 VSS.n1977 0.2705
R33625 VSS.n1979 VSS.n1978 0.2705
R33626 VSS.n1980 VSS.n1979 0.2705
R33627 VSS.n1981 VSS.n1980 0.2705
R33628 VSS.n1982 VSS.n1981 0.2705
R33629 VSS.n1983 VSS.n1982 0.2705
R33630 VSS.n1984 VSS.n1983 0.2705
R33631 VSS.n1985 VSS.n1984 0.2705
R33632 VSS.n1986 VSS.n1985 0.2705
R33633 VSS.n1987 VSS.n1986 0.2705
R33634 VSS.n1988 VSS.n1987 0.2705
R33635 VSS.n1857 VSS.n1856 0.2705
R33636 VSS.n1859 VSS.n1857 0.2705
R33637 VSS.n1861 VSS.n1859 0.2705
R33638 VSS.n1863 VSS.n1861 0.2705
R33639 VSS.n1864 VSS.n1863 0.2705
R33640 VSS.n1920 VSS.n1864 0.2705
R33641 VSS.n1922 VSS.n1920 0.2705
R33642 VSS.n1924 VSS.n1922 0.2705
R33643 VSS.n1928 VSS.n1924 0.2705
R33644 VSS.n1930 VSS.n1928 0.2705
R33645 VSS.n1932 VSS.n1930 0.2705
R33646 VSS.n1934 VSS.n1932 0.2705
R33647 VSS.n1936 VSS.n1934 0.2705
R33648 VSS.n1938 VSS.n1936 0.2705
R33649 VSS.n1941 VSS.n1938 0.2705
R33650 VSS.n1943 VSS.n1941 0.2705
R33651 VSS.n1946 VSS.n1943 0.2705
R33652 VSS.n1948 VSS.n1946 0.2705
R33653 VSS.n1949 VSS.n1948 0.2705
R33654 VSS.n2157 VSS.n2156 0.2705
R33655 VSS.n2156 VSS.n2155 0.2705
R33656 VSS.n2155 VSS.n2154 0.2705
R33657 VSS.n2154 VSS.n2153 0.2705
R33658 VSS.n2153 VSS.n2152 0.2705
R33659 VSS.n2152 VSS.n2151 0.2705
R33660 VSS.n2151 VSS.n2150 0.2705
R33661 VSS.n2150 VSS.n2149 0.2705
R33662 VSS.n2149 VSS.n2148 0.2705
R33663 VSS.n2148 VSS.n2147 0.2705
R33664 VSS.n2147 VSS.n2146 0.2705
R33665 VSS.n2146 VSS.n2145 0.2705
R33666 VSS.n2145 VSS.n2144 0.2705
R33667 VSS.n2144 VSS.n2143 0.2705
R33668 VSS.n2143 VSS.n2142 0.2705
R33669 VSS.n2142 VSS.n2141 0.2705
R33670 VSS.n2141 VSS.n2140 0.2705
R33671 VSS.n2140 VSS.n2139 0.2705
R33672 VSS.n2139 VSS.n2138 0.2705
R33673 VSS.n1947 VSS.n1945 0.2705
R33674 VSS.n2137 VSS.n1947 0.2705
R33675 VSS.n2001 VSS.n1995 0.2705
R33676 VSS.n1995 VSS.n1992 0.2705
R33677 VSS.n2132 VSS.n1996 0.2705
R33678 VSS.n2133 VSS.n2132 0.2705
R33679 VSS.n2131 VSS.n2130 0.2705
R33680 VSS.n2131 VSS.n1994 0.2705
R33681 VSS.n1998 VSS.n1997 0.2705
R33682 VSS.n2015 VSS.n1997 0.2705
R33683 VSS.n2020 VSS.n2019 0.2705
R33684 VSS.n2019 VSS.n2018 0.2705
R33685 VSS.n2024 VSS.n2023 0.2705
R33686 VSS.n2025 VSS.n2024 0.2705
R33687 VSS.n2011 VSS.n2010 0.2705
R33688 VSS.n2026 VSS.n2011 0.2705
R33689 VSS.n2122 VSS.n2121 0.2705
R33690 VSS.n2121 VSS.n2012 0.2705
R33691 VSS.n2120 VSS.n2009 0.2705
R33692 VSS.n2120 VSS.n2119 0.2705
R33693 VSS.n2102 VSS.n2013 0.2705
R33694 VSS.n2118 VSS.n2013 0.2705
R33695 VSS.n2103 VSS.n2033 0.2705
R33696 VSS.n2033 VSS.n2030 0.2705
R33697 VSS.n2113 VSS.n2034 0.2705
R33698 VSS.n2114 VSS.n2113 0.2705
R33699 VSS.n2112 VSS.n2111 0.2705
R33700 VSS.n2112 VSS.n2032 0.2705
R33701 VSS.n2036 VSS.n2035 0.2705
R33702 VSS.n2046 VSS.n2035 0.2705
R33703 VSS.n2042 VSS.n2041 0.2705
R33704 VSS.n2047 VSS.n2042 0.2705
R33705 VSS.n2095 VSS.n2094 0.2705
R33706 VSS.n2094 VSS.n2043 0.2705
R33707 VSS.n2093 VSS.n2040 0.2705
R33708 VSS.n2093 VSS.n2092 0.2705
R33709 VSS.n2079 VSS.n2044 0.2705
R33710 VSS.n2091 VSS.n2044 0.2705
R33711 VSS.n2080 VSS.n2054 0.2705
R33712 VSS.n2054 VSS.n2051 0.2705
R33713 VSS.n2086 VSS.n2055 0.2705
R33714 VSS.n2087 VSS.n2086 0.2705
R33715 VSS.n2085 VSS.n2084 0.2705
R33716 VSS.n2085 VSS.n2053 0.2705
R33717 VSS.n2057 VSS.n2056 0.2705
R33718 VSS.n2061 VSS.n2056 0.2705
R33719 VSS.n2074 VSS.n2073 0.2705
R33720 VSS.n2073 VSS.n2072 0.2705
R33721 VSS.n2060 VSS.n2059 0.2705
R33722 VSS.n2071 VSS.n2060 0.2705
R33723 VSS.n2066 VSS.n2065 0.2705
R33724 VSS.n2067 VSS.n2066 0.2705
R33725 VSS.n1634 VSS.n1632 0.2705
R33726 VSS.n1635 VSS.n1634 0.2705
R33727 VSS.n2211 VSS.n2210 0.2705
R33728 VSS.n2210 VSS.n2209 0.2705
R33729 VSS.n2209 VSS.n2208 0.2705
R33730 VSS.n2208 VSS.n2207 0.2705
R33731 VSS.n2207 VSS.n2206 0.2705
R33732 VSS.n2206 VSS.n2205 0.2705
R33733 VSS.n2205 VSS.n2204 0.2705
R33734 VSS.n2204 VSS.n2203 0.2705
R33735 VSS.n2203 VSS.n1627 0.2705
R33736 VSS.n2235 VSS.n1627 0.2705
R33737 VSS.n2235 VSS.n2234 0.2705
R33738 VSS.n2234 VSS.n2233 0.2705
R33739 VSS.n2233 VSS.n2232 0.2705
R33740 VSS.n2232 VSS.n2231 0.2705
R33741 VSS.n2231 VSS.n2230 0.2705
R33742 VSS.n2212 VSS.n1645 0.2705
R33743 VSS.n1645 VSS.n1644 0.2705
R33744 VSS.n1644 VSS.n1643 0.2705
R33745 VSS.n1643 VSS.n1642 0.2705
R33746 VSS.n1642 VSS.n1641 0.2705
R33747 VSS.n1641 VSS.n1640 0.2705
R33748 VSS.n1640 VSS.n1639 0.2705
R33749 VSS.n1639 VSS.n1638 0.2705
R33750 VSS.n1638 VSS.n1637 0.2705
R33751 VSS.n1637 VSS.n1626 0.2705
R33752 VSS.n1628 VSS.n1626 0.2705
R33753 VSS.n1629 VSS.n1628 0.2705
R33754 VSS.n1631 VSS.n1629 0.2705
R33755 VSS.n1633 VSS.n1631 0.2705
R33756 VSS.n2229 VSS.n1633 0.2705
R33757 VSS.n1647 VSS.n1646 0.2705
R33758 VSS.n1818 VSS.n1688 0.2705
R33759 VSS.n1818 VSS.n1817 0.2705
R33760 VSS.n1817 VSS.n1816 0.2705
R33761 VSS.n1816 VSS.n1815 0.2705
R33762 VSS.n1815 VSS.n1814 0.2705
R33763 VSS.n1814 VSS.n1813 0.2705
R33764 VSS.n1813 VSS.n1812 0.2705
R33765 VSS.n1812 VSS.n1811 0.2705
R33766 VSS.n1811 VSS.n1810 0.2705
R33767 VSS.n1810 VSS.n1809 0.2705
R33768 VSS.n1809 VSS.n1808 0.2705
R33769 VSS.n1808 VSS.n1807 0.2705
R33770 VSS.n1807 VSS.n1806 0.2705
R33771 VSS.n1806 VSS.n1805 0.2705
R33772 VSS.n1805 VSS.n1804 0.2705
R33773 VSS.n1804 VSS.n1803 0.2705
R33774 VSS.n1803 VSS.n1802 0.2705
R33775 VSS.n1820 VSS.n1819 0.2705
R33776 VSS.n1819 VSS.n1680 0.2705
R33777 VSS.n1680 VSS.n1679 0.2705
R33778 VSS.n1679 VSS.n1677 0.2705
R33779 VSS.n1677 VSS.n1676 0.2705
R33780 VSS.n1676 VSS.n1675 0.2705
R33781 VSS.n1675 VSS.n1674 0.2705
R33782 VSS.n1674 VSS.n1673 0.2705
R33783 VSS.n1673 VSS.n1672 0.2705
R33784 VSS.n1672 VSS.n1671 0.2705
R33785 VSS.n1671 VSS.n1670 0.2705
R33786 VSS.n1670 VSS.n1669 0.2705
R33787 VSS.n1669 VSS.n1668 0.2705
R33788 VSS.n1668 VSS.n1666 0.2705
R33789 VSS.n1666 VSS.n1665 0.2705
R33790 VSS.n1665 VSS.n1664 0.2705
R33791 VSS.n1801 VSS.n1664 0.2705
R33792 VSS.n1821 VSS.n1681 0.2705
R33793 VSS.n1829 VSS.n1681 0.2705
R33794 VSS.n1827 VSS.n1683 0.2705
R33795 VSS.n1828 VSS.n1827 0.2705
R33796 VSS.n1826 VSS.n1825 0.2705
R33797 VSS.n1826 VSS.n1682 0.2705
R33798 VSS.n1685 VSS.n1684 0.2705
R33799 VSS.n1720 VSS.n1684 0.2705
R33800 VSS.n1723 VSS.n1722 0.2705
R33801 VSS.n1722 VSS.n1721 0.2705
R33802 VSS.n1728 VSS.n1727 0.2705
R33803 VSS.n1729 VSS.n1728 0.2705
R33804 VSS.n1715 VSS.n1714 0.2705
R33805 VSS.n1716 VSS.n1715 0.2705
R33806 VSS.n1735 VSS.n1734 0.2705
R33807 VSS.n1734 VSS.n1733 0.2705
R33808 VSS.n1712 VSS.n1711 0.2705
R33809 VSS.n1711 VSS.n1710 0.2705
R33810 VSS.n1741 VSS.n1740 0.2705
R33811 VSS.n1742 VSS.n1741 0.2705
R33812 VSS.n1706 VSS.n1705 0.2705
R33813 VSS.n1707 VSS.n1706 0.2705
R33814 VSS.n1750 VSS.n1749 0.2705
R33815 VSS.n1749 VSS.n1748 0.2705
R33816 VSS.n805 VSS.n804 0.2705
R33817 VSS.n1708 VSS.n805 0.2705
R33818 VSS.n925 VSS.n876 0.2705
R33819 VSS.n952 VSS.n925 0.2705
R33820 VSS.n952 VSS.n900 0.2705
R33821 VSS.n901 VSS.n900 0.2705
R33822 VSS.n902 VSS.n901 0.2705
R33823 VSS.n903 VSS.n902 0.2705
R33824 VSS.n904 VSS.n903 0.2705
R33825 VSS.n905 VSS.n904 0.2705
R33826 VSS.n906 VSS.n905 0.2705
R33827 VSS.n907 VSS.n906 0.2705
R33828 VSS.n908 VSS.n907 0.2705
R33829 VSS.n909 VSS.n908 0.2705
R33830 VSS.n910 VSS.n909 0.2705
R33831 VSS.n1012 VSS.n910 0.2705
R33832 VSS.n1012 VSS.n780 0.2705
R33833 VSS.n3502 VSS.n780 0.2705
R33834 VSS.n3502 VSS.n3501 0.2705
R33835 VSS.n3501 VSS.n3500 0.2705
R33836 VSS.n3500 VSS.n3499 0.2705
R33837 VSS.n3499 VSS.n3498 0.2705
R33838 VSS.n3498 VSS.n3497 0.2705
R33839 VSS.n3497 VSS.n3496 0.2705
R33840 VSS.n3496 VSS.n3495 0.2705
R33841 VSS.n3495 VSS.n3494 0.2705
R33842 VSS.n3494 VSS.n3493 0.2705
R33843 VSS.n3493 VSS.n3492 0.2705
R33844 VSS.n3492 VSS.n3491 0.2705
R33845 VSS.n3491 VSS.n3490 0.2705
R33846 VSS.n3490 VSS.n3489 0.2705
R33847 VSS.n3489 VSS.n3488 0.2705
R33848 VSS.n3488 VSS.n806 0.2705
R33849 VSS.n964 VSS.n875 0.2705
R33850 VSS.n964 VSS.n963 0.2705
R33851 VSS.n963 VSS.n962 0.2705
R33852 VSS.n962 VSS.n961 0.2705
R33853 VSS.n961 VSS.n960 0.2705
R33854 VSS.n960 VSS.n959 0.2705
R33855 VSS.n959 VSS.n958 0.2705
R33856 VSS.n958 VSS.n957 0.2705
R33857 VSS.n957 VSS.n956 0.2705
R33858 VSS.n956 VSS.n955 0.2705
R33859 VSS.n955 VSS.n954 0.2705
R33860 VSS.n954 VSS.n953 0.2705
R33861 VSS.n953 VSS.n912 0.2705
R33862 VSS.n1011 VSS.n912 0.2705
R33863 VSS.n1011 VSS.n1010 0.2705
R33864 VSS.n1010 VSS.n779 0.2705
R33865 VSS.n781 VSS.n779 0.2705
R33866 VSS.n782 VSS.n781 0.2705
R33867 VSS.n784 VSS.n782 0.2705
R33868 VSS.n786 VSS.n784 0.2705
R33869 VSS.n788 VSS.n786 0.2705
R33870 VSS.n790 VSS.n788 0.2705
R33871 VSS.n792 VSS.n790 0.2705
R33872 VSS.n794 VSS.n792 0.2705
R33873 VSS.n796 VSS.n794 0.2705
R33874 VSS.n798 VSS.n796 0.2705
R33875 VSS.n800 VSS.n798 0.2705
R33876 VSS.n802 VSS.n800 0.2705
R33877 VSS.n803 VSS.n802 0.2705
R33878 VSS.n3487 VSS.n803 0.2705
R33879 VSS.n3487 VSS.n3486 0.2705
R33880 VSS.n965 VSS.n874 0.2705
R33881 VSS.n965 VSS.n924 0.2705
R33882 VSS.n924 VSS.n923 0.2705
R33883 VSS.n923 VSS.n922 0.2705
R33884 VSS.n922 VSS.n921 0.2705
R33885 VSS.n921 VSS.n920 0.2705
R33886 VSS.n920 VSS.n919 0.2705
R33887 VSS.n919 VSS.n918 0.2705
R33888 VSS.n918 VSS.n917 0.2705
R33889 VSS.n917 VSS.n916 0.2705
R33890 VSS.n916 VSS.n915 0.2705
R33891 VSS.n915 VSS.n914 0.2705
R33892 VSS.n914 VSS.n913 0.2705
R33893 VSS.n913 VSS.n911 0.2705
R33894 VSS.n1009 VSS.n911 0.2705
R33895 VSS.n1009 VSS.n1008 0.2705
R33896 VSS.n1008 VSS.n1007 0.2705
R33897 VSS.n1007 VSS.n1006 0.2705
R33898 VSS.n1006 VSS.n1005 0.2705
R33899 VSS.n1005 VSS.n1004 0.2705
R33900 VSS.n1004 VSS.n1003 0.2705
R33901 VSS.n1003 VSS.n1002 0.2705
R33902 VSS.n1002 VSS.n1001 0.2705
R33903 VSS.n1001 VSS.n1000 0.2705
R33904 VSS.n1000 VSS.n999 0.2705
R33905 VSS.n999 VSS.n998 0.2705
R33906 VSS.n998 VSS.n997 0.2705
R33907 VSS.n997 VSS.n996 0.2705
R33908 VSS.n996 VSS.n995 0.2705
R33909 VSS.n995 VSS.n807 0.2705
R33910 VSS.n3485 VSS.n807 0.2705
R33911 VSS.n966 VSS.n873 0.2705
R33912 VSS.n967 VSS.n966 0.2705
R33913 VSS.n968 VSS.n967 0.2705
R33914 VSS.n969 VSS.n968 0.2705
R33915 VSS.n970 VSS.n969 0.2705
R33916 VSS.n971 VSS.n970 0.2705
R33917 VSS.n972 VSS.n971 0.2705
R33918 VSS.n973 VSS.n972 0.2705
R33919 VSS.n974 VSS.n973 0.2705
R33920 VSS.n975 VSS.n974 0.2705
R33921 VSS.n976 VSS.n975 0.2705
R33922 VSS.n977 VSS.n976 0.2705
R33923 VSS.n978 VSS.n977 0.2705
R33924 VSS.n979 VSS.n978 0.2705
R33925 VSS.n980 VSS.n979 0.2705
R33926 VSS.n981 VSS.n980 0.2705
R33927 VSS.n982 VSS.n981 0.2705
R33928 VSS.n983 VSS.n982 0.2705
R33929 VSS.n984 VSS.n983 0.2705
R33930 VSS.n985 VSS.n984 0.2705
R33931 VSS.n986 VSS.n985 0.2705
R33932 VSS.n987 VSS.n986 0.2705
R33933 VSS.n988 VSS.n987 0.2705
R33934 VSS.n989 VSS.n988 0.2705
R33935 VSS.n990 VSS.n989 0.2705
R33936 VSS.n991 VSS.n990 0.2705
R33937 VSS.n992 VSS.n991 0.2705
R33938 VSS.n993 VSS.n992 0.2705
R33939 VSS.n994 VSS.n993 0.2705
R33940 VSS.n994 VSS.n812 0.2705
R33941 VSS.n812 VSS.n809 0.2705
R33942 VSS.n3448 VSS.n871 0.2705
R33943 VSS.n871 VSS.n869 0.2705
R33944 VSS.n869 VSS.n867 0.2705
R33945 VSS.n867 VSS.n865 0.2705
R33946 VSS.n865 VSS.n863 0.2705
R33947 VSS.n863 VSS.n861 0.2705
R33948 VSS.n861 VSS.n859 0.2705
R33949 VSS.n859 VSS.n857 0.2705
R33950 VSS.n857 VSS.n855 0.2705
R33951 VSS.n855 VSS.n853 0.2705
R33952 VSS.n853 VSS.n851 0.2705
R33953 VSS.n851 VSS.n849 0.2705
R33954 VSS.n849 VSS.n847 0.2705
R33955 VSS.n847 VSS.n845 0.2705
R33956 VSS.n845 VSS.n843 0.2705
R33957 VSS.n843 VSS.n841 0.2705
R33958 VSS.n841 VSS.n839 0.2705
R33959 VSS.n839 VSS.n837 0.2705
R33960 VSS.n837 VSS.n835 0.2705
R33961 VSS.n835 VSS.n833 0.2705
R33962 VSS.n833 VSS.n831 0.2705
R33963 VSS.n831 VSS.n829 0.2705
R33964 VSS.n829 VSS.n827 0.2705
R33965 VSS.n827 VSS.n825 0.2705
R33966 VSS.n825 VSS.n823 0.2705
R33967 VSS.n823 VSS.n821 0.2705
R33968 VSS.n821 VSS.n819 0.2705
R33969 VSS.n819 VSS.n817 0.2705
R33970 VSS.n817 VSS.n813 0.2705
R33971 VSS.n3480 VSS.n813 0.2705
R33972 VSS.n3481 VSS.n3480 0.2705
R33973 VSS.n3450 VSS.n3449 0.2705
R33974 VSS.n3451 VSS.n3450 0.2705
R33975 VSS.n3452 VSS.n3451 0.2705
R33976 VSS.n3453 VSS.n3452 0.2705
R33977 VSS.n3454 VSS.n3453 0.2705
R33978 VSS.n3455 VSS.n3454 0.2705
R33979 VSS.n3456 VSS.n3455 0.2705
R33980 VSS.n3457 VSS.n3456 0.2705
R33981 VSS.n3458 VSS.n3457 0.2705
R33982 VSS.n3459 VSS.n3458 0.2705
R33983 VSS.n3460 VSS.n3459 0.2705
R33984 VSS.n3461 VSS.n3460 0.2705
R33985 VSS.n3462 VSS.n3461 0.2705
R33986 VSS.n3463 VSS.n3462 0.2705
R33987 VSS.n3464 VSS.n3463 0.2705
R33988 VSS.n3465 VSS.n3464 0.2705
R33989 VSS.n3466 VSS.n3465 0.2705
R33990 VSS.n3467 VSS.n3466 0.2705
R33991 VSS.n3468 VSS.n3467 0.2705
R33992 VSS.n3469 VSS.n3468 0.2705
R33993 VSS.n3470 VSS.n3469 0.2705
R33994 VSS.n3471 VSS.n3470 0.2705
R33995 VSS.n3472 VSS.n3471 0.2705
R33996 VSS.n3473 VSS.n3472 0.2705
R33997 VSS.n3474 VSS.n3473 0.2705
R33998 VSS.n3475 VSS.n3474 0.2705
R33999 VSS.n3476 VSS.n3475 0.2705
R34000 VSS.n3477 VSS.n3476 0.2705
R34001 VSS.n3478 VSS.n3477 0.2705
R34002 VSS.n3479 VSS.n3478 0.2705
R34003 VSS.n3479 VSS.n811 0.2705
R34004 VSS.n3871 VSS.n714 0.2705
R34005 VSS.n3871 VSS.n3870 0.2705
R34006 VSS.n3858 VSS.n716 0.2705
R34007 VSS.n3869 VSS.n716 0.2705
R34008 VSS.n3553 VSS.n3550 0.2705
R34009 VSS.n3865 VSS.n3864 0.2705
R34010 VSS.n3863 VSS.n3862 0.2705
R34011 VSS.n3863 VSS.n3552 0.2705
R34012 VSS.n3556 VSS.n3555 0.2705
R34013 VSS.n3812 VSS.n3555 0.2705
R34014 VSS.n3808 VSS.n3807 0.2705
R34015 VSS.n3813 VSS.n3808 0.2705
R34016 VSS.n3849 VSS.n3848 0.2705
R34017 VSS.n3848 VSS.n3809 0.2705
R34018 VSS.n3847 VSS.n3806 0.2705
R34019 VSS.n3847 VSS.n3846 0.2705
R34020 VSS.n3833 VSS.n3810 0.2705
R34021 VSS.n3845 VSS.n3810 0.2705
R34022 VSS.n3834 VSS.n3820 0.2705
R34023 VSS.n3820 VSS.n3817 0.2705
R34024 VSS.n3840 VSS.n3821 0.2705
R34025 VSS.n3841 VSS.n3840 0.2705
R34026 VSS.n3839 VSS.n3838 0.2705
R34027 VSS.n3839 VSS.n3819 0.2705
R34028 VSS.n3828 VSS.n3827 0.2705
R34029 VSS.n3827 VSS.n3822 0.2705
R34030 VSS.n3826 VSS.n603 0.2705
R34031 VSS.n3826 VSS.n3825 0.2705
R34032 VSS.n4035 VSS.n602 0.2705
R34033 VSS.n602 VSS.n601 0.2705
R34034 VSS.n4037 VSS.n4036 0.2705
R34035 VSS.n4038 VSS.n4037 0.2705
R34036 VSS.n528 VSS.n526 0.2705
R34037 VSS.n530 VSS.n528 0.2705
R34038 VSS.n532 VSS.n530 0.2705
R34039 VSS.n534 VSS.n532 0.2705
R34040 VSS.n536 VSS.n534 0.2705
R34041 VSS.n538 VSS.n536 0.2705
R34042 VSS.n540 VSS.n538 0.2705
R34043 VSS.n542 VSS.n540 0.2705
R34044 VSS.n544 VSS.n542 0.2705
R34045 VSS.n546 VSS.n544 0.2705
R34046 VSS.n548 VSS.n546 0.2705
R34047 VSS.n550 VSS.n548 0.2705
R34048 VSS.n552 VSS.n550 0.2705
R34049 VSS.n554 VSS.n552 0.2705
R34050 VSS.n556 VSS.n554 0.2705
R34051 VSS.n558 VSS.n556 0.2705
R34052 VSS.n560 VSS.n558 0.2705
R34053 VSS.n562 VSS.n560 0.2705
R34054 VSS.n564 VSS.n562 0.2705
R34055 VSS.n566 VSS.n564 0.2705
R34056 VSS.n568 VSS.n566 0.2705
R34057 VSS.n570 VSS.n568 0.2705
R34058 VSS.n572 VSS.n570 0.2705
R34059 VSS.n574 VSS.n572 0.2705
R34060 VSS.n576 VSS.n574 0.2705
R34061 VSS.n578 VSS.n576 0.2705
R34062 VSS.n580 VSS.n578 0.2705
R34063 VSS.n582 VSS.n580 0.2705
R34064 VSS.n584 VSS.n582 0.2705
R34065 VSS.n586 VSS.n584 0.2705
R34066 VSS.n588 VSS.n586 0.2705
R34067 VSS.n590 VSS.n588 0.2705
R34068 VSS.n592 VSS.n590 0.2705
R34069 VSS.n594 VSS.n592 0.2705
R34070 VSS.n596 VSS.n594 0.2705
R34071 VSS.n597 VSS.n596 0.2705
R34072 VSS.n599 VSS.n597 0.2705
R34073 VSS.n4079 VSS.n4078 0.2705
R34074 VSS.n4078 VSS.n4077 0.2705
R34075 VSS.n4077 VSS.n4076 0.2705
R34076 VSS.n4076 VSS.n4075 0.2705
R34077 VSS.n4075 VSS.n4074 0.2705
R34078 VSS.n4074 VSS.n4073 0.2705
R34079 VSS.n4073 VSS.n4072 0.2705
R34080 VSS.n4072 VSS.n4071 0.2705
R34081 VSS.n4071 VSS.n4070 0.2705
R34082 VSS.n4070 VSS.n4069 0.2705
R34083 VSS.n4069 VSS.n4068 0.2705
R34084 VSS.n4068 VSS.n4067 0.2705
R34085 VSS.n4067 VSS.n4066 0.2705
R34086 VSS.n4066 VSS.n4065 0.2705
R34087 VSS.n4065 VSS.n4064 0.2705
R34088 VSS.n4064 VSS.n4063 0.2705
R34089 VSS.n4063 VSS.n4062 0.2705
R34090 VSS.n4062 VSS.n4061 0.2705
R34091 VSS.n4061 VSS.n4060 0.2705
R34092 VSS.n4060 VSS.n4059 0.2705
R34093 VSS.n4059 VSS.n4058 0.2705
R34094 VSS.n4058 VSS.n4057 0.2705
R34095 VSS.n4057 VSS.n4056 0.2705
R34096 VSS.n4056 VSS.n4055 0.2705
R34097 VSS.n4055 VSS.n4054 0.2705
R34098 VSS.n4054 VSS.n4053 0.2705
R34099 VSS.n4053 VSS.n4052 0.2705
R34100 VSS.n4052 VSS.n4051 0.2705
R34101 VSS.n4051 VSS.n4050 0.2705
R34102 VSS.n4050 VSS.n4049 0.2705
R34103 VSS.n4049 VSS.n4048 0.2705
R34104 VSS.n4048 VSS.n4047 0.2705
R34105 VSS.n4047 VSS.n4046 0.2705
R34106 VSS.n4046 VSS.n4045 0.2705
R34107 VSS.n4045 VSS.n4044 0.2705
R34108 VSS.n4044 VSS.n4043 0.2705
R34109 VSS.n4043 VSS.n4042 0.2705
R34110 VSS.n3931 VSS.n3930 0.2705
R34111 VSS.n3930 VSS.n3929 0.2705
R34112 VSS.n3929 VSS.n3928 0.2705
R34113 VSS.n3928 VSS.n3922 0.2705
R34114 VSS.n3923 VSS.n3922 0.2705
R34115 VSS.n3924 VSS.n3923 0.2705
R34116 VSS.n3925 VSS.n3924 0.2705
R34117 VSS.n3926 VSS.n3925 0.2705
R34118 VSS.n3927 VSS.n3926 0.2705
R34119 VSS.n3963 VSS.n3927 0.2705
R34120 VSS.n3963 VSS.n3962 0.2705
R34121 VSS.n3962 VSS.n3961 0.2705
R34122 VSS.n3961 VSS.n3960 0.2705
R34123 VSS.n3960 VSS.n3959 0.2705
R34124 VSS.n3959 VSS.n3958 0.2705
R34125 VSS.n3958 VSS.n3957 0.2705
R34126 VSS.n3957 VSS.n3956 0.2705
R34127 VSS.n3956 VSS.n3955 0.2705
R34128 VSS.n3955 VSS.n3954 0.2705
R34129 VSS.n3954 VSS.n3953 0.2705
R34130 VSS.n3917 VSS.n3916 0.2705
R34131 VSS.n3919 VSS.n3917 0.2705
R34132 VSS.n3921 VSS.n3919 0.2705
R34133 VSS.n3970 VSS.n3921 0.2705
R34134 VSS.n3970 VSS.n3969 0.2705
R34135 VSS.n3969 VSS.n3968 0.2705
R34136 VSS.n3968 VSS.n3967 0.2705
R34137 VSS.n3967 VSS.n3966 0.2705
R34138 VSS.n3966 VSS.n3965 0.2705
R34139 VSS.n3965 VSS.n3964 0.2705
R34140 VSS.n3964 VSS.n3897 0.2705
R34141 VSS.n3897 VSS.n3895 0.2705
R34142 VSS.n3895 VSS.n3893 0.2705
R34143 VSS.n3893 VSS.n3891 0.2705
R34144 VSS.n3891 VSS.n3889 0.2705
R34145 VSS.n3889 VSS.n3887 0.2705
R34146 VSS.n3887 VSS.n3885 0.2705
R34147 VSS.n3885 VSS.n3883 0.2705
R34148 VSS.n3883 VSS.n3882 0.2705
R34149 VSS.n3882 VSS.n3881 0.2705
R34150 VSS.n3975 VSS.n3974 0.2705
R34151 VSS.n3974 VSS.n3973 0.2705
R34152 VSS.n3973 VSS.n3972 0.2705
R34153 VSS.n3972 VSS.n3971 0.2705
R34154 VSS.n3971 VSS.n3903 0.2705
R34155 VSS.n3903 VSS.n3902 0.2705
R34156 VSS.n3902 VSS.n3901 0.2705
R34157 VSS.n3901 VSS.n3900 0.2705
R34158 VSS.n3900 VSS.n3899 0.2705
R34159 VSS.n3899 VSS.n3898 0.2705
R34160 VSS.n3999 VSS.n3898 0.2705
R34161 VSS.n4000 VSS.n3999 0.2705
R34162 VSS.n4001 VSS.n4000 0.2705
R34163 VSS.n4002 VSS.n4001 0.2705
R34164 VSS.n4003 VSS.n4002 0.2705
R34165 VSS.n4004 VSS.n4003 0.2705
R34166 VSS.n4005 VSS.n4004 0.2705
R34167 VSS.n4006 VSS.n4005 0.2705
R34168 VSS.n4007 VSS.n4006 0.2705
R34169 VSS.n4008 VSS.n4007 0.2705
R34170 VSS.n1205 VSS.n1170 0.2705
R34171 VSS.n1170 VSS.n1166 0.2705
R34172 VSS.n1204 VSS.n1203 0.2705
R34173 VSS.n1203 VSS.n1165 0.2705
R34174 VSS.n1202 VSS.n1172 0.2705
R34175 VSS.n1202 VSS.n1164 0.2705
R34176 VSS.n1201 VSS.n1200 0.2705
R34177 VSS.n1201 VSS.n1163 0.2705
R34178 VSS.n1199 VSS.n1173 0.2705
R34179 VSS.n1173 VSS.n1162 0.2705
R34180 VSS.n1198 VSS.n1197 0.2705
R34181 VSS.n1197 VSS.n1161 0.2705
R34182 VSS.n1196 VSS.n1174 0.2705
R34183 VSS.n1196 VSS.n1160 0.2705
R34184 VSS.n1195 VSS.n1194 0.2705
R34185 VSS.n1195 VSS.n1159 0.2705
R34186 VSS.n1193 VSS.n1175 0.2705
R34187 VSS.n1175 VSS.n1158 0.2705
R34188 VSS.n1192 VSS.n1191 0.2705
R34189 VSS.n1191 VSS.n1157 0.2705
R34190 VSS.n1190 VSS.n1176 0.2705
R34191 VSS.n1190 VSS.n1156 0.2705
R34192 VSS.n1189 VSS.n1188 0.2705
R34193 VSS.n1189 VSS.n1155 0.2705
R34194 VSS.n1187 VSS.n1177 0.2705
R34195 VSS.n1177 VSS.n1154 0.2705
R34196 VSS.n1186 VSS.n1185 0.2705
R34197 VSS.n1185 VSS.n1153 0.2705
R34198 VSS.n1184 VSS.n1178 0.2705
R34199 VSS.n1184 VSS.n1152 0.2705
R34200 VSS.n1183 VSS.n1182 0.2705
R34201 VSS.n1183 VSS.n1151 0.2705
R34202 VSS.n1179 VSS.n1150 0.2705
R34203 VSS.n1373 VSS.n1372 0.2705
R34204 VSS.n1374 VSS.n1373 0.2705
R34205 VSS.n1362 VSS.n1361 0.2705
R34206 VSS.n1363 VSS.n1362 0.2705
R34207 VSS.n1364 VSS.n1363 0.2705
R34208 VSS.n1365 VSS.n1364 0.2705
R34209 VSS.n1366 VSS.n1365 0.2705
R34210 VSS.n1367 VSS.n1366 0.2705
R34211 VSS.n1368 VSS.n1367 0.2705
R34212 VSS.n1369 VSS.n1368 0.2705
R34213 VSS.n1370 VSS.n1369 0.2705
R34214 VSS.n3214 VSS.n1370 0.2705
R34215 VSS.n3213 VSS.n3212 0.2705
R34216 VSS.n3212 VSS.n3211 0.2705
R34217 VSS.n3211 VSS.n3210 0.2705
R34218 VSS.n1138 VSS.n1137 0.2705
R34219 VSS.n1137 VSS.n1136 0.2705
R34220 VSS.n1136 VSS.n1135 0.2705
R34221 VSS.n1135 VSS.n1134 0.2705
R34222 VSS.n1134 VSS.n1133 0.2705
R34223 VSS.n1133 VSS.n1132 0.2705
R34224 VSS.n1132 VSS.n1131 0.2705
R34225 VSS.n1131 VSS.n1130 0.2705
R34226 VSS.n1130 VSS.n1129 0.2705
R34227 VSS.n1129 VSS.n1128 0.2705
R34228 VSS.n1128 VSS.n1125 0.2705
R34229 VSS.n1126 VSS.n1125 0.2705
R34230 VSS.n1127 VSS.n1126 0.2705
R34231 VSS.n3215 VSS.n1127 0.2705
R34232 VSS.n3317 VSS.n3316 0.2705
R34233 VSS.n3316 VSS.n3216 0.2705
R34234 VSS.n3315 VSS.n1123 0.2705
R34235 VSS.n3315 VSS.n3314 0.2705
R34236 VSS.n3217 VSS.n1122 0.2705
R34237 VSS.n3313 VSS.n3217 0.2705
R34238 VSS.n3218 VSS.n1121 0.2705
R34239 VSS.n3312 VSS.n3218 0.2705
R34240 VSS.n3310 VSS.n1120 0.2705
R34241 VSS.n3311 VSS.n3310 0.2705
R34242 VSS.n3309 VSS.n1119 0.2705
R34243 VSS.n3309 VSS.n3219 0.2705
R34244 VSS.n3308 VSS.n1118 0.2705
R34245 VSS.n3308 VSS.n3220 0.2705
R34246 VSS.n3307 VSS.n1117 0.2705
R34247 VSS.n3307 VSS.n3306 0.2705
R34248 VSS.n3221 VSS.n1116 0.2705
R34249 VSS.n3305 VSS.n3221 0.2705
R34250 VSS.n3222 VSS.n1115 0.2705
R34251 VSS.n3304 VSS.n3222 0.2705
R34252 VSS.n3302 VSS.n1114 0.2705
R34253 VSS.n3303 VSS.n3302 0.2705
R34254 VSS.n3301 VSS.n1113 0.2705
R34255 VSS.n3301 VSS.n3223 0.2705
R34256 VSS.n3300 VSS.n1112 0.2705
R34257 VSS.n3300 VSS.n3224 0.2705
R34258 VSS.n3299 VSS.n1111 0.2705
R34259 VSS.n3299 VSS.n3298 0.2705
R34260 VSS.n3225 VSS.n1110 0.2705
R34261 VSS.n3297 VSS.n3225 0.2705
R34262 VSS.n3297 VSS.n3296 0.2705
R34263 VSS.n3296 VSS.n3295 0.2705
R34264 VSS.n3295 VSS.n3294 0.2705
R34265 VSS.n3294 VSS.n3293 0.2705
R34266 VSS.n3293 VSS.n1015 0.2705
R34267 VSS.n3399 VSS.n3398 0.2705
R34268 VSS.n3398 VSS.n3397 0.2705
R34269 VSS.n3397 VSS.n3396 0.2705
R34270 VSS.n3396 VSS.n3395 0.2705
R34271 VSS.n3395 VSS.n3394 0.2705
R34272 VSS.n3394 VSS.n3393 0.2705
R34273 VSS.n3393 VSS.n3392 0.2705
R34274 VSS.n3392 VSS.n3391 0.2705
R34275 VSS.n3391 VSS.n3390 0.2705
R34276 VSS.n3390 VSS.n3389 0.2705
R34277 VSS.n1439 VSS.n1435 0.2705
R34278 VSS.n3086 VSS.n1435 0.2705
R34279 VSS.n3087 VSS.n3086 0.2705
R34280 VSS.n3084 VSS.n3083 0.2705
R34281 VSS.n3085 VSS.n3084 0.2705
R34282 VSS.n3085 VSS.n1434 0.2705
R34283 VSS.n1438 VSS.n1437 0.2705
R34284 VSS.n1437 VSS.n1436 0.2705
R34285 VSS.n1525 VSS.n1436 0.2705
R34286 VSS.n1528 VSS.n1441 0.2705
R34287 VSS.n1528 VSS.n1527 0.2705
R34288 VSS.n1527 VSS.n1526 0.2705
R34289 VSS.n1603 VSS.n1602 0.2705
R34290 VSS.n1602 VSS.n1601 0.2705
R34291 VSS.n1601 VSS.n1600 0.2705
R34292 VSS.n1600 VSS.n1599 0.2705
R34293 VSS.n1599 VSS.n1598 0.2705
R34294 VSS.n1598 VSS.n1597 0.2705
R34295 VSS.n1597 VSS.n1596 0.2705
R34296 VSS.n1596 VSS.n1595 0.2705
R34297 VSS.n1595 VSS.n1594 0.2705
R34298 VSS.n1594 VSS.n1593 0.2705
R34299 VSS.n1593 VSS.n1592 0.2705
R34300 VSS.n1592 VSS.n1591 0.2705
R34301 VSS.n1591 VSS.n1509 0.2705
R34302 VSS.n2260 VSS.n1509 0.2705
R34303 VSS.n2261 VSS.n2260 0.2705
R34304 VSS.n2246 VSS.n2245 0.2705
R34305 VSS.n2247 VSS.n2246 0.2705
R34306 VSS.n2248 VSS.n2247 0.2705
R34307 VSS.n2249 VSS.n2248 0.2705
R34308 VSS.n2250 VSS.n2249 0.2705
R34309 VSS.n2251 VSS.n2250 0.2705
R34310 VSS.n2252 VSS.n2251 0.2705
R34311 VSS.n2253 VSS.n2252 0.2705
R34312 VSS.n2254 VSS.n2253 0.2705
R34313 VSS.n2255 VSS.n2254 0.2705
R34314 VSS.n2256 VSS.n2255 0.2705
R34315 VSS.n2257 VSS.n2256 0.2705
R34316 VSS.n2258 VSS.n2257 0.2705
R34317 VSS.n2259 VSS.n2258 0.2705
R34318 VSS.n2259 VSS.n1507 0.2705
R34319 VSS.n1590 VSS.n1510 0.2705
R34320 VSS.n1510 VSS.n1506 0.2705
R34321 VSS.n1589 VSS.n1588 0.2705
R34322 VSS.n1588 VSS.n1505 0.2705
R34323 VSS.n1587 VSS.n1511 0.2705
R34324 VSS.n1587 VSS.n1504 0.2705
R34325 VSS.n1586 VSS.n1585 0.2705
R34326 VSS.n1586 VSS.n1503 0.2705
R34327 VSS.n1584 VSS.n1512 0.2705
R34328 VSS.n1512 VSS.n1502 0.2705
R34329 VSS.n1583 VSS.n1582 0.2705
R34330 VSS.n1582 VSS.n1501 0.2705
R34331 VSS.n1581 VSS.n1513 0.2705
R34332 VSS.n1581 VSS.n1500 0.2705
R34333 VSS.n1580 VSS.n1579 0.2705
R34334 VSS.n1580 VSS.n1499 0.2705
R34335 VSS.n1578 VSS.n1514 0.2705
R34336 VSS.n1514 VSS.n1498 0.2705
R34337 VSS.n1577 VSS.n1576 0.2705
R34338 VSS.n1576 VSS.n1497 0.2705
R34339 VSS.n1575 VSS.n1515 0.2705
R34340 VSS.n1575 VSS.n1496 0.2705
R34341 VSS.n1574 VSS.n1573 0.2705
R34342 VSS.n1574 VSS.n1495 0.2705
R34343 VSS.n1572 VSS.n1516 0.2705
R34344 VSS.n1516 VSS.n1494 0.2705
R34345 VSS.n1571 VSS.n1570 0.2705
R34346 VSS.n1570 VSS.n1493 0.2705
R34347 VSS.n1569 VSS.n1517 0.2705
R34348 VSS.n1569 VSS.n1492 0.2705
R34349 VSS.n1568 VSS.n1567 0.2705
R34350 VSS.n1568 VSS.n1491 0.2705
R34351 VSS.n1566 VSS.n1518 0.2705
R34352 VSS.n1518 VSS.n1490 0.2705
R34353 VSS.n1565 VSS.n1564 0.2705
R34354 VSS.n1564 VSS.n1489 0.2705
R34355 VSS.n1563 VSS.n1519 0.2705
R34356 VSS.n1563 VSS.n1488 0.2705
R34357 VSS.n1562 VSS.n1561 0.2705
R34358 VSS.n1562 VSS.n1487 0.2705
R34359 VSS.n1560 VSS.n1520 0.2705
R34360 VSS.n1520 VSS.n1486 0.2705
R34361 VSS.n1559 VSS.n1558 0.2705
R34362 VSS.n1558 VSS.n1485 0.2705
R34363 VSS.n1557 VSS.n1521 0.2705
R34364 VSS.n1557 VSS.n1484 0.2705
R34365 VSS.n1556 VSS.n1555 0.2705
R34366 VSS.n1556 VSS.n1481 0.2705
R34367 VSS.n1554 VSS.n1523 0.2705
R34368 VSS.n1523 VSS.n1522 0.2705
R34369 VSS.n1553 VSS.n1552 0.2705
R34370 VSS.n1552 VSS.n1551 0.2705
R34371 VSS.n1549 VSS.n1524 0.2705
R34372 VSS.n1550 VSS.n1549 0.2705
R34373 VSS.n1529 VSS.n1442 0.2705
R34374 VSS.n1530 VSS.n1529 0.2705
R34375 VSS.n1531 VSS.n1530 0.2705
R34376 VSS.n1532 VSS.n1531 0.2705
R34377 VSS.n1533 VSS.n1532 0.2705
R34378 VSS.n1534 VSS.n1533 0.2705
R34379 VSS.n1535 VSS.n1534 0.2705
R34380 VSS.n1536 VSS.n1535 0.2705
R34381 VSS.n1537 VSS.n1536 0.2705
R34382 VSS.n1538 VSS.n1537 0.2705
R34383 VSS.n1539 VSS.n1538 0.2705
R34384 VSS.n1540 VSS.n1539 0.2705
R34385 VSS.n1541 VSS.n1540 0.2705
R34386 VSS.n1542 VSS.n1541 0.2705
R34387 VSS.n1543 VSS.n1542 0.2705
R34388 VSS.n1544 VSS.n1543 0.2705
R34389 VSS.n1545 VSS.n1544 0.2705
R34390 VSS.n1548 VSS.n1545 0.2705
R34391 VSS.n1548 VSS.n1547 0.2705
R34392 VSS.n1445 VSS.n1443 0.2705
R34393 VSS.n1447 VSS.n1445 0.2705
R34394 VSS.n1449 VSS.n1447 0.2705
R34395 VSS.n1451 VSS.n1449 0.2705
R34396 VSS.n1453 VSS.n1451 0.2705
R34397 VSS.n1455 VSS.n1453 0.2705
R34398 VSS.n1457 VSS.n1455 0.2705
R34399 VSS.n1459 VSS.n1457 0.2705
R34400 VSS.n1461 VSS.n1459 0.2705
R34401 VSS.n1463 VSS.n1461 0.2705
R34402 VSS.n1465 VSS.n1463 0.2705
R34403 VSS.n1467 VSS.n1465 0.2705
R34404 VSS.n1469 VSS.n1467 0.2705
R34405 VSS.n1471 VSS.n1469 0.2705
R34406 VSS.n1473 VSS.n1471 0.2705
R34407 VSS.n1475 VSS.n1473 0.2705
R34408 VSS.n1477 VSS.n1475 0.2705
R34409 VSS.n1478 VSS.n1477 0.2705
R34410 VSS.n1546 VSS.n1478 0.2705
R34411 VSS.n3076 VSS.n3075 0.2705
R34412 VSS.n3075 VSS.n3074 0.2705
R34413 VSS.n3074 VSS.n3073 0.2705
R34414 VSS.n3073 VSS.n3072 0.2705
R34415 VSS.n3072 VSS.n3071 0.2705
R34416 VSS.n3071 VSS.n3070 0.2705
R34417 VSS.n3070 VSS.n3069 0.2705
R34418 VSS.n3069 VSS.n3068 0.2705
R34419 VSS.n3068 VSS.n3067 0.2705
R34420 VSS.n3067 VSS.n3066 0.2705
R34421 VSS.n3066 VSS.n3065 0.2705
R34422 VSS.n3065 VSS.n3064 0.2705
R34423 VSS.n3064 VSS.n3063 0.2705
R34424 VSS.n3063 VSS.n3062 0.2705
R34425 VSS.n3062 VSS.n3061 0.2705
R34426 VSS.n3061 VSS.n3060 0.2705
R34427 VSS.n3060 VSS.n3059 0.2705
R34428 VSS.n3059 VSS.n3058 0.2705
R34429 VSS.n3058 VSS.n3057 0.2705
R34430 VSS.n3122 VSS.n3120 0.2705
R34431 VSS.n3168 VSS.n3120 0.2705
R34432 VSS.n3166 VSS.n3123 0.2705
R34433 VSS.n3167 VSS.n3166 0.2705
R34434 VSS.n3165 VSS.n3164 0.2705
R34435 VSS.n3165 VSS.n3121 0.2705
R34436 VSS.n3163 VSS.n3124 0.2705
R34437 VSS.n3127 VSS.n3124 0.2705
R34438 VSS.n3162 VSS.n3161 0.2705
R34439 VSS.n3161 VSS.n3160 0.2705
R34440 VSS.n3126 VSS.n3125 0.2705
R34441 VSS.n3159 VSS.n3126 0.2705
R34442 VSS.n3135 VSS.n3134 0.2705
R34443 VSS.n3134 VSS.n3131 0.2705
R34444 VSS.n3154 VSS.n3136 0.2705
R34445 VSS.n3155 VSS.n3154 0.2705
R34446 VSS.n3153 VSS.n3152 0.2705
R34447 VSS.n3153 VSS.n3133 0.2705
R34448 VSS.n3151 VSS.n3137 0.2705
R34449 VSS.n3140 VSS.n3137 0.2705
R34450 VSS.n3150 VSS.n3149 0.2705
R34451 VSS.n3149 VSS.n3148 0.2705
R34452 VSS.n3139 VSS.n3138 0.2705
R34453 VSS.n3147 VSS.n3139 0.2705
R34454 VSS.n1039 VSS.n1038 0.2705
R34455 VSS.n3143 VSS.n1039 0.2705
R34456 VSS.n3384 VSS.n3383 0.2705
R34457 VSS.n3383 VSS.n3382 0.2705
R34458 VSS.n3382 VSS.n3381 0.2705
R34459 VSS.n3381 VSS.n3380 0.2705
R34460 VSS.n3380 VSS.n3379 0.2705
R34461 VSS.n3379 VSS.n3378 0.2705
R34462 VSS.n3378 VSS.n1040 0.2705
R34463 VSS.n3236 VSS.n1109 0.2705
R34464 VSS.n3236 VSS.n3226 0.2705
R34465 VSS.n3227 VSS.n3226 0.2705
R34466 VSS.n3228 VSS.n3227 0.2705
R34467 VSS.n3229 VSS.n3228 0.2705
R34468 VSS.n3292 VSS.n3229 0.2705
R34469 VSS.n3292 VSS.n3291 0.2705
R34470 VSS.n3291 VSS.n3290 0.2705
R34471 VSS.n3247 VSS.n1017 0.2705
R34472 VSS.n1018 VSS.n1017 0.2705
R34473 VSS.n1019 VSS.n1018 0.2705
R34474 VSS.n1020 VSS.n1019 0.2705
R34475 VSS.n1021 VSS.n1020 0.2705
R34476 VSS.n1022 VSS.n1021 0.2705
R34477 VSS.n1023 VSS.n1022 0.2705
R34478 VSS.n1024 VSS.n1023 0.2705
R34479 VSS.n1025 VSS.n1024 0.2705
R34480 VSS.n1026 VSS.n1025 0.2705
R34481 VSS.n1027 VSS.n1026 0.2705
R34482 VSS.n1028 VSS.n1027 0.2705
R34483 VSS.n1029 VSS.n1028 0.2705
R34484 VSS.n1031 VSS.n1029 0.2705
R34485 VSS.n1032 VSS.n1031 0.2705
R34486 VSS.n1033 VSS.n1032 0.2705
R34487 VSS.n1034 VSS.n1033 0.2705
R34488 VSS.n1035 VSS.n1034 0.2705
R34489 VSS.n1036 VSS.n1035 0.2705
R34490 VSS.n1037 VSS.n1036 0.2705
R34491 VSS.n3377 VSS.n1037 0.2705
R34492 VSS.n3377 VSS.n3376 0.2705
R34493 VSS.n3237 VSS.n1108 0.2705
R34494 VSS.n3237 VSS.n3235 0.2705
R34495 VSS.n3235 VSS.n3234 0.2705
R34496 VSS.n3234 VSS.n3233 0.2705
R34497 VSS.n3233 VSS.n3232 0.2705
R34498 VSS.n3232 VSS.n3230 0.2705
R34499 VSS.n3231 VSS.n3230 0.2705
R34500 VSS.n3289 VSS.n3231 0.2705
R34501 VSS.n3289 VSS.n3288 0.2705
R34502 VSS.n3288 VSS.n3287 0.2705
R34503 VSS.n3287 VSS.n3286 0.2705
R34504 VSS.n3286 VSS.n3285 0.2705
R34505 VSS.n3285 VSS.n3284 0.2705
R34506 VSS.n3284 VSS.n3283 0.2705
R34507 VSS.n3283 VSS.n3282 0.2705
R34508 VSS.n3282 VSS.n3281 0.2705
R34509 VSS.n3281 VSS.n3280 0.2705
R34510 VSS.n3280 VSS.n3279 0.2705
R34511 VSS.n3279 VSS.n3278 0.2705
R34512 VSS.n3278 VSS.n3277 0.2705
R34513 VSS.n3277 VSS.n3276 0.2705
R34514 VSS.n3276 VSS.n3275 0.2705
R34515 VSS.n3275 VSS.n3274 0.2705
R34516 VSS.n3274 VSS.n3273 0.2705
R34517 VSS.n3273 VSS.n3272 0.2705
R34518 VSS.n3272 VSS.n3271 0.2705
R34519 VSS.n3271 VSS.n3270 0.2705
R34520 VSS.n3270 VSS.n3269 0.2705
R34521 VSS.n3269 VSS.n3268 0.2705
R34522 VSS.n3268 VSS.n1041 0.2705
R34523 VSS.n3375 VSS.n1041 0.2705
R34524 VSS.n3238 VSS.n1107 0.2705
R34525 VSS.n3239 VSS.n3238 0.2705
R34526 VSS.n3240 VSS.n3239 0.2705
R34527 VSS.n3241 VSS.n3240 0.2705
R34528 VSS.n3242 VSS.n3241 0.2705
R34529 VSS.n3243 VSS.n3242 0.2705
R34530 VSS.n3244 VSS.n3243 0.2705
R34531 VSS.n3245 VSS.n3244 0.2705
R34532 VSS.n3246 VSS.n3245 0.2705
R34533 VSS.n3248 VSS.n3246 0.2705
R34534 VSS.n3249 VSS.n3248 0.2705
R34535 VSS.n3250 VSS.n3249 0.2705
R34536 VSS.n3251 VSS.n3250 0.2705
R34537 VSS.n3252 VSS.n3251 0.2705
R34538 VSS.n3253 VSS.n3252 0.2705
R34539 VSS.n3254 VSS.n3253 0.2705
R34540 VSS.n3255 VSS.n3254 0.2705
R34541 VSS.n3256 VSS.n3255 0.2705
R34542 VSS.n3257 VSS.n3256 0.2705
R34543 VSS.n3258 VSS.n3257 0.2705
R34544 VSS.n3259 VSS.n3258 0.2705
R34545 VSS.n3260 VSS.n3259 0.2705
R34546 VSS.n3261 VSS.n3260 0.2705
R34547 VSS.n3262 VSS.n3261 0.2705
R34548 VSS.n3263 VSS.n3262 0.2705
R34549 VSS.n3264 VSS.n3263 0.2705
R34550 VSS.n3265 VSS.n3264 0.2705
R34551 VSS.n3266 VSS.n3265 0.2705
R34552 VSS.n3267 VSS.n3266 0.2705
R34553 VSS.n3267 VSS.n1046 0.2705
R34554 VSS.n1046 VSS.n1043 0.2705
R34555 VSS.n3338 VSS.n1105 0.2705
R34556 VSS.n1105 VSS.n1103 0.2705
R34557 VSS.n1103 VSS.n1101 0.2705
R34558 VSS.n1101 VSS.n1099 0.2705
R34559 VSS.n1099 VSS.n1097 0.2705
R34560 VSS.n1097 VSS.n1095 0.2705
R34561 VSS.n1095 VSS.n1093 0.2705
R34562 VSS.n1093 VSS.n1091 0.2705
R34563 VSS.n1091 VSS.n1089 0.2705
R34564 VSS.n1089 VSS.n1087 0.2705
R34565 VSS.n1087 VSS.n1085 0.2705
R34566 VSS.n1085 VSS.n1083 0.2705
R34567 VSS.n1083 VSS.n1081 0.2705
R34568 VSS.n1081 VSS.n1079 0.2705
R34569 VSS.n1079 VSS.n1077 0.2705
R34570 VSS.n1077 VSS.n1075 0.2705
R34571 VSS.n1075 VSS.n1073 0.2705
R34572 VSS.n1073 VSS.n1071 0.2705
R34573 VSS.n1071 VSS.n1069 0.2705
R34574 VSS.n1069 VSS.n1067 0.2705
R34575 VSS.n1067 VSS.n1065 0.2705
R34576 VSS.n1065 VSS.n1063 0.2705
R34577 VSS.n1063 VSS.n1061 0.2705
R34578 VSS.n1061 VSS.n1059 0.2705
R34579 VSS.n1059 VSS.n1057 0.2705
R34580 VSS.n1057 VSS.n1055 0.2705
R34581 VSS.n1055 VSS.n1053 0.2705
R34582 VSS.n1053 VSS.n1051 0.2705
R34583 VSS.n1051 VSS.n1047 0.2705
R34584 VSS.n3370 VSS.n1047 0.2705
R34585 VSS.n3371 VSS.n3370 0.2705
R34586 VSS.n3340 VSS.n3339 0.2705
R34587 VSS.n3341 VSS.n3340 0.2705
R34588 VSS.n3342 VSS.n3341 0.2705
R34589 VSS.n3343 VSS.n3342 0.2705
R34590 VSS.n3344 VSS.n3343 0.2705
R34591 VSS.n3345 VSS.n3344 0.2705
R34592 VSS.n3346 VSS.n3345 0.2705
R34593 VSS.n3347 VSS.n3346 0.2705
R34594 VSS.n3348 VSS.n3347 0.2705
R34595 VSS.n3349 VSS.n3348 0.2705
R34596 VSS.n3350 VSS.n3349 0.2705
R34597 VSS.n3351 VSS.n3350 0.2705
R34598 VSS.n3352 VSS.n3351 0.2705
R34599 VSS.n3353 VSS.n3352 0.2705
R34600 VSS.n3354 VSS.n3353 0.2705
R34601 VSS.n3355 VSS.n3354 0.2705
R34602 VSS.n3356 VSS.n3355 0.2705
R34603 VSS.n3357 VSS.n3356 0.2705
R34604 VSS.n3358 VSS.n3357 0.2705
R34605 VSS.n3359 VSS.n3358 0.2705
R34606 VSS.n3360 VSS.n3359 0.2705
R34607 VSS.n3361 VSS.n3360 0.2705
R34608 VSS.n3362 VSS.n3361 0.2705
R34609 VSS.n3363 VSS.n3362 0.2705
R34610 VSS.n3364 VSS.n3363 0.2705
R34611 VSS.n3365 VSS.n3364 0.2705
R34612 VSS.n3366 VSS.n3365 0.2705
R34613 VSS.n3367 VSS.n3366 0.2705
R34614 VSS.n3368 VSS.n3367 0.2705
R34615 VSS.n3369 VSS.n3368 0.2705
R34616 VSS.n3369 VSS.n1045 0.2705
R34617 VSS.n1298 VSS.n1297 0.2705
R34618 VSS.n1299 VSS.n1298 0.2705
R34619 VSS.n1300 VSS.n1299 0.2705
R34620 VSS.n1301 VSS.n1300 0.2705
R34621 VSS.n1302 VSS.n1301 0.2705
R34622 VSS.n1303 VSS.n1302 0.2705
R34623 VSS.n1304 VSS.n1303 0.2705
R34624 VSS.n1305 VSS.n1304 0.2705
R34625 VSS.n1306 VSS.n1305 0.2705
R34626 VSS.n1307 VSS.n1306 0.2705
R34627 VSS.n1308 VSS.n1307 0.2705
R34628 VSS.n1309 VSS.n1308 0.2705
R34629 VSS.n1310 VSS.n1309 0.2705
R34630 VSS.n1311 VSS.n1310 0.2705
R34631 VSS.n1312 VSS.n1311 0.2705
R34632 VSS.n1313 VSS.n1312 0.2705
R34633 VSS.n1314 VSS.n1313 0.2705
R34634 VSS.n1315 VSS.n1314 0.2705
R34635 VSS.n1316 VSS.n1315 0.2705
R34636 VSS.n1317 VSS.n1316 0.2705
R34637 VSS.n1318 VSS.n1317 0.2705
R34638 VSS.n1319 VSS.n1318 0.2705
R34639 VSS.n1320 VSS.n1319 0.2705
R34640 VSS.n1321 VSS.n1320 0.2705
R34641 VSS.n1322 VSS.n1321 0.2705
R34642 VSS.n1323 VSS.n1322 0.2705
R34643 VSS.n1324 VSS.n1323 0.2705
R34644 VSS.n1325 VSS.n1324 0.2705
R34645 VSS.n1326 VSS.n1325 0.2705
R34646 VSS.n1327 VSS.n1326 0.2705
R34647 VSS.n1328 VSS.n1327 0.2705
R34648 VSS.n1329 VSS.n1328 0.2705
R34649 VSS.n1330 VSS.n1329 0.2705
R34650 VSS.n1331 VSS.n1330 0.2705
R34651 VSS.n1332 VSS.n1331 0.2705
R34652 VSS.n1333 VSS.n1332 0.2705
R34653 VSS.n1334 VSS.n1333 0.2705
R34654 VSS.n1256 VSS.n1255 0.2705
R34655 VSS.n1255 VSS.n1254 0.2705
R34656 VSS.n1254 VSS.n1253 0.2705
R34657 VSS.n1249 VSS.n1248 0.2705
R34658 VSS.n1250 VSS.n1249 0.2705
R34659 VSS.n1251 VSS.n1250 0.2705
R34660 VSS.n451 VSS.n450 0.2705
R34661 VSS.n454 VSS.n451 0.2705
R34662 VSS.n455 VSS.n454 0.2705
R34663 VSS.n1247 VSS.n1244 0.2705
R34664 VSS.n1245 VSS.n1244 0.2705
R34665 VSS.n1252 VSS.n1245 0.2705
R34666 VSS.n1257 VSS.n1241 0.2705
R34667 VSS.n1241 VSS.n1239 0.2705
R34668 VSS.n1239 VSS.n1237 0.2705
R34669 VSS.n1296 VSS.n1242 0.2705
R34670 VSS.n1242 VSS.n1240 0.2705
R34671 VSS.n1240 VSS.n1238 0.2705
R34672 VSS.n1238 VSS.n1236 0.2705
R34673 VSS.n1236 VSS.n1235 0.2705
R34674 VSS.n1235 VSS.n1234 0.2705
R34675 VSS.n1234 VSS.n1233 0.2705
R34676 VSS.n1233 VSS.n1232 0.2705
R34677 VSS.n1232 VSS.n1231 0.2705
R34678 VSS.n1231 VSS.n1230 0.2705
R34679 VSS.n1230 VSS.n1229 0.2705
R34680 VSS.n1229 VSS.n1228 0.2705
R34681 VSS.n1228 VSS.n1227 0.2705
R34682 VSS.n1227 VSS.n1226 0.2705
R34683 VSS.n1226 VSS.n1225 0.2705
R34684 VSS.n1225 VSS.n1224 0.2705
R34685 VSS.n1224 VSS.n1223 0.2705
R34686 VSS.n1223 VSS.n1222 0.2705
R34687 VSS.n1222 VSS.n1221 0.2705
R34688 VSS.n1221 VSS.n1220 0.2705
R34689 VSS.n1220 VSS.n1219 0.2705
R34690 VSS.n1219 VSS.n1218 0.2705
R34691 VSS.n1218 VSS.n1217 0.2705
R34692 VSS.n1217 VSS.n1216 0.2705
R34693 VSS.n1216 VSS.n1215 0.2705
R34694 VSS.n1215 VSS.n1214 0.2705
R34695 VSS.n1214 VSS.n1213 0.2705
R34696 VSS.n1213 VSS.n1212 0.2705
R34697 VSS.n1212 VSS.n1211 0.2705
R34698 VSS.n1211 VSS.n1210 0.2705
R34699 VSS.n1210 VSS.n1209 0.2705
R34700 VSS.n1209 VSS.n1208 0.2705
R34701 VSS.n1208 VSS.n1207 0.2705
R34702 VSS.n1207 VSS.n1206 0.2705
R34703 VSS.n1206 VSS.n1171 0.2705
R34704 VSS.n1171 VSS.n1169 0.2705
R34705 VSS.n1169 VSS.n1168 0.2705
R34706 VSS.n3588 VSS.n3587 0.2705
R34707 VSS.n3589 VSS.n3588 0.2705
R34708 VSS.n3590 VSS.n3589 0.2705
R34709 VSS.n3592 VSS.n3590 0.2705
R34710 VSS.n3594 VSS.n3592 0.2705
R34711 VSS.n3596 VSS.n3594 0.2705
R34712 VSS.n3598 VSS.n3596 0.2705
R34713 VSS.n3600 VSS.n3598 0.2705
R34714 VSS.n3602 VSS.n3600 0.2705
R34715 VSS.n3604 VSS.n3602 0.2705
R34716 VSS.n3606 VSS.n3604 0.2705
R34717 VSS.n3608 VSS.n3606 0.2705
R34718 VSS.n3610 VSS.n3608 0.2705
R34719 VSS.n3612 VSS.n3610 0.2705
R34720 VSS.n3614 VSS.n3612 0.2705
R34721 VSS.n3616 VSS.n3614 0.2705
R34722 VSS.n3618 VSS.n3616 0.2705
R34723 VSS.n3620 VSS.n3618 0.2705
R34724 VSS.n3621 VSS.n3620 0.2705
R34725 VSS.n3623 VSS.n3621 0.2705
R34726 VSS.n3665 VSS.n3664 0.2705
R34727 VSS.n3664 VSS.n3663 0.2705
R34728 VSS.n3663 VSS.n3662 0.2705
R34729 VSS.n3662 VSS.n3661 0.2705
R34730 VSS.n3661 VSS.n3660 0.2705
R34731 VSS.n3660 VSS.n3659 0.2705
R34732 VSS.n3659 VSS.n3658 0.2705
R34733 VSS.n3658 VSS.n3657 0.2705
R34734 VSS.n3657 VSS.n3656 0.2705
R34735 VSS.n3656 VSS.n3655 0.2705
R34736 VSS.n3655 VSS.n3654 0.2705
R34737 VSS.n3654 VSS.n3653 0.2705
R34738 VSS.n3653 VSS.n3652 0.2705
R34739 VSS.n3652 VSS.n3651 0.2705
R34740 VSS.n3651 VSS.n3650 0.2705
R34741 VSS.n3650 VSS.n3649 0.2705
R34742 VSS.n3649 VSS.n3648 0.2705
R34743 VSS.n3648 VSS.n3647 0.2705
R34744 VSS.n3647 VSS.n3646 0.2705
R34745 VSS.n3646 VSS.n3645 0.2705
R34746 VSS.n3585 VSS.n3584 0.2705
R34747 VSS.n3584 VSS.n3583 0.2705
R34748 VSS.n3583 VSS.n3582 0.2705
R34749 VSS.n3591 VSS.n3582 0.2705
R34750 VSS.n3593 VSS.n3591 0.2705
R34751 VSS.n3595 VSS.n3593 0.2705
R34752 VSS.n3597 VSS.n3595 0.2705
R34753 VSS.n3599 VSS.n3597 0.2705
R34754 VSS.n3601 VSS.n3599 0.2705
R34755 VSS.n3603 VSS.n3601 0.2705
R34756 VSS.n3605 VSS.n3603 0.2705
R34757 VSS.n3607 VSS.n3605 0.2705
R34758 VSS.n3609 VSS.n3607 0.2705
R34759 VSS.n3611 VSS.n3609 0.2705
R34760 VSS.n3613 VSS.n3611 0.2705
R34761 VSS.n3615 VSS.n3613 0.2705
R34762 VSS.n3617 VSS.n3615 0.2705
R34763 VSS.n3619 VSS.n3617 0.2705
R34764 VSS.n3622 VSS.n3619 0.2705
R34765 VSS.n3670 VSS.n3669 0.2705
R34766 VSS.n3671 VSS.n3670 0.2705
R34767 VSS.n3672 VSS.n3671 0.2705
R34768 VSS.n3580 VSS.n3579 0.2705
R34769 VSS.n3581 VSS.n3580 0.2705
R34770 VSS.n3673 VSS.n3581 0.2705
R34771 VSS.n3677 VSS.n3676 0.2705
R34772 VSS.n3676 VSS.n3675 0.2705
R34773 VSS.n3675 VSS.n3674 0.2705
R34774 VSS.n3577 VSS.n3575 0.2705
R34775 VSS.n3575 VSS.n3574 0.2705
R34776 VSS.n3574 VSS.n3573 0.2705
R34777 VSS.n3683 VSS.n3682 0.2705
R34778 VSS.n3684 VSS.n3683 0.2705
R34779 VSS.n3685 VSS.n3684 0.2705
R34780 VSS.n3576 VSS.n3571 0.2705
R34781 VSS.n3572 VSS.n3571 0.2705
R34782 VSS.n3686 VSS.n3572 0.2705
R34783 VSS.n3689 VSS.n3570 0.2705
R34784 VSS.n3689 VSS.n3688 0.2705
R34785 VSS.n3691 VSS.n3690 0.2705
R34786 VSS.n3690 VSS.n3563 0.2705
R34787 VSS.n3568 VSS.n3564 0.2705
R34788 VSS.n3791 VSS.n3564 0.2705
R34789 VSS.n3789 VSS.n3788 0.2705
R34790 VSS.n3790 VSS.n3789 0.2705
R34791 VSS.n3790 VSS.n3562 0.2705
R34792 VSS.n3567 VSS.n3566 0.2705
R34793 VSS.n3566 VSS.n3565 0.2705
R34794 VSS.n3779 VSS.n3565 0.2705
R34795 VSS.n3764 VSS.n3763 0.2705
R34796 VSS.n3765 VSS.n3764 0.2705
R34797 VSS.n3766 VSS.n3765 0.2705
R34798 VSS.n3767 VSS.n3766 0.2705
R34799 VSS.n3768 VSS.n3767 0.2705
R34800 VSS.n3769 VSS.n3768 0.2705
R34801 VSS.n3770 VSS.n3769 0.2705
R34802 VSS.n3771 VSS.n3770 0.2705
R34803 VSS.n3772 VSS.n3771 0.2705
R34804 VSS.n3773 VSS.n3772 0.2705
R34805 VSS.n3774 VSS.n3773 0.2705
R34806 VSS.n3775 VSS.n3774 0.2705
R34807 VSS.n3776 VSS.n3775 0.2705
R34808 VSS.n3784 VSS.n3776 0.2705
R34809 VSS.n3784 VSS.n3783 0.2705
R34810 VSS.n3783 VSS.n3782 0.2705
R34811 VSS.n3782 VSS.n3781 0.2705
R34812 VSS.n3721 VSS.n3719 0.2705
R34813 VSS.n3719 VSS.n3717 0.2705
R34814 VSS.n3717 VSS.n3715 0.2705
R34815 VSS.n3715 VSS.n3713 0.2705
R34816 VSS.n3713 VSS.n3711 0.2705
R34817 VSS.n3711 VSS.n3709 0.2705
R34818 VSS.n3709 VSS.n3707 0.2705
R34819 VSS.n3707 VSS.n3705 0.2705
R34820 VSS.n3705 VSS.n3703 0.2705
R34821 VSS.n3703 VSS.n3701 0.2705
R34822 VSS.n3701 VSS.n3699 0.2705
R34823 VSS.n3699 VSS.n3697 0.2705
R34824 VSS.n3697 VSS.n3696 0.2705
R34825 VSS.n3696 VSS.n3695 0.2705
R34826 VSS.n3777 VSS.n3695 0.2705
R34827 VSS.n3778 VSS.n3777 0.2705
R34828 VSS.n3759 VSS.n3758 0.2705
R34829 VSS.n3758 VSS.n3757 0.2705
R34830 VSS.n3757 VSS.n3756 0.2705
R34831 VSS.n3724 VSS.n3723 0.2705
R34832 VSS.n3725 VSS.n3724 0.2705
R34833 VSS.n3755 VSS.n3725 0.2705
R34834 VSS.n3734 VSS.n3733 0.2705
R34835 VSS.n3733 VSS.n3726 0.2705
R34836 VSS.n3754 VSS.n3726 0.2705
R34837 VSS.n3732 VSS.n3728 0.2705
R34838 VSS.n3752 VSS.n3728 0.2705
R34839 VSS.n3753 VSS.n3752 0.2705
R34840 VSS.n3750 VSS.n3749 0.2705
R34841 VSS.n3751 VSS.n3750 0.2705
R34842 VSS.n3751 VSS.n3727 0.2705
R34843 VSS.n3731 VSS.n3730 0.2705
R34844 VSS.n3730 VSS.n3729 0.2705
R34845 VSS.n3740 VSS.n3729 0.2705
R34846 VSS.n3745 VSS.n3744 0.2705
R34847 VSS.n3744 VSS.n3743 0.2705
R34848 VSS.n3739 VSS.n3738 0.2705
R34849 VSS.n3742 VSS.n3739 0.2705
R34850 VSS.n452 VSS.n449 0.2705
R34851 VSS.n453 VSS.n452 0.2705
R34852 VSS.n4186 VSS.n4185 0.2705
R34853 VSS.n4185 VSS.n4184 0.2705
R34854 VSS.n4184 VSS.n4183 0.2705
R34855 VSS.n1430 VSS.n1429 0.2705
R34856 VSS.n1431 VSS.n1430 0.2705
R34857 VSS.n3088 VSS.n1431 0.2705
R34858 VSS.n3092 VSS.n3091 0.2705
R34859 VSS.n3091 VSS.n3090 0.2705
R34860 VSS.n1427 VSS.n1426 0.2705
R34861 VSS.n1426 VSS.n1425 0.2705
R34862 VSS.n3097 VSS.n3096 0.2705
R34863 VSS.n3098 VSS.n3097 0.2705
R34864 VSS.n1422 VSS.n1421 0.2705
R34865 VSS.n1423 VSS.n1422 0.2705
R34866 VSS.n3100 VSS.n1423 0.2705
R34867 VSS.n3104 VSS.n3103 0.2705
R34868 VSS.n3103 VSS.n3102 0.2705
R34869 VSS.n3102 VSS.n3101 0.2705
R34870 VSS.n1419 VSS.n1418 0.2705
R34871 VSS.n1418 VSS.n1417 0.2705
R34872 VSS.n1417 VSS.n1416 0.2705
R34873 VSS.n3109 VSS.n3108 0.2705
R34874 VSS.n3110 VSS.n3109 0.2705
R34875 VSS.n3111 VSS.n3110 0.2705
R34876 VSS.n1414 VSS.n1413 0.2705
R34877 VSS.n1415 VSS.n1414 0.2705
R34878 VSS.n3112 VSS.n1415 0.2705
R34879 VSS.n3116 VSS.n3115 0.2705
R34880 VSS.n3115 VSS.n3114 0.2705
R34881 VSS.n3114 VSS.n3113 0.2705
R34882 VSS.n1411 VSS.n1410 0.2705
R34883 VSS.n1410 VSS.n1409 0.2705
R34884 VSS.n1409 VSS.n1408 0.2705
R34885 VSS.n3183 VSS.n3182 0.2705
R34886 VSS.n3184 VSS.n3183 0.2705
R34887 VSS.n3185 VSS.n3184 0.2705
R34888 VSS.n1378 VSS.n1377 0.2705
R34889 VSS.n1380 VSS.n1378 0.2705
R34890 VSS.n1382 VSS.n1380 0.2705
R34891 VSS.n1384 VSS.n1382 0.2705
R34892 VSS.n1386 VSS.n1384 0.2705
R34893 VSS.n1388 VSS.n1386 0.2705
R34894 VSS.n1390 VSS.n1388 0.2705
R34895 VSS.n1392 VSS.n1390 0.2705
R34896 VSS.n1394 VSS.n1392 0.2705
R34897 VSS.n1396 VSS.n1394 0.2705
R34898 VSS.n1398 VSS.n1396 0.2705
R34899 VSS.n1400 VSS.n1398 0.2705
R34900 VSS.n1402 VSS.n1400 0.2705
R34901 VSS.n1404 VSS.n1402 0.2705
R34902 VSS.n1406 VSS.n1404 0.2705
R34903 VSS.n1407 VSS.n1406 0.2705
R34904 VSS.n3186 VSS.n1407 0.2705
R34905 VSS.n3204 VSS.n3203 0.2705
R34906 VSS.n3203 VSS.n3202 0.2705
R34907 VSS.n3202 VSS.n3201 0.2705
R34908 VSS.n3201 VSS.n3200 0.2705
R34909 VSS.n3200 VSS.n3199 0.2705
R34910 VSS.n3199 VSS.n3198 0.2705
R34911 VSS.n3198 VSS.n3197 0.2705
R34912 VSS.n3197 VSS.n3196 0.2705
R34913 VSS.n3196 VSS.n3195 0.2705
R34914 VSS.n3195 VSS.n3194 0.2705
R34915 VSS.n3194 VSS.n3193 0.2705
R34916 VSS.n3193 VSS.n3192 0.2705
R34917 VSS.n3192 VSS.n3191 0.2705
R34918 VSS.n3191 VSS.n3190 0.2705
R34919 VSS.n3190 VSS.n3189 0.2705
R34920 VSS.n3189 VSS.n3188 0.2705
R34921 VSS.n3530 VSS.n3529 0.26825
R34922 VSS.n3991 VSS.n3990 0.261026
R34923 VSS.n3801 VSS.n3800 0.2605
R34924 VSS.n3801 VSS.n707 0.2605
R34925 VSS.n3864 VSS.n3554 0.252366
R34926 VSS.n3519 VSS.n3518 0.2485
R34927 VSS.n3213 VSS.n1371 0.2485
R34928 VSS.n4131 VSS.n4130 0.248
R34929 VSS.n3535 VSS.n3534 0.248
R34930 VSS.n744 VSS.n743 0.248
R34931 VSS.n1783 VSS.n1782 0.248
R34932 VSS.n2176 VSS.n2175 0.248
R34933 VSS.n1830 VSS.n1829 0.248
R34934 VSS.n1361 VSS.n1360 0.248
R34935 VSS.n3318 VSS.n3317 0.248
R34936 VSS.n3169 VSS.n3168 0.248
R34937 VSS.n3182 VSS.n3181 0.248
R34938 VSS.n3785 VSS.n3567 0.248
R34939 VSS.n1357 VSS.n1356 0.247929
R34940 VSS.n740 VSS.n739 0.246929
R34941 VSS.n3859 VSS.n3553 0.244855
R34942 VSS.n1919 VSS.n1918 0.242079
R34943 VSS.n1391 VSS.n1375 0.242
R34944 VSS.n3861 VSS.n3860 0.24169
R34945 VSS.n1799 VSS.n1798 0.240895
R34946 VSS.n4181 VSS.n4180 0.238278
R34947 VSS.n1013 VSS.n777 0.237342
R34948 VSS.n3512 VSS.n770 0.237342
R34949 VSS.n890 VSS.n735 0.23675
R34950 VSS.n3428 VSS.n3427 0.23675
R34951 VSS.n3426 VSS.n889 0.23675
R34952 VSS.n933 VSS.n891 0.23675
R34953 VSS.n935 VSS.n934 0.23675
R34954 VSS.n937 VSS.n936 0.23675
R34955 VSS.n929 VSS.n928 0.23675
R34956 VSS.n942 VSS.n941 0.23675
R34957 VSS.n943 VSS.n927 0.23675
R34958 VSS.n946 VSS.n945 0.23675
R34959 VSS.n947 VSS.n898 0.23675
R34960 VSS.n3419 VSS.n899 0.23675
R34961 VSS.n3532 VSS.n736 0.23675
R34962 VSS.n3389 VSS.n3388 0.235126
R34963 VSS.n3385 VSS.n3384 0.235126
R34964 VSS.n2182 VSS.n2181 0.22775
R34965 VSS.n2180 VSS.n1658 0.22775
R34966 VSS.n1798 VSS.n1662 0.22775
R34967 VSS.n1802 VSS.n1797 0.22775
R34968 VSS.n1801 VSS.n1800 0.22775
R34969 VSS.n4097 VSS.n510 0.226
R34970 VSS.n3952 VSS.n3880 0.226
R34971 VSS.n4021 VSS.n4020 0.226
R34972 VSS.n3516 VSS.n768 0.226
R34973 VSS.n2228 VSS.n1636 0.226
R34974 VSS.n1990 VSS.n1989 0.226
R34975 VSS.n3482 VSS.n810 0.226
R34976 VSS.n1968 VSS.n1855 0.226
R34977 VSS.n2213 VSS.n1646 0.226
R34978 VSS.n3447 VSS.n872 0.226
R34979 VSS.n4041 VSS.n4040 0.226
R34980 VSS.n4081 VSS.n4080 0.226
R34981 VSS.n3932 VSS.n3915 0.226
R34982 VSS.n3209 VSS.n3208 0.226
R34983 VSS.n2244 VSS.n1617 0.226
R34984 VSS.n2263 VSS.n2262 0.226
R34985 VSS.n3078 VSS.n3077 0.226
R34986 VSS.n3372 VSS.n1044 0.226
R34987 VSS.n3337 VSS.n1106 0.226
R34988 VSS.n1335 VSS.n1167 0.226
R34989 VSS.n3762 VSS.n3761 0.226
R34990 VSS.n3666 VSS.n3586 0.226
R34991 VSS.n4082 VSS.n525 0.2255
R34992 VSS.n4083 VSS.n524 0.2255
R34993 VSS.n4084 VSS.n523 0.2255
R34994 VSS.n4085 VSS.n522 0.2255
R34995 VSS.n4086 VSS.n521 0.2255
R34996 VSS.n4087 VSS.n520 0.2255
R34997 VSS.n4088 VSS.n519 0.2255
R34998 VSS.n4089 VSS.n518 0.2255
R34999 VSS.n4090 VSS.n517 0.2255
R35000 VSS.n4091 VSS.n516 0.2255
R35001 VSS.n4092 VSS.n515 0.2255
R35002 VSS.n4093 VSS.n514 0.2255
R35003 VSS.n4094 VSS.n513 0.2255
R35004 VSS.n4096 VSS.n511 0.2255
R35005 VSS.n4095 VSS.n512 0.2255
R35006 VSS.n3977 VSS.n3914 0.2255
R35007 VSS.n3978 VSS.n3913 0.2255
R35008 VSS.n3985 VSS.n3984 0.2255
R35009 VSS.n3983 VSS.n3912 0.2255
R35010 VSS.n3982 VSS.n3981 0.2255
R35011 VSS.n482 VSS.n481 0.2255
R35012 VSS.n4137 VSS.n4136 0.2255
R35013 VSS.n4135 VSS.n480 0.2255
R35014 VSS.n4134 VSS.n483 0.2255
R35015 VSS.n4133 VSS.n484 0.2255
R35016 VSS.n4098 VSS.n4097 0.2255
R35017 VSS.n4010 VSS.n3879 0.2255
R35018 VSS.n4013 VSS.n4012 0.2255
R35019 VSS.n4011 VSS.n3877 0.2255
R35020 VSS.n4017 VSS.n3876 0.2255
R35021 VSS.n4019 VSS.n4018 0.2255
R35022 VSS.n4020 VSS.n712 0.2255
R35023 VSS.n3442 VSS.n877 0.2255
R35024 VSS.n732 VSS.n729 0.2255
R35025 VSS.n3431 VSS.n3430 0.2255
R35026 VSS.n3432 VSS.n887 0.2255
R35027 VSS.n3433 VSS.n886 0.2255
R35028 VSS.n3434 VSS.n885 0.2255
R35029 VSS.n3435 VSS.n884 0.2255
R35030 VSS.n3436 VSS.n883 0.2255
R35031 VSS.n3437 VSS.n882 0.2255
R35032 VSS.n3438 VSS.n881 0.2255
R35033 VSS.n3439 VSS.n880 0.2255
R35034 VSS.n3440 VSS.n879 0.2255
R35035 VSS.n3441 VSS.n878 0.2255
R35036 VSS.n737 VSS.n718 0.2255
R35037 VSS.n3514 VSS.n768 0.2255
R35038 VSS.n2159 VSS.n1854 0.2255
R35039 VSS.n2160 VSS.n1853 0.2255
R35040 VSS.n2161 VSS.n1852 0.2255
R35041 VSS.n2162 VSS.n1851 0.2255
R35042 VSS.n2163 VSS.n1850 0.2255
R35043 VSS.n2164 VSS.n1849 0.2255
R35044 VSS.n2165 VSS.n1848 0.2255
R35045 VSS.n2166 VSS.n1847 0.2255
R35046 VSS.n2167 VSS.n1846 0.2255
R35047 VSS.n2168 VSS.n1845 0.2255
R35048 VSS.n2169 VSS.n1844 0.2255
R35049 VSS.n2170 VSS.n1843 0.2255
R35050 VSS.n2171 VSS.n1842 0.2255
R35051 VSS.n2172 VSS.n1841 0.2255
R35052 VSS.n2173 VSS.n1667 0.2255
R35053 VSS.n1856 VSS.n1855 0.2255
R35054 VSS.n1990 VSS.n1949 0.2255
R35055 VSS.n2158 VSS.n2157 0.2255
R35056 VSS.n2138 VSS.n1991 0.2255
R35057 VSS.n2137 VSS.n2136 0.2255
R35058 VSS.n2135 VSS.n1992 0.2255
R35059 VSS.n2134 VSS.n2133 0.2255
R35060 VSS.n1994 VSS.n1993 0.2255
R35061 VSS.n2016 VSS.n2015 0.2255
R35062 VSS.n2018 VSS.n2017 0.2255
R35063 VSS.n2025 VSS.n2014 0.2255
R35064 VSS.n2027 VSS.n2026 0.2255
R35065 VSS.n2028 VSS.n2012 0.2255
R35066 VSS.n2119 VSS.n2029 0.2255
R35067 VSS.n2118 VSS.n2117 0.2255
R35068 VSS.n2116 VSS.n2030 0.2255
R35069 VSS.n2115 VSS.n2114 0.2255
R35070 VSS.n2032 VSS.n2031 0.2255
R35071 VSS.n2046 VSS.n2045 0.2255
R35072 VSS.n2048 VSS.n2047 0.2255
R35073 VSS.n2049 VSS.n2043 0.2255
R35074 VSS.n2092 VSS.n2050 0.2255
R35075 VSS.n2091 VSS.n2090 0.2255
R35076 VSS.n2089 VSS.n2051 0.2255
R35077 VSS.n2088 VSS.n2087 0.2255
R35078 VSS.n2053 VSS.n2052 0.2255
R35079 VSS.n2062 VSS.n2061 0.2255
R35080 VSS.n2072 VSS.n2063 0.2255
R35081 VSS.n2071 VSS.n2070 0.2255
R35082 VSS.n2069 VSS.n2067 0.2255
R35083 VSS.n2068 VSS.n1635 0.2255
R35084 VSS.n2211 VSS.n1646 0.2255
R35085 VSS.n2230 VSS.n1636 0.2255
R35086 VSS.n1828 VSS.n1678 0.2255
R35087 VSS.n1718 VSS.n1682 0.2255
R35088 VSS.n1720 VSS.n1719 0.2255
R35089 VSS.n1721 VSS.n1717 0.2255
R35090 VSS.n1730 VSS.n1729 0.2255
R35091 VSS.n1731 VSS.n1716 0.2255
R35092 VSS.n1733 VSS.n1732 0.2255
R35093 VSS.n1710 VSS.n1709 0.2255
R35094 VSS.n1743 VSS.n1742 0.2255
R35095 VSS.n1744 VSS.n1707 0.2255
R35096 VSS.n1748 VSS.n1747 0.2255
R35097 VSS.n1746 VSS.n1708 0.2255
R35098 VSS.n3443 VSS.n876 0.2255
R35099 VSS.n1745 VSS.n806 0.2255
R35100 VSS.n3444 VSS.n875 0.2255
R35101 VSS.n3486 VSS.n808 0.2255
R35102 VSS.n3445 VSS.n874 0.2255
R35103 VSS.n3485 VSS.n3484 0.2255
R35104 VSS.n3446 VSS.n873 0.2255
R35105 VSS.n3483 VSS.n809 0.2255
R35106 VSS.n3448 VSS.n3447 0.2255
R35107 VSS.n3482 VSS.n3481 0.2255
R35108 VSS.n3870 VSS.n3549 0.2255
R35109 VSS.n3869 VSS.n3868 0.2255
R35110 VSS.n3867 VSS.n3550 0.2255
R35111 VSS.n3866 VSS.n3865 0.2255
R35112 VSS.n3552 VSS.n3551 0.2255
R35113 VSS.n3812 VSS.n3811 0.2255
R35114 VSS.n3814 VSS.n3813 0.2255
R35115 VSS.n3815 VSS.n3809 0.2255
R35116 VSS.n3846 VSS.n3816 0.2255
R35117 VSS.n3845 VSS.n3844 0.2255
R35118 VSS.n3843 VSS.n3817 0.2255
R35119 VSS.n3842 VSS.n3841 0.2255
R35120 VSS.n3819 VSS.n3818 0.2255
R35121 VSS.n3823 VSS.n3822 0.2255
R35122 VSS.n3825 VSS.n3824 0.2255
R35123 VSS.n601 VSS.n600 0.2255
R35124 VSS.n4039 VSS.n4038 0.2255
R35125 VSS.n4081 VSS.n526 0.2255
R35126 VSS.n4040 VSS.n599 0.2255
R35127 VSS.n3916 VSS.n3915 0.2255
R35128 VSS.n3881 VSS.n3880 0.2255
R35129 VSS.n3976 VSS.n3975 0.2255
R35130 VSS.n4009 VSS.n4008 0.2255
R35131 VSS.n1336 VSS.n1166 0.2255
R35132 VSS.n1337 VSS.n1165 0.2255
R35133 VSS.n1338 VSS.n1164 0.2255
R35134 VSS.n1339 VSS.n1163 0.2255
R35135 VSS.n1340 VSS.n1162 0.2255
R35136 VSS.n1341 VSS.n1161 0.2255
R35137 VSS.n1342 VSS.n1160 0.2255
R35138 VSS.n1343 VSS.n1159 0.2255
R35139 VSS.n1344 VSS.n1158 0.2255
R35140 VSS.n1345 VSS.n1157 0.2255
R35141 VSS.n1346 VSS.n1156 0.2255
R35142 VSS.n1347 VSS.n1155 0.2255
R35143 VSS.n1348 VSS.n1154 0.2255
R35144 VSS.n1349 VSS.n1153 0.2255
R35145 VSS.n1350 VSS.n1152 0.2255
R35146 VSS.n1351 VSS.n1151 0.2255
R35147 VSS.n1352 VSS.n1150 0.2255
R35148 VSS.n3210 VSS.n3209 0.2255
R35149 VSS.n1355 VSS.n1138 0.2255
R35150 VSS.n3320 VSS.n1123 0.2255
R35151 VSS.n3321 VSS.n1122 0.2255
R35152 VSS.n3322 VSS.n1121 0.2255
R35153 VSS.n3323 VSS.n1120 0.2255
R35154 VSS.n3324 VSS.n1119 0.2255
R35155 VSS.n3325 VSS.n1118 0.2255
R35156 VSS.n3326 VSS.n1117 0.2255
R35157 VSS.n3327 VSS.n1116 0.2255
R35158 VSS.n3328 VSS.n1115 0.2255
R35159 VSS.n3329 VSS.n1114 0.2255
R35160 VSS.n3330 VSS.n1113 0.2255
R35161 VSS.n3331 VSS.n1112 0.2255
R35162 VSS.n3332 VSS.n1111 0.2255
R35163 VSS.n3333 VSS.n1110 0.2255
R35164 VSS.n3400 VSS.n1015 0.2255
R35165 VSS.n3400 VSS.n3399 0.2255
R35166 VSS.n1440 VSS.n1439 0.2255
R35167 VSS.n3083 VSS.n3082 0.2255
R35168 VSS.n3081 VSS.n1438 0.2255
R35169 VSS.n3080 VSS.n1441 0.2255
R35170 VSS.n2245 VSS.n2244 0.2255
R35171 VSS.n2263 VSS.n1507 0.2255
R35172 VSS.n2264 VSS.n1506 0.2255
R35173 VSS.n2265 VSS.n1505 0.2255
R35174 VSS.n2266 VSS.n1504 0.2255
R35175 VSS.n2267 VSS.n1503 0.2255
R35176 VSS.n2268 VSS.n1502 0.2255
R35177 VSS.n2269 VSS.n1501 0.2255
R35178 VSS.n2270 VSS.n1500 0.2255
R35179 VSS.n2271 VSS.n1499 0.2255
R35180 VSS.n2272 VSS.n1498 0.2255
R35181 VSS.n2273 VSS.n1497 0.2255
R35182 VSS.n2274 VSS.n1496 0.2255
R35183 VSS.n2275 VSS.n1495 0.2255
R35184 VSS.n2276 VSS.n1494 0.2255
R35185 VSS.n2277 VSS.n1493 0.2255
R35186 VSS.n2278 VSS.n1492 0.2255
R35187 VSS.n2279 VSS.n1491 0.2255
R35188 VSS.n2280 VSS.n1490 0.2255
R35189 VSS.n2281 VSS.n1489 0.2255
R35190 VSS.n2282 VSS.n1488 0.2255
R35191 VSS.n2283 VSS.n1487 0.2255
R35192 VSS.n2284 VSS.n1486 0.2255
R35193 VSS.n2285 VSS.n1485 0.2255
R35194 VSS.n2286 VSS.n1484 0.2255
R35195 VSS.n3055 VSS.n1481 0.2255
R35196 VSS.n3079 VSS.n1442 0.2255
R35197 VSS.n3078 VSS.n1443 0.2255
R35198 VSS.n3167 VSS.n3119 0.2255
R35199 VSS.n3128 VSS.n3121 0.2255
R35200 VSS.n3129 VSS.n3127 0.2255
R35201 VSS.n3160 VSS.n3130 0.2255
R35202 VSS.n3159 VSS.n3158 0.2255
R35203 VSS.n3157 VSS.n3131 0.2255
R35204 VSS.n3156 VSS.n3155 0.2255
R35205 VSS.n3133 VSS.n3132 0.2255
R35206 VSS.n3141 VSS.n3140 0.2255
R35207 VSS.n3148 VSS.n3142 0.2255
R35208 VSS.n3147 VSS.n3146 0.2255
R35209 VSS.n3145 VSS.n3143 0.2255
R35210 VSS.n3144 VSS.n1040 0.2255
R35211 VSS.n3334 VSS.n1109 0.2255
R35212 VSS.n3376 VSS.n1042 0.2255
R35213 VSS.n3335 VSS.n1108 0.2255
R35214 VSS.n3375 VSS.n3374 0.2255
R35215 VSS.n3336 VSS.n1107 0.2255
R35216 VSS.n3373 VSS.n1043 0.2255
R35217 VSS.n3338 VSS.n3337 0.2255
R35218 VSS.n3372 VSS.n3371 0.2255
R35219 VSS.n1335 VSS.n1334 0.2255
R35220 VSS.n3666 VSS.n3665 0.2255
R35221 VSS.n3667 VSS.n3585 0.2255
R35222 VSS.n3669 VSS.n3668 0.2255
R35223 VSS.n3579 VSS.n3578 0.2255
R35224 VSS.n3678 VSS.n3677 0.2255
R35225 VSS.n3679 VSS.n3577 0.2255
R35226 VSS.n3682 VSS.n3681 0.2255
R35227 VSS.n3680 VSS.n3576 0.2255
R35228 VSS.n3570 VSS.n3569 0.2255
R35229 VSS.n3688 VSS.n3687 0.2255
R35230 VSS.n3692 VSS.n3691 0.2255
R35231 VSS.n3563 VSS.n3561 0.2255
R35232 VSS.n3693 VSS.n3568 0.2255
R35233 VSS.n3792 VSS.n3791 0.2255
R35234 VSS.n3788 VSS.n3787 0.2255
R35235 VSS.n3761 VSS.n3721 0.2255
R35236 VSS.n3760 VSS.n3759 0.2255
R35237 VSS.n3723 VSS.n3722 0.2255
R35238 VSS.n3735 VSS.n3734 0.2255
R35239 VSS.n3736 VSS.n3732 0.2255
R35240 VSS.n3749 VSS.n3748 0.2255
R35241 VSS.n3747 VSS.n3731 0.2255
R35242 VSS.n3746 VSS.n3745 0.2255
R35243 VSS.n3743 VSS.n3741 0.2255
R35244 VSS.n3738 VSS.n3737 0.2255
R35245 VSS.n3742 VSS.n456 0.2255
R35246 VSS.n449 VSS.n448 0.2255
R35247 VSS.n4182 VSS.n453 0.2255
R35248 VSS.n4187 VSS.n4186 0.2255
R35249 VSS.n1429 VSS.n1428 0.2255
R35250 VSS.n3093 VSS.n3092 0.2255
R35251 VSS.n3090 VSS.n3089 0.2255
R35252 VSS.n3094 VSS.n1427 0.2255
R35253 VSS.n1432 VSS.n1425 0.2255
R35254 VSS.n3096 VSS.n3095 0.2255
R35255 VSS.n3099 VSS.n3098 0.2255
R35256 VSS.n1421 VSS.n1420 0.2255
R35257 VSS.n3105 VSS.n3104 0.2255
R35258 VSS.n3106 VSS.n1419 0.2255
R35259 VSS.n3108 VSS.n3107 0.2255
R35260 VSS.n1413 VSS.n1412 0.2255
R35261 VSS.n3117 VSS.n3116 0.2255
R35262 VSS.n3118 VSS.n1411 0.2255
R35263 VSS.n2193 VSS.n2192 0.219609
R35264 VSS.n642 VSS.n641 0.218395
R35265 VSS.n1181 VSS.n1180 0.210118
R35266 VSS.n3933 VSS.n3932 0.208
R35267 VSS.n3518 VSS.n3517 0.208
R35268 VSS.n3517 VSS.n3516 0.208
R35269 VSS.n1968 VSS.n1967 0.208
R35270 VSS.n1989 VSS.n1950 0.208
R35271 VSS.n2228 VSS.n2227 0.208
R35272 VSS.n2214 VSS.n2213 0.208
R35273 VSS.n814 VSS.n810 0.208
R35274 VSS.n872 VSS.n870 0.208
R35275 VSS.n4041 VSS.n598 0.208
R35276 VSS.n4080 VSS.n527 0.208
R35277 VSS.n510 VSS.n508 0.208
R35278 VSS.n3952 VSS.n3951 0.208
R35279 VSS.n3624 VSS.n3586 0.208
R35280 VSS.n3762 VSS.n3720 0.208
R35281 VSS.n3208 VSS.n3207 0.208
R35282 VSS.n3207 VSS.n1371 0.208
R35283 VSS.n3077 VSS.n1444 0.208
R35284 VSS.n1048 VSS.n1044 0.208
R35285 VSS.n1106 VSS.n1104 0.208
R35286 VSS.n1259 VSS.n1167 0.208
R35287 VSS.n3643 VSS.n3642 0.208
R35288 VSS.n1617 VSS.n1616 0.208
R35289 VSS.n2262 VSS.n1508 0.208
R35290 VSS.n677 VSS.n676 0.206553
R35291 VSS.n1796 VSS.n1789 0.20525
R35292 VSS.n3100 VSS.n3099 0.195376
R35293 VSS.n3089 VSS.n3088 0.195376
R35294 VSS.n2240 VSS.n1424 0.194912
R35295 VSS.n1689 VSS.n1687 0.194711
R35296 VSS.n3792 VSS.n3562 0.192914
R35297 VSS.n3687 VSS.n3686 0.192914
R35298 VSS.n3741 VSS.n3740 0.192038
R35299 VSS.n4183 VSS.n4182 0.192038
R35300 VSS.n3830 VSS.n3829 0.189974
R35301 VSS.n3837 VSS.n3836 0.189974
R35302 VSS.n3836 VSS.n3835 0.189974
R35303 VSS.n3835 VSS.n3832 0.189974
R35304 VSS.n3832 VSS.n3805 0.189974
R35305 VSS.n3850 VSS.n3805 0.189974
R35306 VSS.n3804 VSS.n3557 0.189974
R35307 VSS.n3861 VSS.n3557 0.189974
R35308 VSS.n4033 VSS.n4032 0.189974
R35309 VSS.n4032 VSS.n4031 0.189974
R35310 VSS.n689 VSS.n605 0.189974
R35311 VSS.n690 VSS.n689 0.189974
R35312 VSS.n691 VSS.n690 0.189974
R35313 VSS.n692 VSS.n691 0.189974
R35314 VSS.n693 VSS.n692 0.189974
R35315 VSS.n694 VSS.n693 0.189974
R35316 VSS.n695 VSS.n694 0.189974
R35317 VSS.n696 VSS.n695 0.189974
R35318 VSS.n697 VSS.n696 0.189974
R35319 VSS.n698 VSS.n697 0.189974
R35320 VSS.n699 VSS.n698 0.189974
R35321 VSS.n700 VSS.n699 0.189974
R35322 VSS.n701 VSS.n700 0.189974
R35323 VSS.n702 VSS.n701 0.189974
R35324 VSS.n688 VSS.n687 0.189974
R35325 VSS.n687 VSS.n686 0.189974
R35326 VSS.n686 VSS.n685 0.189974
R35327 VSS.n685 VSS.n684 0.189974
R35328 VSS.n684 VSS.n683 0.189974
R35329 VSS.n683 VSS.n682 0.189974
R35330 VSS.n682 VSS.n681 0.189974
R35331 VSS.n681 VSS.n680 0.189974
R35332 VSS.n680 VSS.n679 0.189974
R35333 VSS.n679 VSS.n678 0.189974
R35334 VSS.n678 VSS.n677 0.189974
R35335 VSS.n674 VSS.n608 0.189974
R35336 VSS.n659 VSS.n618 0.189974
R35337 VSS.n658 VSS.n657 0.189974
R35338 VSS.n659 VSS.n658 0.189974
R35339 VSS.n656 VSS.n620 0.189974
R35340 VSS.n657 VSS.n656 0.189974
R35341 VSS.n644 VSS.n628 0.189974
R35342 VSS.n643 VSS.n642 0.189974
R35343 VSS.n644 VSS.n643 0.189974
R35344 VSS.n641 VSS.n640 0.189974
R35345 VSS.n640 VSS.n639 0.189974
R35346 VSS.n639 VSS.n638 0.189974
R35347 VSS.n638 VSS.n637 0.189974
R35348 VSS.n637 VSS.n636 0.189974
R35349 VSS.n636 VSS.n635 0.189974
R35350 VSS.n635 VSS.n460 0.189974
R35351 VSS.n4156 VSS.n4155 0.189974
R35352 VSS.n4155 VSS.n4154 0.189974
R35353 VSS.n4154 VSS.n4153 0.189974
R35354 VSS.n4152 VSS.n465 0.189974
R35355 VSS.n4153 VSS.n4152 0.189974
R35356 VSS.n3998 VSS.n3996 0.189974
R35357 VSS.n3996 VSS.n3995 0.189974
R35358 VSS.n3995 VSS.n3994 0.189974
R35359 VSS.n3994 VSS.n3993 0.189974
R35360 VSS.n3993 VSS.n3992 0.189974
R35361 VSS.n3992 VSS.n3991 0.189974
R35362 VSS.n3990 VSS.n3904 0.189974
R35363 VSS.n3907 VSS.n3904 0.189974
R35364 VSS.n3907 VSS.n472 0.189974
R35365 VSS.n4142 VSS.n473 0.189974
R35366 VSS.n4119 VSS.n473 0.189974
R35367 VSS.n4123 VSS.n4119 0.189974
R35368 VSS.n4124 VSS.n4123 0.189974
R35369 VSS.n4126 VSS.n4124 0.189974
R35370 VSS.n4149 VSS.n468 0.189974
R35371 VSS.n3857 VSS.n3856 0.189974
R35372 VSS.n3896 VSS.n3894 0.189974
R35373 VSS.n3894 VSS.n3892 0.189974
R35374 VSS.n3892 VSS.n3890 0.189974
R35375 VSS.n3890 VSS.n3888 0.189974
R35376 VSS.n3888 VSS.n3886 0.189974
R35377 VSS.n3886 VSS.n3884 0.189974
R35378 VSS.n3884 VSS.n3878 0.189974
R35379 VSS.n4015 VSS.n4014 0.189974
R35380 VSS.n4016 VSS.n4015 0.189974
R35381 VSS.n4016 VSS.n711 0.189974
R35382 VSS.n4024 VSS.n4023 0.189974
R35383 VSS.n4023 VSS.n3875 0.189974
R35384 VSS.n1739 VSS.n1704 0.189974
R35385 VSS.n1737 VSS.n1736 0.189974
R35386 VSS.n1736 VSS.n1713 0.189974
R35387 VSS.n1726 VSS.n1713 0.189974
R35388 VSS.n1726 VSS.n1725 0.189974
R35389 VSS.n1725 VSS.n1724 0.189974
R35390 VSS.n1824 VSS.n1823 0.189974
R35391 VSS.n1823 VSS.n1822 0.189974
R35392 VSS.n1822 VSS.n1687 0.189974
R35393 VSS.n1760 VSS.n769 0.189974
R35394 VSS.n801 VSS.n799 0.189974
R35395 VSS.n799 VSS.n797 0.189974
R35396 VSS.n797 VSS.n795 0.189974
R35397 VSS.n795 VSS.n793 0.189974
R35398 VSS.n793 VSS.n791 0.189974
R35399 VSS.n791 VSS.n789 0.189974
R35400 VSS.n789 VSS.n787 0.189974
R35401 VSS.n787 VSS.n785 0.189974
R35402 VSS.n783 VSS.n778 0.189974
R35403 VSS.n3503 VSS.n778 0.189974
R35404 VSS.n3427 VSS.n890 0.189974
R35405 VSS.n3427 VSS.n3426 0.189974
R35406 VSS.n935 VSS.n891 0.189974
R35407 VSS.n936 VSS.n935 0.189974
R35408 VSS.n936 VSS.n928 0.189974
R35409 VSS.n942 VSS.n928 0.189974
R35410 VSS.n943 VSS.n942 0.189974
R35411 VSS.n945 VSS.n898 0.189974
R35412 VSS.n3418 VSS.n3417 0.189974
R35413 VSS.n3417 VSS.n3416 0.189974
R35414 VSS.n3416 VSS.n3415 0.189974
R35415 VSS.n3413 VSS.n3412 0.189974
R35416 VSS.n3412 VSS.n3411 0.189974
R35417 VSS.n3411 VSS.n3410 0.189974
R35418 VSS.n3410 VSS.n3409 0.189974
R35419 VSS.n3409 VSS.n3408 0.189974
R35420 VSS.n1014 VSS.n1013 0.189974
R35421 VSS.n770 VSS.n764 0.189974
R35422 VSS.n763 VSS.n762 0.189974
R35423 VSS.n762 VSS.n761 0.189974
R35424 VSS.n761 VSS.n760 0.189974
R35425 VSS.n760 VSS.n759 0.189974
R35426 VSS.n759 VSS.n758 0.189974
R35427 VSS.n757 VSS.n756 0.189974
R35428 VSS.n756 VSS.n755 0.189974
R35429 VSS.n755 VSS.n754 0.189974
R35430 VSS.n890 VSS.n736 0.189974
R35431 VSS.n1690 VSS.n1689 0.189974
R35432 VSS.n1691 VSS.n1690 0.189974
R35433 VSS.n1692 VSS.n1691 0.189974
R35434 VSS.n1693 VSS.n1692 0.189974
R35435 VSS.n1694 VSS.n1693 0.189974
R35436 VSS.n1695 VSS.n1694 0.189974
R35437 VSS.n1696 VSS.n1695 0.189974
R35438 VSS.n1697 VSS.n1696 0.189974
R35439 VSS.n1761 VSS.n1760 0.189974
R35440 VSS.n2064 VSS.n2058 0.189974
R35441 VSS.n2075 VSS.n2058 0.189974
R35442 VSS.n2076 VSS.n2075 0.189974
R35443 VSS.n2083 VSS.n2082 0.189974
R35444 VSS.n2082 VSS.n2081 0.189974
R35445 VSS.n2081 VSS.n2078 0.189974
R35446 VSS.n2078 VSS.n2038 0.189974
R35447 VSS.n2096 VSS.n2038 0.189974
R35448 VSS.n2096 VSS.n2039 0.189974
R35449 VSS.n2039 VSS.n2037 0.189974
R35450 VSS.n2105 VSS.n2104 0.189974
R35451 VSS.n2104 VSS.n2101 0.189974
R35452 VSS.n2101 VSS.n2007 0.189974
R35453 VSS.n2123 VSS.n2008 0.189974
R35454 VSS.n2022 VSS.n2008 0.189974
R35455 VSS.n2022 VSS.n2021 0.189974
R35456 VSS.n2021 VSS.n1999 0.189974
R35457 VSS.n2129 VSS.n1999 0.189974
R35458 VSS.n2002 VSS.n2000 0.189974
R35459 VSS.n1944 VSS.n1942 0.189974
R35460 VSS.n1942 VSS.n1940 0.189974
R35461 VSS.n1937 VSS.n1935 0.189974
R35462 VSS.n1935 VSS.n1933 0.189974
R35463 VSS.n1933 VSS.n1931 0.189974
R35464 VSS.n1931 VSS.n1929 0.189974
R35465 VSS.n1929 VSS.n1927 0.189974
R35466 VSS.n1923 VSS.n1921 0.189974
R35467 VSS.n1921 VSS.n1919 0.189974
R35468 VSS.n1916 VSS.n1915 0.189974
R35469 VSS.n1911 VSS.n1910 0.189974
R35470 VSS.n1912 VSS.n1911 0.189974
R35471 VSS.n1909 VSS.n1872 0.189974
R35472 VSS.n1910 VSS.n1909 0.189974
R35473 VSS.n1879 VSS.n1872 0.189974
R35474 VSS.n1890 VSS.n1889 0.189974
R35475 VSS.n1891 VSS.n1890 0.189974
R35476 VSS.n1630 VSS.n1625 0.189974
R35477 VSS.n2236 VSS.n1625 0.189974
R35478 VSS.n2202 VSS.n1624 0.189974
R35479 VSS.n2202 VSS.n2201 0.189974
R35480 VSS.n2201 VSS.n2200 0.189974
R35481 VSS.n2200 VSS.n2199 0.189974
R35482 VSS.n2199 VSS.n2198 0.189974
R35483 VSS.n2196 VSS.n2195 0.189974
R35484 VSS.n2195 VSS.n2194 0.189974
R35485 VSS.n2194 VSS.n2193 0.189974
R35486 VSS.n1889 VSS.n1888 0.189974
R35487 VSS.n2192 VSS.n1647 0.18275
R35488 VSS.n2191 VSS.n1648 0.18275
R35489 VSS.n2190 VSS.n1649 0.18275
R35490 VSS.n2189 VSS.n1650 0.18275
R35491 VSS.n1792 VSS.n1651 0.18275
R35492 VSS.n1794 VSS.n1793 0.18275
R35493 VSS.n1795 VSS.n1791 0.18275
R35494 VSS.n1700 VSS.n785 0.181684
R35495 VSS.n3203 VSS.n1376 0.1805
R35496 VSS.n3202 VSS.n1379 0.1805
R35497 VSS.n3201 VSS.n1381 0.1805
R35498 VSS.n3200 VSS.n1383 0.1805
R35499 VSS.n3199 VSS.n1385 0.1805
R35500 VSS.n3198 VSS.n1387 0.1805
R35501 VSS.n3197 VSS.n1389 0.1805
R35502 VSS.n3196 VSS.n1391 0.1805
R35503 VSS.n3195 VSS.n1393 0.1805
R35504 VSS.n3194 VSS.n1395 0.1805
R35505 VSS.n3193 VSS.n1397 0.1805
R35506 VSS.n3192 VSS.n1399 0.1805
R35507 VSS.n3191 VSS.n1401 0.1805
R35508 VSS.n3190 VSS.n1403 0.1805
R35509 VSS.n3189 VSS.n1405 0.1805
R35510 VSS.n3204 VSS.n1377 0.1805
R35511 VSS.n3203 VSS.n1378 0.1805
R35512 VSS.n3202 VSS.n1380 0.1805
R35513 VSS.n3201 VSS.n1382 0.1805
R35514 VSS.n3200 VSS.n1384 0.1805
R35515 VSS.n3199 VSS.n1386 0.1805
R35516 VSS.n3198 VSS.n1388 0.1805
R35517 VSS.n3197 VSS.n1390 0.1805
R35518 VSS.n3196 VSS.n1392 0.1805
R35519 VSS.n3195 VSS.n1394 0.1805
R35520 VSS.n3194 VSS.n1396 0.1805
R35521 VSS.n3193 VSS.n1398 0.1805
R35522 VSS.n3192 VSS.n1400 0.1805
R35523 VSS.n3191 VSS.n1402 0.1805
R35524 VSS.n3190 VSS.n1404 0.1805
R35525 VSS.n3189 VSS.n1406 0.1805
R35526 VSS.n3182 VSS.n1404 0.1805
R35527 VSS.n3183 VSS.n1406 0.1805
R35528 VSS.n3182 VSS.n1411 0.1805
R35529 VSS.n3183 VSS.n1410 0.1805
R35530 VSS.n3116 VSS.n1411 0.1805
R35531 VSS.n3115 VSS.n1410 0.1805
R35532 VSS.n3116 VSS.n1413 0.1805
R35533 VSS.n3115 VSS.n1414 0.1805
R35534 VSS.n3108 VSS.n1413 0.1805
R35535 VSS.n3109 VSS.n1414 0.1805
R35536 VSS.n3108 VSS.n1419 0.1805
R35537 VSS.n3109 VSS.n1418 0.1805
R35538 VSS.n3104 VSS.n1419 0.1805
R35539 VSS.n3103 VSS.n1418 0.1805
R35540 VSS.n3104 VSS.n1421 0.1805
R35541 VSS.n3103 VSS.n1422 0.1805
R35542 VSS.n3096 VSS.n1421 0.1805
R35543 VSS.n3096 VSS.n1427 0.1805
R35544 VSS.n3092 VSS.n1427 0.1805
R35545 VSS.n3092 VSS.n1429 0.1805
R35546 VSS.n3090 VSS.n1431 0.1805
R35547 VSS.n3975 VSS.n3916 0.1805
R35548 VSS.n3974 VSS.n3917 0.1805
R35549 VSS.n3973 VSS.n3919 0.1805
R35550 VSS.n3972 VSS.n3921 0.1805
R35551 VSS.n3971 VSS.n3970 0.1805
R35552 VSS.n3969 VSS.n3903 0.1805
R35553 VSS.n3968 VSS.n3902 0.1805
R35554 VSS.n3967 VSS.n3901 0.1805
R35555 VSS.n3966 VSS.n3900 0.1805
R35556 VSS.n3965 VSS.n3899 0.1805
R35557 VSS.n3964 VSS.n3898 0.1805
R35558 VSS.n3999 VSS.n3897 0.1805
R35559 VSS.n4000 VSS.n3895 0.1805
R35560 VSS.n4001 VSS.n3893 0.1805
R35561 VSS.n4002 VSS.n3891 0.1805
R35562 VSS.n4003 VSS.n3889 0.1805
R35563 VSS.n4004 VSS.n3887 0.1805
R35564 VSS.n4005 VSS.n3885 0.1805
R35565 VSS.n4006 VSS.n3883 0.1805
R35566 VSS.n3931 VSS.n3916 0.1805
R35567 VSS.n3930 VSS.n3917 0.1805
R35568 VSS.n3929 VSS.n3919 0.1805
R35569 VSS.n3928 VSS.n3921 0.1805
R35570 VSS.n3970 VSS.n3922 0.1805
R35571 VSS.n3969 VSS.n3923 0.1805
R35572 VSS.n3968 VSS.n3924 0.1805
R35573 VSS.n3967 VSS.n3925 0.1805
R35574 VSS.n3966 VSS.n3926 0.1805
R35575 VSS.n3965 VSS.n3927 0.1805
R35576 VSS.n3964 VSS.n3963 0.1805
R35577 VSS.n3962 VSS.n3897 0.1805
R35578 VSS.n3961 VSS.n3895 0.1805
R35579 VSS.n3960 VSS.n3893 0.1805
R35580 VSS.n3959 VSS.n3891 0.1805
R35581 VSS.n3958 VSS.n3889 0.1805
R35582 VSS.n3957 VSS.n3887 0.1805
R35583 VSS.n3956 VSS.n3885 0.1805
R35584 VSS.n3955 VSS.n3883 0.1805
R35585 VSS.n3954 VSS.n3951 0.1805
R35586 VSS.n3955 VSS.n3950 0.1805
R35587 VSS.n3956 VSS.n3949 0.1805
R35588 VSS.n3957 VSS.n3948 0.1805
R35589 VSS.n3958 VSS.n3947 0.1805
R35590 VSS.n3959 VSS.n3946 0.1805
R35591 VSS.n3960 VSS.n3945 0.1805
R35592 VSS.n3961 VSS.n3944 0.1805
R35593 VSS.n3962 VSS.n3943 0.1805
R35594 VSS.n3963 VSS.n3942 0.1805
R35595 VSS.n3941 VSS.n3927 0.1805
R35596 VSS.n3940 VSS.n3926 0.1805
R35597 VSS.n3939 VSS.n3925 0.1805
R35598 VSS.n3938 VSS.n3924 0.1805
R35599 VSS.n3937 VSS.n3923 0.1805
R35600 VSS.n3936 VSS.n3922 0.1805
R35601 VSS.n3935 VSS.n3928 0.1805
R35602 VSS.n3934 VSS.n3929 0.1805
R35603 VSS.n3933 VSS.n3930 0.1805
R35604 VSS.n4078 VSS.n527 0.1805
R35605 VSS.n4077 VSS.n529 0.1805
R35606 VSS.n4076 VSS.n531 0.1805
R35607 VSS.n4075 VSS.n533 0.1805
R35608 VSS.n4074 VSS.n535 0.1805
R35609 VSS.n4073 VSS.n537 0.1805
R35610 VSS.n4072 VSS.n539 0.1805
R35611 VSS.n4071 VSS.n541 0.1805
R35612 VSS.n4070 VSS.n543 0.1805
R35613 VSS.n4069 VSS.n545 0.1805
R35614 VSS.n4068 VSS.n547 0.1805
R35615 VSS.n4067 VSS.n549 0.1805
R35616 VSS.n4066 VSS.n551 0.1805
R35617 VSS.n4065 VSS.n553 0.1805
R35618 VSS.n4064 VSS.n555 0.1805
R35619 VSS.n4063 VSS.n557 0.1805
R35620 VSS.n4062 VSS.n559 0.1805
R35621 VSS.n4061 VSS.n561 0.1805
R35622 VSS.n4060 VSS.n563 0.1805
R35623 VSS.n4059 VSS.n565 0.1805
R35624 VSS.n4058 VSS.n567 0.1805
R35625 VSS.n4057 VSS.n569 0.1805
R35626 VSS.n4056 VSS.n571 0.1805
R35627 VSS.n4055 VSS.n573 0.1805
R35628 VSS.n4054 VSS.n575 0.1805
R35629 VSS.n4053 VSS.n577 0.1805
R35630 VSS.n4052 VSS.n579 0.1805
R35631 VSS.n4051 VSS.n581 0.1805
R35632 VSS.n4050 VSS.n583 0.1805
R35633 VSS.n4049 VSS.n585 0.1805
R35634 VSS.n4048 VSS.n587 0.1805
R35635 VSS.n4047 VSS.n589 0.1805
R35636 VSS.n4046 VSS.n591 0.1805
R35637 VSS.n4045 VSS.n593 0.1805
R35638 VSS.n4044 VSS.n595 0.1805
R35639 VSS.n4079 VSS.n526 0.1805
R35640 VSS.n4078 VSS.n528 0.1805
R35641 VSS.n4077 VSS.n530 0.1805
R35642 VSS.n4076 VSS.n532 0.1805
R35643 VSS.n4074 VSS.n536 0.1805
R35644 VSS.n4073 VSS.n538 0.1805
R35645 VSS.n4072 VSS.n540 0.1805
R35646 VSS.n4071 VSS.n542 0.1805
R35647 VSS.n4070 VSS.n544 0.1805
R35648 VSS.n4069 VSS.n546 0.1805
R35649 VSS.n4068 VSS.n548 0.1805
R35650 VSS.n4067 VSS.n550 0.1805
R35651 VSS.n4066 VSS.n552 0.1805
R35652 VSS.n4065 VSS.n554 0.1805
R35653 VSS.n4064 VSS.n556 0.1805
R35654 VSS.n4063 VSS.n558 0.1805
R35655 VSS.n4062 VSS.n560 0.1805
R35656 VSS.n4061 VSS.n562 0.1805
R35657 VSS.n4060 VSS.n564 0.1805
R35658 VSS.n4059 VSS.n566 0.1805
R35659 VSS.n4058 VSS.n568 0.1805
R35660 VSS.n4057 VSS.n570 0.1805
R35661 VSS.n4056 VSS.n572 0.1805
R35662 VSS.n4055 VSS.n574 0.1805
R35663 VSS.n4054 VSS.n576 0.1805
R35664 VSS.n4053 VSS.n578 0.1805
R35665 VSS.n4052 VSS.n580 0.1805
R35666 VSS.n4051 VSS.n582 0.1805
R35667 VSS.n4050 VSS.n584 0.1805
R35668 VSS.n4049 VSS.n586 0.1805
R35669 VSS.n4048 VSS.n588 0.1805
R35670 VSS.n4047 VSS.n590 0.1805
R35671 VSS.n4046 VSS.n592 0.1805
R35672 VSS.n4045 VSS.n594 0.1805
R35673 VSS.n4044 VSS.n596 0.1805
R35674 VSS.n4036 VSS.n596 0.1805
R35675 VSS.n4036 VSS.n4035 0.1805
R35676 VSS.n4035 VSS.n603 0.1805
R35677 VSS.n3828 VSS.n603 0.1805
R35678 VSS.n3838 VSS.n3828 0.1805
R35679 VSS.n3838 VSS.n3821 0.1805
R35680 VSS.n3834 VSS.n3821 0.1805
R35681 VSS.n3834 VSS.n3833 0.1805
R35682 VSS.n3833 VSS.n3806 0.1805
R35683 VSS.n3849 VSS.n3806 0.1805
R35684 VSS.n3849 VSS.n3807 0.1805
R35685 VSS.n3807 VSS.n3556 0.1805
R35686 VSS.n3862 VSS.n3556 0.1805
R35687 VSS.n513 VSS.n512 0.1805
R35688 VSS.n632 VSS.n624 0.1805
R35689 VSS.n633 VSS.n625 0.1805
R35690 VSS.n514 VSS.n513 0.1805
R35691 VSS.n647 VSS.n624 0.1805
R35692 VSS.n646 VSS.n625 0.1805
R35693 VSS.n515 VSS.n514 0.1805
R35694 VSS.n648 VSS.n647 0.1805
R35695 VSS.n646 VSS.n623 0.1805
R35696 VSS.n516 VSS.n515 0.1805
R35697 VSS.n652 VSS.n648 0.1805
R35698 VSS.n653 VSS.n623 0.1805
R35699 VSS.n517 VSS.n516 0.1805
R35700 VSS.n652 VSS.n651 0.1805
R35701 VSS.n653 VSS.n621 0.1805
R35702 VSS.n518 VSS.n517 0.1805
R35703 VSS.n651 VSS.n650 0.1805
R35704 VSS.n649 VSS.n621 0.1805
R35705 VSS.n519 VSS.n518 0.1805
R35706 VSS.n650 VSS.n612 0.1805
R35707 VSS.n649 VSS.n613 0.1805
R35708 VSS.n520 VSS.n519 0.1805
R35709 VSS.n662 VSS.n612 0.1805
R35710 VSS.n661 VSS.n613 0.1805
R35711 VSS.n521 VSS.n520 0.1805
R35712 VSS.n663 VSS.n662 0.1805
R35713 VSS.n661 VSS.n611 0.1805
R35714 VSS.n522 VSS.n521 0.1805
R35715 VSS.n670 VSS.n663 0.1805
R35716 VSS.n671 VSS.n611 0.1805
R35717 VSS.n523 VSS.n522 0.1805
R35718 VSS.n670 VSS.n669 0.1805
R35719 VSS.n671 VSS.n609 0.1805
R35720 VSS.n524 VSS.n523 0.1805
R35721 VSS.n669 VSS.n668 0.1805
R35722 VSS.n667 VSS.n609 0.1805
R35723 VSS.n665 VSS.n532 0.1805
R35724 VSS.n525 VSS.n524 0.1805
R35725 VSS.n526 VSS.n525 0.1805
R35726 VSS.n668 VSS.n664 0.1805
R35727 VSS.n664 VSS.n528 0.1805
R35728 VSS.n667 VSS.n666 0.1805
R35729 VSS.n666 VSS.n530 0.1805
R35730 VSS.n673 VSS.n607 0.1805
R35731 VSS.n665 VSS.n607 0.1805
R35732 VSS.n672 VSS.n610 0.1805
R35733 VSS.n673 VSS.n672 0.1805
R35734 VSS.n660 VSS.n614 0.1805
R35735 VSS.n660 VSS.n610 0.1805
R35736 VSS.n655 VSS.n619 0.1805
R35737 VSS.n619 VSS.n614 0.1805
R35738 VSS.n654 VSS.n622 0.1805
R35739 VSS.n655 VSS.n654 0.1805
R35740 VSS.n645 VSS.n626 0.1805
R35741 VSS.n645 VSS.n622 0.1805
R35742 VSS.n629 VSS.n505 0.1805
R35743 VSS.n4098 VSS.n511 0.1805
R35744 VSS.n512 VSS.n511 0.1805
R35745 VSS.n631 VSS.n509 0.1805
R35746 VSS.n632 VSS.n631 0.1805
R35747 VSS.n630 VSS.n507 0.1805
R35748 VSS.n633 VSS.n630 0.1805
R35749 VSS.n634 VSS.n629 0.1805
R35750 VSS.n634 VSS.n626 0.1805
R35751 VSS.n4099 VSS.n4098 0.1805
R35752 VSS.n4100 VSS.n508 0.1805
R35753 VSS.n4100 VSS.n509 0.1805
R35754 VSS.n4101 VSS.n506 0.1805
R35755 VSS.n4101 VSS.n507 0.1805
R35756 VSS.n4102 VSS.n504 0.1805
R35757 VSS.n4102 VSS.n505 0.1805
R35758 VSS.n4103 VSS.n502 0.1805
R35759 VSS.n4103 VSS.n503 0.1805
R35760 VSS.n4104 VSS.n500 0.1805
R35761 VSS.n4104 VSS.n501 0.1805
R35762 VSS.n4105 VSS.n498 0.1805
R35763 VSS.n4105 VSS.n499 0.1805
R35764 VSS.n4106 VSS.n496 0.1805
R35765 VSS.n4106 VSS.n497 0.1805
R35766 VSS.n4107 VSS.n494 0.1805
R35767 VSS.n4107 VSS.n495 0.1805
R35768 VSS.n4108 VSS.n492 0.1805
R35769 VSS.n4108 VSS.n493 0.1805
R35770 VSS.n4109 VSS.n490 0.1805
R35771 VSS.n4109 VSS.n491 0.1805
R35772 VSS.n4110 VSS.n488 0.1805
R35773 VSS.n4110 VSS.n489 0.1805
R35774 VSS.n4111 VSS.n486 0.1805
R35775 VSS.n4111 VSS.n487 0.1805
R35776 VSS.n4112 VSS.n485 0.1805
R35777 VSS.n4112 VSS.n461 0.1805
R35778 VSS.n4131 VSS.n4113 0.1805
R35779 VSS.n4113 VSS.n462 0.1805
R35780 VSS.n4114 VSS.n463 0.1805
R35781 VSS.n4115 VSS.n464 0.1805
R35782 VSS.n4151 VSS.n466 0.1805
R35783 VSS.n4130 VSS.n4114 0.1805
R35784 VSS.n4129 VSS.n4115 0.1805
R35785 VSS.n4128 VSS.n466 0.1805
R35786 VSS.n4130 VSS.n484 0.1805
R35787 VSS.n4129 VSS.n4116 0.1805
R35788 VSS.n4128 VSS.n4117 0.1805
R35789 VSS.n484 VSS.n483 0.1805
R35790 VSS.n4120 VSS.n4116 0.1805
R35791 VSS.n4121 VSS.n4117 0.1805
R35792 VSS.n483 VSS.n480 0.1805
R35793 VSS.n4120 VSS.n478 0.1805
R35794 VSS.n4121 VSS.n477 0.1805
R35795 VSS.n4137 VSS.n480 0.1805
R35796 VSS.n4138 VSS.n478 0.1805
R35797 VSS.n4139 VSS.n477 0.1805
R35798 VSS.n4137 VSS.n481 0.1805
R35799 VSS.n4138 VSS.n479 0.1805
R35800 VSS.n4139 VSS.n475 0.1805
R35801 VSS.n3981 VSS.n481 0.1805
R35802 VSS.n3980 VSS.n479 0.1805
R35803 VSS.n3979 VSS.n475 0.1805
R35804 VSS.n3981 VSS.n3912 0.1805
R35805 VSS.n3980 VSS.n3910 0.1805
R35806 VSS.n3979 VSS.n3909 0.1805
R35807 VSS.n3985 VSS.n3912 0.1805
R35808 VSS.n3986 VSS.n3910 0.1805
R35809 VSS.n3987 VSS.n3909 0.1805
R35810 VSS.n3985 VSS.n3913 0.1805
R35811 VSS.n3986 VSS.n3911 0.1805
R35812 VSS.n3973 VSS.n3920 0.1805
R35813 VSS.n3975 VSS.n3914 0.1805
R35814 VSS.n3914 VSS.n3913 0.1805
R35815 VSS.n3974 VSS.n3918 0.1805
R35816 VSS.n3918 VSS.n3911 0.1805
R35817 VSS.n3972 VSS.n3905 0.1805
R35818 VSS.n3989 VSS.n3905 0.1805
R35819 VSS.n3920 VSS.n3906 0.1805
R35820 VSS.n3987 VSS.n3906 0.1805
R35821 VSS.n3989 VSS.n3988 0.1805
R35822 VSS.n3988 VSS.n3908 0.1805
R35823 VSS.n3908 VSS.n474 0.1805
R35824 VSS.n4141 VSS.n474 0.1805
R35825 VSS.n4141 VSS.n4140 0.1805
R35826 VSS.n4140 VSS.n476 0.1805
R35827 VSS.n4122 VSS.n476 0.1805
R35828 VSS.n4122 VSS.n4118 0.1805
R35829 VSS.n4127 VSS.n4118 0.1805
R35830 VSS.n4127 VSS.n467 0.1805
R35831 VSS.n4150 VSS.n467 0.1805
R35832 VSS.n4148 VSS.n469 0.1805
R35833 VSS.n3862 VSS.n3554 0.1805
R35834 VSS.n3859 VSS.n3858 0.1805
R35835 VSS.n3858 VSS.n714 0.1805
R35836 VSS.n4013 VSS.n3879 0.1805
R35837 VSS.n4013 VSS.n3877 0.1805
R35838 VSS.n4017 VSS.n3877 0.1805
R35839 VSS.n4018 VSS.n4017 0.1805
R35840 VSS.n4018 VSS.n712 0.1805
R35841 VSS.n4022 VSS.n712 0.1805
R35842 VSS.n3450 VSS.n870 0.1805
R35843 VSS.n3451 VSS.n868 0.1805
R35844 VSS.n3452 VSS.n866 0.1805
R35845 VSS.n3453 VSS.n864 0.1805
R35846 VSS.n3454 VSS.n862 0.1805
R35847 VSS.n3455 VSS.n860 0.1805
R35848 VSS.n3456 VSS.n858 0.1805
R35849 VSS.n3457 VSS.n856 0.1805
R35850 VSS.n3458 VSS.n854 0.1805
R35851 VSS.n3459 VSS.n852 0.1805
R35852 VSS.n3460 VSS.n850 0.1805
R35853 VSS.n3461 VSS.n848 0.1805
R35854 VSS.n3462 VSS.n846 0.1805
R35855 VSS.n3463 VSS.n844 0.1805
R35856 VSS.n3464 VSS.n842 0.1805
R35857 VSS.n3465 VSS.n840 0.1805
R35858 VSS.n3466 VSS.n838 0.1805
R35859 VSS.n3467 VSS.n836 0.1805
R35860 VSS.n3468 VSS.n834 0.1805
R35861 VSS.n3469 VSS.n832 0.1805
R35862 VSS.n3470 VSS.n830 0.1805
R35863 VSS.n3471 VSS.n828 0.1805
R35864 VSS.n3472 VSS.n826 0.1805
R35865 VSS.n3473 VSS.n824 0.1805
R35866 VSS.n3474 VSS.n822 0.1805
R35867 VSS.n3475 VSS.n820 0.1805
R35868 VSS.n3476 VSS.n818 0.1805
R35869 VSS.n3477 VSS.n816 0.1805
R35870 VSS.n3478 VSS.n815 0.1805
R35871 VSS.n3449 VSS.n3448 0.1805
R35872 VSS.n3450 VSS.n871 0.1805
R35873 VSS.n3451 VSS.n869 0.1805
R35874 VSS.n3452 VSS.n867 0.1805
R35875 VSS.n3453 VSS.n865 0.1805
R35876 VSS.n3454 VSS.n863 0.1805
R35877 VSS.n3455 VSS.n861 0.1805
R35878 VSS.n3456 VSS.n859 0.1805
R35879 VSS.n3457 VSS.n857 0.1805
R35880 VSS.n3458 VSS.n855 0.1805
R35881 VSS.n3459 VSS.n853 0.1805
R35882 VSS.n3460 VSS.n851 0.1805
R35883 VSS.n3461 VSS.n849 0.1805
R35884 VSS.n3462 VSS.n847 0.1805
R35885 VSS.n3463 VSS.n845 0.1805
R35886 VSS.n3464 VSS.n843 0.1805
R35887 VSS.n3465 VSS.n841 0.1805
R35888 VSS.n3466 VSS.n839 0.1805
R35889 VSS.n3467 VSS.n837 0.1805
R35890 VSS.n3468 VSS.n835 0.1805
R35891 VSS.n3469 VSS.n833 0.1805
R35892 VSS.n3470 VSS.n831 0.1805
R35893 VSS.n3471 VSS.n829 0.1805
R35894 VSS.n3472 VSS.n827 0.1805
R35895 VSS.n3473 VSS.n825 0.1805
R35896 VSS.n3474 VSS.n823 0.1805
R35897 VSS.n3475 VSS.n821 0.1805
R35898 VSS.n3476 VSS.n819 0.1805
R35899 VSS.n3477 VSS.n817 0.1805
R35900 VSS.n3478 VSS.n813 0.1805
R35901 VSS.n3448 VSS.n873 0.1805
R35902 VSS.n966 VSS.n871 0.1805
R35903 VSS.n967 VSS.n869 0.1805
R35904 VSS.n968 VSS.n867 0.1805
R35905 VSS.n969 VSS.n865 0.1805
R35906 VSS.n970 VSS.n863 0.1805
R35907 VSS.n971 VSS.n861 0.1805
R35908 VSS.n972 VSS.n859 0.1805
R35909 VSS.n973 VSS.n857 0.1805
R35910 VSS.n974 VSS.n855 0.1805
R35911 VSS.n975 VSS.n853 0.1805
R35912 VSS.n976 VSS.n851 0.1805
R35913 VSS.n977 VSS.n849 0.1805
R35914 VSS.n978 VSS.n847 0.1805
R35915 VSS.n979 VSS.n845 0.1805
R35916 VSS.n980 VSS.n843 0.1805
R35917 VSS.n981 VSS.n841 0.1805
R35918 VSS.n982 VSS.n839 0.1805
R35919 VSS.n983 VSS.n837 0.1805
R35920 VSS.n984 VSS.n835 0.1805
R35921 VSS.n985 VSS.n833 0.1805
R35922 VSS.n986 VSS.n831 0.1805
R35923 VSS.n987 VSS.n829 0.1805
R35924 VSS.n988 VSS.n827 0.1805
R35925 VSS.n989 VSS.n825 0.1805
R35926 VSS.n990 VSS.n823 0.1805
R35927 VSS.n991 VSS.n821 0.1805
R35928 VSS.n992 VSS.n819 0.1805
R35929 VSS.n993 VSS.n817 0.1805
R35930 VSS.n994 VSS.n813 0.1805
R35931 VSS.n874 VSS.n873 0.1805
R35932 VSS.n966 VSS.n965 0.1805
R35933 VSS.n967 VSS.n924 0.1805
R35934 VSS.n968 VSS.n923 0.1805
R35935 VSS.n969 VSS.n922 0.1805
R35936 VSS.n970 VSS.n921 0.1805
R35937 VSS.n971 VSS.n920 0.1805
R35938 VSS.n972 VSS.n919 0.1805
R35939 VSS.n973 VSS.n918 0.1805
R35940 VSS.n974 VSS.n917 0.1805
R35941 VSS.n975 VSS.n916 0.1805
R35942 VSS.n976 VSS.n915 0.1805
R35943 VSS.n977 VSS.n914 0.1805
R35944 VSS.n978 VSS.n913 0.1805
R35945 VSS.n979 VSS.n911 0.1805
R35946 VSS.n1009 VSS.n980 0.1805
R35947 VSS.n1008 VSS.n981 0.1805
R35948 VSS.n1007 VSS.n982 0.1805
R35949 VSS.n1006 VSS.n983 0.1805
R35950 VSS.n1005 VSS.n984 0.1805
R35951 VSS.n1004 VSS.n985 0.1805
R35952 VSS.n1003 VSS.n986 0.1805
R35953 VSS.n1002 VSS.n987 0.1805
R35954 VSS.n1001 VSS.n988 0.1805
R35955 VSS.n1000 VSS.n989 0.1805
R35956 VSS.n999 VSS.n990 0.1805
R35957 VSS.n998 VSS.n991 0.1805
R35958 VSS.n997 VSS.n992 0.1805
R35959 VSS.n996 VSS.n993 0.1805
R35960 VSS.n995 VSS.n994 0.1805
R35961 VSS.n875 VSS.n874 0.1805
R35962 VSS.n965 VSS.n964 0.1805
R35963 VSS.n963 VSS.n924 0.1805
R35964 VSS.n962 VSS.n923 0.1805
R35965 VSS.n961 VSS.n922 0.1805
R35966 VSS.n960 VSS.n921 0.1805
R35967 VSS.n959 VSS.n920 0.1805
R35968 VSS.n958 VSS.n919 0.1805
R35969 VSS.n957 VSS.n918 0.1805
R35970 VSS.n956 VSS.n917 0.1805
R35971 VSS.n955 VSS.n916 0.1805
R35972 VSS.n954 VSS.n915 0.1805
R35973 VSS.n953 VSS.n914 0.1805
R35974 VSS.n913 VSS.n912 0.1805
R35975 VSS.n1011 VSS.n911 0.1805
R35976 VSS.n1010 VSS.n1009 0.1805
R35977 VSS.n1008 VSS.n779 0.1805
R35978 VSS.n1007 VSS.n781 0.1805
R35979 VSS.n1006 VSS.n782 0.1805
R35980 VSS.n1005 VSS.n784 0.1805
R35981 VSS.n1004 VSS.n786 0.1805
R35982 VSS.n1003 VSS.n788 0.1805
R35983 VSS.n1002 VSS.n790 0.1805
R35984 VSS.n1001 VSS.n792 0.1805
R35985 VSS.n1000 VSS.n794 0.1805
R35986 VSS.n999 VSS.n796 0.1805
R35987 VSS.n998 VSS.n798 0.1805
R35988 VSS.n997 VSS.n800 0.1805
R35989 VSS.n996 VSS.n802 0.1805
R35990 VSS.n995 VSS.n803 0.1805
R35991 VSS.n876 VSS.n875 0.1805
R35992 VSS.n964 VSS.n925 0.1805
R35993 VSS.n963 VSS.n952 0.1805
R35994 VSS.n962 VSS.n900 0.1805
R35995 VSS.n961 VSS.n901 0.1805
R35996 VSS.n960 VSS.n902 0.1805
R35997 VSS.n959 VSS.n903 0.1805
R35998 VSS.n958 VSS.n904 0.1805
R35999 VSS.n957 VSS.n905 0.1805
R36000 VSS.n956 VSS.n906 0.1805
R36001 VSS.n955 VSS.n907 0.1805
R36002 VSS.n954 VSS.n908 0.1805
R36003 VSS.n953 VSS.n909 0.1805
R36004 VSS.n912 VSS.n910 0.1805
R36005 VSS.n1012 VSS.n1011 0.1805
R36006 VSS.n1010 VSS.n780 0.1805
R36007 VSS.n3502 VSS.n779 0.1805
R36008 VSS.n3501 VSS.n781 0.1805
R36009 VSS.n3500 VSS.n782 0.1805
R36010 VSS.n3499 VSS.n784 0.1805
R36011 VSS.n3498 VSS.n786 0.1805
R36012 VSS.n3497 VSS.n788 0.1805
R36013 VSS.n3496 VSS.n790 0.1805
R36014 VSS.n3495 VSS.n792 0.1805
R36015 VSS.n3494 VSS.n794 0.1805
R36016 VSS.n3493 VSS.n796 0.1805
R36017 VSS.n3492 VSS.n798 0.1805
R36018 VSS.n3491 VSS.n800 0.1805
R36019 VSS.n3489 VSS.n803 0.1805
R36020 VSS.n3489 VSS.n804 0.1805
R36021 VSS.n1750 VSS.n804 0.1805
R36022 VSS.n1750 VSS.n1705 0.1805
R36023 VSS.n1740 VSS.n1705 0.1805
R36024 VSS.n1740 VSS.n1712 0.1805
R36025 VSS.n1735 VSS.n1712 0.1805
R36026 VSS.n1735 VSS.n1714 0.1805
R36027 VSS.n1727 VSS.n1714 0.1805
R36028 VSS.n1727 VSS.n1723 0.1805
R36029 VSS.n1723 VSS.n1685 0.1805
R36030 VSS.n1825 VSS.n1685 0.1805
R36031 VSS.n1825 VSS.n1683 0.1805
R36032 VSS.n1821 VSS.n1683 0.1805
R36033 VSS.n1821 VSS.n1820 0.1805
R36034 VSS.n1829 VSS.n1680 0.1805
R36035 VSS.n1820 VSS.n1688 0.1805
R36036 VSS.n1819 VSS.n1818 0.1805
R36037 VSS.n1817 VSS.n1680 0.1805
R36038 VSS.n1816 VSS.n1679 0.1805
R36039 VSS.n1815 VSS.n1677 0.1805
R36040 VSS.n1814 VSS.n1676 0.1805
R36041 VSS.n1813 VSS.n1675 0.1805
R36042 VSS.n1812 VSS.n1674 0.1805
R36043 VSS.n1811 VSS.n1673 0.1805
R36044 VSS.n1810 VSS.n1672 0.1805
R36045 VSS.n1809 VSS.n1671 0.1805
R36046 VSS.n1808 VSS.n1670 0.1805
R36047 VSS.n1807 VSS.n1669 0.1805
R36048 VSS.n1806 VSS.n1668 0.1805
R36049 VSS.n1805 VSS.n1666 0.1805
R36050 VSS.n1804 VSS.n1665 0.1805
R36051 VSS.n3517 VSS.n767 0.1805
R36052 VSS.n766 VSS.n765 0.1805
R36053 VSS.n3513 VSS.n767 0.1805
R36054 VSS.n3543 VSS.n722 0.1805
R36055 VSS.n740 VSS.n718 0.1805
R36056 VSS.n3547 VSS.n718 0.1805
R36057 VSS.n741 VSS.n719 0.1805
R36058 VSS.n3546 VSS.n719 0.1805
R36059 VSS.n742 VSS.n720 0.1805
R36060 VSS.n3545 VSS.n720 0.1805
R36061 VSS.n743 VSS.n721 0.1805
R36062 VSS.n3544 VSS.n721 0.1805
R36063 VSS.n745 VSS.n723 0.1805
R36064 VSS.n3542 VSS.n723 0.1805
R36065 VSS.n746 VSS.n724 0.1805
R36066 VSS.n3541 VSS.n724 0.1805
R36067 VSS.n747 VSS.n725 0.1805
R36068 VSS.n3540 VSS.n725 0.1805
R36069 VSS.n748 VSS.n726 0.1805
R36070 VSS.n3539 VSS.n726 0.1805
R36071 VSS.n749 VSS.n727 0.1805
R36072 VSS.n3538 VSS.n727 0.1805
R36073 VSS.n750 VSS.n728 0.1805
R36074 VSS.n3537 VSS.n728 0.1805
R36075 VSS.n751 VSS.n730 0.1805
R36076 VSS.n3535 VSS.n730 0.1805
R36077 VSS.n752 VSS.n731 0.1805
R36078 VSS.n753 VSS.n733 0.1805
R36079 VSS.n3534 VSS.n731 0.1805
R36080 VSS.n3533 VSS.n733 0.1805
R36081 VSS.n952 VSS.n951 0.1805
R36082 VSS.n878 VSS.n877 0.1805
R36083 VSS.n877 VSS.n876 0.1805
R36084 VSS.n950 VSS.n949 0.1805
R36085 VSS.n950 VSS.n925 0.1805
R36086 VSS.n879 VSS.n878 0.1805
R36087 VSS.n949 VSS.n948 0.1805
R36088 VSS.n880 VSS.n879 0.1805
R36089 VSS.n948 VSS.n926 0.1805
R36090 VSS.n881 VSS.n880 0.1805
R36091 VSS.n930 VSS.n926 0.1805
R36092 VSS.n882 VSS.n881 0.1805
R36093 VSS.n940 VSS.n930 0.1805
R36094 VSS.n883 VSS.n882 0.1805
R36095 VSS.n940 VSS.n939 0.1805
R36096 VSS.n884 VSS.n883 0.1805
R36097 VSS.n939 VSS.n938 0.1805
R36098 VSS.n885 VSS.n884 0.1805
R36099 VSS.n938 VSS.n931 0.1805
R36100 VSS.n886 VSS.n885 0.1805
R36101 VSS.n932 VSS.n931 0.1805
R36102 VSS.n887 VSS.n886 0.1805
R36103 VSS.n932 VSS.n888 0.1805
R36104 VSS.n3430 VSS.n887 0.1805
R36105 VSS.n3429 VSS.n888 0.1805
R36106 VSS.n3532 VSS.n735 0.1805
R36107 VSS.n3534 VSS.n732 0.1805
R36108 VSS.n3430 VSS.n732 0.1805
R36109 VSS.n3533 VSS.n734 0.1805
R36110 VSS.n3429 VSS.n734 0.1805
R36111 VSS.n3428 VSS.n735 0.1805
R36112 VSS.n3428 VSS.n889 0.1805
R36113 VSS.n933 VSS.n889 0.1805
R36114 VSS.n934 VSS.n933 0.1805
R36115 VSS.n937 VSS.n934 0.1805
R36116 VSS.n937 VSS.n929 0.1805
R36117 VSS.n941 VSS.n929 0.1805
R36118 VSS.n941 VSS.n927 0.1805
R36119 VSS.n946 VSS.n927 0.1805
R36120 VSS.n947 VSS.n946 0.1805
R36121 VSS.n947 VSS.n899 0.1805
R36122 VSS.n951 VSS.n899 0.1805
R36123 VSS.n3505 VSS.n3504 0.1805
R36124 VSS.n3531 VSS.n3530 0.1805
R36125 VSS.n3532 VSS.n3531 0.1805
R36126 VSS.n744 VSS.n722 0.1805
R36127 VSS.n3515 VSS.n3514 0.1805
R36128 VSS.n1809 VSS.n1782 0.1805
R36129 VSS.n1810 VSS.n1781 0.1805
R36130 VSS.n1811 VSS.n1780 0.1805
R36131 VSS.n1812 VSS.n1779 0.1805
R36132 VSS.n1813 VSS.n1778 0.1805
R36133 VSS.n1814 VSS.n1777 0.1805
R36134 VSS.n1815 VSS.n1776 0.1805
R36135 VSS.n1816 VSS.n1775 0.1805
R36136 VSS.n1817 VSS.n1774 0.1805
R36137 VSS.n1818 VSS.n1773 0.1805
R36138 VSS.n2214 VSS.n1645 0.1805
R36139 VSS.n2215 VSS.n1644 0.1805
R36140 VSS.n2216 VSS.n1643 0.1805
R36141 VSS.n2217 VSS.n1642 0.1805
R36142 VSS.n2218 VSS.n1641 0.1805
R36143 VSS.n2219 VSS.n1640 0.1805
R36144 VSS.n2220 VSS.n1639 0.1805
R36145 VSS.n2221 VSS.n1638 0.1805
R36146 VSS.n2222 VSS.n1637 0.1805
R36147 VSS.n2223 VSS.n1626 0.1805
R36148 VSS.n2224 VSS.n1628 0.1805
R36149 VSS.n2225 VSS.n1629 0.1805
R36150 VSS.n2226 VSS.n1631 0.1805
R36151 VSS.n2227 VSS.n1633 0.1805
R36152 VSS.n2212 VSS.n2211 0.1805
R36153 VSS.n2210 VSS.n1645 0.1805
R36154 VSS.n2209 VSS.n1644 0.1805
R36155 VSS.n2208 VSS.n1643 0.1805
R36156 VSS.n2207 VSS.n1642 0.1805
R36157 VSS.n2206 VSS.n1641 0.1805
R36158 VSS.n2205 VSS.n1640 0.1805
R36159 VSS.n2204 VSS.n1639 0.1805
R36160 VSS.n2203 VSS.n1638 0.1805
R36161 VSS.n1637 VSS.n1627 0.1805
R36162 VSS.n2235 VSS.n1626 0.1805
R36163 VSS.n2234 VSS.n1628 0.1805
R36164 VSS.n2233 VSS.n1629 0.1805
R36165 VSS.n2232 VSS.n1631 0.1805
R36166 VSS.n2232 VSS.n1632 0.1805
R36167 VSS.n2065 VSS.n1632 0.1805
R36168 VSS.n2065 VSS.n2059 0.1805
R36169 VSS.n2074 VSS.n2059 0.1805
R36170 VSS.n2074 VSS.n2057 0.1805
R36171 VSS.n2084 VSS.n2057 0.1805
R36172 VSS.n2084 VSS.n2055 0.1805
R36173 VSS.n2080 VSS.n2055 0.1805
R36174 VSS.n2080 VSS.n2079 0.1805
R36175 VSS.n2079 VSS.n2040 0.1805
R36176 VSS.n2095 VSS.n2040 0.1805
R36177 VSS.n2095 VSS.n2041 0.1805
R36178 VSS.n2041 VSS.n2036 0.1805
R36179 VSS.n2111 VSS.n2036 0.1805
R36180 VSS.n2111 VSS.n2034 0.1805
R36181 VSS.n2103 VSS.n2034 0.1805
R36182 VSS.n2103 VSS.n2102 0.1805
R36183 VSS.n2102 VSS.n2009 0.1805
R36184 VSS.n2122 VSS.n2009 0.1805
R36185 VSS.n2122 VSS.n2010 0.1805
R36186 VSS.n2023 VSS.n2010 0.1805
R36187 VSS.n2023 VSS.n2020 0.1805
R36188 VSS.n2020 VSS.n1998 0.1805
R36189 VSS.n2130 VSS.n1998 0.1805
R36190 VSS.n2130 VSS.n1996 0.1805
R36191 VSS.n2001 VSS.n1996 0.1805
R36192 VSS.n2001 VSS.n1945 0.1805
R36193 VSS.n2140 VSS.n1945 0.1805
R36194 VSS.n2139 VSS.n1947 0.1805
R36195 VSS.n2157 VSS.n1856 0.1805
R36196 VSS.n2156 VSS.n1857 0.1805
R36197 VSS.n2155 VSS.n1859 0.1805
R36198 VSS.n2154 VSS.n1861 0.1805
R36199 VSS.n2152 VSS.n1864 0.1805
R36200 VSS.n2151 VSS.n1920 0.1805
R36201 VSS.n2150 VSS.n1922 0.1805
R36202 VSS.n2149 VSS.n1924 0.1805
R36203 VSS.n2148 VSS.n1928 0.1805
R36204 VSS.n2147 VSS.n1930 0.1805
R36205 VSS.n2146 VSS.n1932 0.1805
R36206 VSS.n2145 VSS.n1934 0.1805
R36207 VSS.n2144 VSS.n1936 0.1805
R36208 VSS.n2143 VSS.n1938 0.1805
R36209 VSS.n2142 VSS.n1941 0.1805
R36210 VSS.n2141 VSS.n1943 0.1805
R36211 VSS.n2140 VSS.n1946 0.1805
R36212 VSS.n2139 VSS.n1948 0.1805
R36213 VSS.n1969 VSS.n1856 0.1805
R36214 VSS.n1970 VSS.n1857 0.1805
R36215 VSS.n1971 VSS.n1859 0.1805
R36216 VSS.n1972 VSS.n1861 0.1805
R36217 VSS.n1973 VSS.n1863 0.1805
R36218 VSS.n1974 VSS.n1864 0.1805
R36219 VSS.n1975 VSS.n1920 0.1805
R36220 VSS.n1976 VSS.n1922 0.1805
R36221 VSS.n1977 VSS.n1924 0.1805
R36222 VSS.n1978 VSS.n1928 0.1805
R36223 VSS.n1979 VSS.n1930 0.1805
R36224 VSS.n1980 VSS.n1932 0.1805
R36225 VSS.n1981 VSS.n1934 0.1805
R36226 VSS.n1982 VSS.n1936 0.1805
R36227 VSS.n1983 VSS.n1938 0.1805
R36228 VSS.n1984 VSS.n1941 0.1805
R36229 VSS.n1985 VSS.n1943 0.1805
R36230 VSS.n1986 VSS.n1946 0.1805
R36231 VSS.n2176 VSS.n1666 0.1805
R36232 VSS.n2177 VSS.n1665 0.1805
R36233 VSS.n2176 VSS.n1667 0.1805
R36234 VSS.n2177 VSS.n1663 0.1805
R36235 VSS.n1841 VSS.n1667 0.1805
R36236 VSS.n1883 VSS.n1663 0.1805
R36237 VSS.n1842 VSS.n1841 0.1805
R36238 VSS.n1884 VSS.n1883 0.1805
R36239 VSS.n2181 VSS.n1660 0.1805
R36240 VSS.n1843 VSS.n1842 0.1805
R36241 VSS.n1885 VSS.n1884 0.1805
R36242 VSS.n1886 VSS.n1882 0.1805
R36243 VSS.n1844 VSS.n1843 0.1805
R36244 VSS.n1885 VSS.n1876 0.1805
R36245 VSS.n1886 VSS.n1877 0.1805
R36246 VSS.n1845 VSS.n1844 0.1805
R36247 VSS.n1894 VSS.n1876 0.1805
R36248 VSS.n1893 VSS.n1877 0.1805
R36249 VSS.n1846 VSS.n1845 0.1805
R36250 VSS.n1895 VSS.n1894 0.1805
R36251 VSS.n1893 VSS.n1875 0.1805
R36252 VSS.n1847 VSS.n1846 0.1805
R36253 VSS.n1905 VSS.n1895 0.1805
R36254 VSS.n1906 VSS.n1875 0.1805
R36255 VSS.n1848 VSS.n1847 0.1805
R36256 VSS.n1905 VSS.n1904 0.1805
R36257 VSS.n1906 VSS.n1873 0.1805
R36258 VSS.n1849 VSS.n1848 0.1805
R36259 VSS.n1904 VSS.n1903 0.1805
R36260 VSS.n1902 VSS.n1873 0.1805
R36261 VSS.n1850 VSS.n1849 0.1805
R36262 VSS.n1903 VSS.n1900 0.1805
R36263 VSS.n1902 VSS.n1901 0.1805
R36264 VSS.n1851 VSS.n1850 0.1805
R36265 VSS.n1900 VSS.n1899 0.1805
R36266 VSS.n1901 VSS.n1870 0.1805
R36267 VSS.n1852 VSS.n1851 0.1805
R36268 VSS.n1899 VSS.n1898 0.1805
R36269 VSS.n1870 VSS.n1868 0.1805
R36270 VSS.n1853 VSS.n1852 0.1805
R36271 VSS.n1898 VSS.n1897 0.1805
R36272 VSS.n1896 VSS.n1868 0.1805
R36273 VSS.n2154 VSS.n1862 0.1805
R36274 VSS.n1854 VSS.n1853 0.1805
R36275 VSS.n2157 VSS.n1854 0.1805
R36276 VSS.n1897 VSS.n1858 0.1805
R36277 VSS.n2156 VSS.n1858 0.1805
R36278 VSS.n1896 VSS.n1860 0.1805
R36279 VSS.n2155 VSS.n1860 0.1805
R36280 VSS.n1914 VSS.n1865 0.1805
R36281 VSS.n1865 VSS.n1862 0.1805
R36282 VSS.n1913 VSS.n1869 0.1805
R36283 VSS.n1914 VSS.n1913 0.1805
R36284 VSS.n1908 VSS.n1871 0.1805
R36285 VSS.n1871 VSS.n1869 0.1805
R36286 VSS.n1907 VSS.n1874 0.1805
R36287 VSS.n1908 VSS.n1907 0.1805
R36288 VSS.n1892 VSS.n1878 0.1805
R36289 VSS.n1892 VSS.n1874 0.1805
R36290 VSS.n1887 VSS.n1660 0.1805
R36291 VSS.n1887 VSS.n1878 0.1805
R36292 VSS.n2179 VSS.n1661 0.1805
R36293 VSS.n1882 VSS.n1661 0.1805
R36294 VSS.n2180 VSS.n1662 0.1805
R36295 VSS.n2181 VSS.n2180 0.1805
R36296 VSS.n2178 VSS.n1664 0.1805
R36297 VSS.n2179 VSS.n2178 0.1805
R36298 VSS.n1830 VSS.n1679 0.1805
R36299 VSS.n1832 VSS.n1677 0.1805
R36300 VSS.n1833 VSS.n1676 0.1805
R36301 VSS.n1834 VSS.n1675 0.1805
R36302 VSS.n1835 VSS.n1674 0.1805
R36303 VSS.n1836 VSS.n1673 0.1805
R36304 VSS.n1837 VSS.n1672 0.1805
R36305 VSS.n1838 VSS.n1671 0.1805
R36306 VSS.n1839 VSS.n1670 0.1805
R36307 VSS.n1840 VSS.n1669 0.1805
R36308 VSS.n2175 VSS.n1668 0.1805
R36309 VSS.n1970 VSS.n1967 0.1805
R36310 VSS.n1971 VSS.n1966 0.1805
R36311 VSS.n1972 VSS.n1965 0.1805
R36312 VSS.n1973 VSS.n1964 0.1805
R36313 VSS.n1974 VSS.n1963 0.1805
R36314 VSS.n1975 VSS.n1962 0.1805
R36315 VSS.n1976 VSS.n1961 0.1805
R36316 VSS.n1977 VSS.n1960 0.1805
R36317 VSS.n1978 VSS.n1959 0.1805
R36318 VSS.n1979 VSS.n1958 0.1805
R36319 VSS.n1980 VSS.n1957 0.1805
R36320 VSS.n1981 VSS.n1956 0.1805
R36321 VSS.n1982 VSS.n1955 0.1805
R36322 VSS.n1983 VSS.n1954 0.1805
R36323 VSS.n1984 VSS.n1953 0.1805
R36324 VSS.n1985 VSS.n1952 0.1805
R36325 VSS.n1986 VSS.n1951 0.1805
R36326 VSS.n1987 VSS.n1948 0.1805
R36327 VSS.n1987 VSS.n1950 0.1805
R36328 VSS.n2138 VSS.n1949 0.1805
R36329 VSS.n1988 VSS.n1949 0.1805
R36330 VSS.n2153 VSS.n1863 0.1805
R36331 VSS.n2137 VSS.n1992 0.1805
R36332 VSS.n2138 VSS.n2137 0.1805
R36333 VSS.n2132 VSS.n1995 0.1805
R36334 VSS.n1995 VSS.n1947 0.1805
R36335 VSS.n2133 VSS.n1994 0.1805
R36336 VSS.n2133 VSS.n1992 0.1805
R36337 VSS.n2131 VSS.n1997 0.1805
R36338 VSS.n2132 VSS.n2131 0.1805
R36339 VSS.n2018 VSS.n2015 0.1805
R36340 VSS.n2015 VSS.n1994 0.1805
R36341 VSS.n2024 VSS.n2019 0.1805
R36342 VSS.n2019 VSS.n1997 0.1805
R36343 VSS.n2026 VSS.n2025 0.1805
R36344 VSS.n2025 VSS.n2018 0.1805
R36345 VSS.n2121 VSS.n2011 0.1805
R36346 VSS.n2024 VSS.n2011 0.1805
R36347 VSS.n2119 VSS.n2012 0.1805
R36348 VSS.n2026 VSS.n2012 0.1805
R36349 VSS.n2120 VSS.n2013 0.1805
R36350 VSS.n2121 VSS.n2120 0.1805
R36351 VSS.n2118 VSS.n2030 0.1805
R36352 VSS.n2119 VSS.n2118 0.1805
R36353 VSS.n2113 VSS.n2033 0.1805
R36354 VSS.n2033 VSS.n2013 0.1805
R36355 VSS.n2114 VSS.n2032 0.1805
R36356 VSS.n2114 VSS.n2030 0.1805
R36357 VSS.n2112 VSS.n2035 0.1805
R36358 VSS.n2113 VSS.n2112 0.1805
R36359 VSS.n2047 VSS.n2046 0.1805
R36360 VSS.n2046 VSS.n2032 0.1805
R36361 VSS.n2094 VSS.n2042 0.1805
R36362 VSS.n2042 VSS.n2035 0.1805
R36363 VSS.n2092 VSS.n2043 0.1805
R36364 VSS.n2047 VSS.n2043 0.1805
R36365 VSS.n2093 VSS.n2044 0.1805
R36366 VSS.n2094 VSS.n2093 0.1805
R36367 VSS.n2091 VSS.n2051 0.1805
R36368 VSS.n2092 VSS.n2091 0.1805
R36369 VSS.n2086 VSS.n2054 0.1805
R36370 VSS.n2054 VSS.n2044 0.1805
R36371 VSS.n2087 VSS.n2053 0.1805
R36372 VSS.n2087 VSS.n2051 0.1805
R36373 VSS.n2085 VSS.n2056 0.1805
R36374 VSS.n2086 VSS.n2085 0.1805
R36375 VSS.n2072 VSS.n2061 0.1805
R36376 VSS.n2061 VSS.n2053 0.1805
R36377 VSS.n2073 VSS.n2060 0.1805
R36378 VSS.n2073 VSS.n2056 0.1805
R36379 VSS.n2071 VSS.n2067 0.1805
R36380 VSS.n2072 VSS.n2071 0.1805
R36381 VSS.n2066 VSS.n1634 0.1805
R36382 VSS.n2066 VSS.n2060 0.1805
R36383 VSS.n2230 VSS.n1635 0.1805
R36384 VSS.n2067 VSS.n1635 0.1805
R36385 VSS.n2231 VSS.n1633 0.1805
R36386 VSS.n2231 VSS.n1634 0.1805
R36387 VSS.n2230 VSS.n2229 0.1805
R36388 VSS.n1802 VSS.n1789 0.1805
R36389 VSS.n1804 VSS.n1787 0.1805
R36390 VSS.n1805 VSS.n1786 0.1805
R36391 VSS.n1806 VSS.n1785 0.1805
R36392 VSS.n1807 VSS.n1784 0.1805
R36393 VSS.n1808 VSS.n1783 0.1805
R36394 VSS.n1803 VSS.n1788 0.1805
R36395 VSS.n1803 VSS.n1664 0.1805
R36396 VSS.n1802 VSS.n1801 0.1805
R36397 VSS.n1801 VSS.n1662 0.1805
R36398 VSS.n1819 VSS.n1681 0.1805
R36399 VSS.n1827 VSS.n1681 0.1805
R36400 VSS.n1829 VSS.n1828 0.1805
R36401 VSS.n1828 VSS.n1682 0.1805
R36402 VSS.n1827 VSS.n1826 0.1805
R36403 VSS.n1826 VSS.n1684 0.1805
R36404 VSS.n1720 VSS.n1682 0.1805
R36405 VSS.n1721 VSS.n1720 0.1805
R36406 VSS.n1722 VSS.n1684 0.1805
R36407 VSS.n1728 VSS.n1722 0.1805
R36408 VSS.n1729 VSS.n1721 0.1805
R36409 VSS.n1729 VSS.n1716 0.1805
R36410 VSS.n1728 VSS.n1715 0.1805
R36411 VSS.n1734 VSS.n1715 0.1805
R36412 VSS.n1733 VSS.n1716 0.1805
R36413 VSS.n1733 VSS.n1710 0.1805
R36414 VSS.n1734 VSS.n1711 0.1805
R36415 VSS.n1741 VSS.n1711 0.1805
R36416 VSS.n1742 VSS.n1710 0.1805
R36417 VSS.n1742 VSS.n1707 0.1805
R36418 VSS.n1741 VSS.n1706 0.1805
R36419 VSS.n1749 VSS.n1706 0.1805
R36420 VSS.n1748 VSS.n1707 0.1805
R36421 VSS.n1748 VSS.n1708 0.1805
R36422 VSS.n1749 VSS.n805 0.1805
R36423 VSS.n3488 VSS.n805 0.1805
R36424 VSS.n1708 VSS.n806 0.1805
R36425 VSS.n3486 VSS.n806 0.1805
R36426 VSS.n3490 VSS.n802 0.1805
R36427 VSS.n3488 VSS.n3487 0.1805
R36428 VSS.n3487 VSS.n807 0.1805
R36429 VSS.n3486 VSS.n3485 0.1805
R36430 VSS.n3485 VSS.n809 0.1805
R36431 VSS.n812 VSS.n807 0.1805
R36432 VSS.n3480 VSS.n812 0.1805
R36433 VSS.n3481 VSS.n809 0.1805
R36434 VSS.n3481 VSS.n811 0.1805
R36435 VSS.n3480 VSS.n3479 0.1805
R36436 VSS.n3479 VSS.n814 0.1805
R36437 VSS.n737 VSS.n717 0.1805
R36438 VSS.n739 VSS.n738 0.1805
R36439 VSS.n3870 VSS.n715 0.1805
R36440 VSS.n3873 VSS.n714 0.1805
R36441 VSS.n3872 VSS.n3871 0.1805
R36442 VSS.n3871 VSS.n716 0.1805
R36443 VSS.n3870 VSS.n3869 0.1805
R36444 VSS.n3869 VSS.n3550 0.1805
R36445 VSS.n3553 VSS.n716 0.1805
R36446 VSS.n3864 VSS.n3553 0.1805
R36447 VSS.n3865 VSS.n3550 0.1805
R36448 VSS.n3865 VSS.n3552 0.1805
R36449 VSS.n3864 VSS.n3863 0.1805
R36450 VSS.n3863 VSS.n3555 0.1805
R36451 VSS.n3812 VSS.n3552 0.1805
R36452 VSS.n3813 VSS.n3812 0.1805
R36453 VSS.n3808 VSS.n3555 0.1805
R36454 VSS.n3848 VSS.n3808 0.1805
R36455 VSS.n3813 VSS.n3809 0.1805
R36456 VSS.n3846 VSS.n3809 0.1805
R36457 VSS.n3848 VSS.n3847 0.1805
R36458 VSS.n3847 VSS.n3810 0.1805
R36459 VSS.n3846 VSS.n3845 0.1805
R36460 VSS.n3845 VSS.n3817 0.1805
R36461 VSS.n3820 VSS.n3810 0.1805
R36462 VSS.n3840 VSS.n3820 0.1805
R36463 VSS.n3841 VSS.n3817 0.1805
R36464 VSS.n3841 VSS.n3819 0.1805
R36465 VSS.n3840 VSS.n3839 0.1805
R36466 VSS.n3839 VSS.n3827 0.1805
R36467 VSS.n3822 VSS.n3819 0.1805
R36468 VSS.n3825 VSS.n3822 0.1805
R36469 VSS.n3827 VSS.n3826 0.1805
R36470 VSS.n3826 VSS.n602 0.1805
R36471 VSS.n3825 VSS.n601 0.1805
R36472 VSS.n4038 VSS.n601 0.1805
R36473 VSS.n4037 VSS.n602 0.1805
R36474 VSS.n4037 VSS.n597 0.1805
R36475 VSS.n4038 VSS.n599 0.1805
R36476 VSS.n4042 VSS.n599 0.1805
R36477 VSS.n4075 VSS.n534 0.1805
R36478 VSS.n4043 VSS.n597 0.1805
R36479 VSS.n4043 VSS.n598 0.1805
R36480 VSS.n3953 VSS.n3881 0.1805
R36481 VSS.n3954 VSS.n3882 0.1805
R36482 VSS.n4007 VSS.n3882 0.1805
R36483 VSS.n4008 VSS.n3881 0.1805
R36484 VSS.n4008 VSS.n3879 0.1805
R36485 VSS.n4186 VSS.n449 0.1805
R36486 VSS.n3738 VSS.n449 0.1805
R36487 VSS.n3745 VSS.n3738 0.1805
R36488 VSS.n3745 VSS.n3731 0.1805
R36489 VSS.n3743 VSS.n3729 0.1805
R36490 VSS.n3749 VSS.n3731 0.1805
R36491 VSS.n3750 VSS.n3730 0.1805
R36492 VSS.n3749 VSS.n3732 0.1805
R36493 VSS.n3750 VSS.n3728 0.1805
R36494 VSS.n3734 VSS.n3732 0.1805
R36495 VSS.n3733 VSS.n3728 0.1805
R36496 VSS.n3734 VSS.n3723 0.1805
R36497 VSS.n3733 VSS.n3724 0.1805
R36498 VSS.n3759 VSS.n3723 0.1805
R36499 VSS.n3758 VSS.n3724 0.1805
R36500 VSS.n3759 VSS.n3721 0.1805
R36501 VSS.n3758 VSS.n3719 0.1805
R36502 VSS.n3756 VSS.n3715 0.1805
R36503 VSS.n3763 VSS.n3721 0.1805
R36504 VSS.n3764 VSS.n3719 0.1805
R36505 VSS.n3765 VSS.n3717 0.1805
R36506 VSS.n3766 VSS.n3715 0.1805
R36507 VSS.n3767 VSS.n3713 0.1805
R36508 VSS.n3768 VSS.n3711 0.1805
R36509 VSS.n3769 VSS.n3709 0.1805
R36510 VSS.n3770 VSS.n3707 0.1805
R36511 VSS.n3771 VSS.n3705 0.1805
R36512 VSS.n3772 VSS.n3703 0.1805
R36513 VSS.n3773 VSS.n3701 0.1805
R36514 VSS.n3774 VSS.n3699 0.1805
R36515 VSS.n3775 VSS.n3697 0.1805
R36516 VSS.n3776 VSS.n3696 0.1805
R36517 VSS.n3784 VSS.n3695 0.1805
R36518 VSS.n3783 VSS.n3777 0.1805
R36519 VSS.n3782 VSS.n3778 0.1805
R36520 VSS.n3783 VSS.n3567 0.1805
R36521 VSS.n3782 VSS.n3566 0.1805
R36522 VSS.n3788 VSS.n3567 0.1805
R36523 VSS.n3789 VSS.n3566 0.1805
R36524 VSS.n3788 VSS.n3568 0.1805
R36525 VSS.n3691 VSS.n3568 0.1805
R36526 VSS.n3691 VSS.n3570 0.1805
R36527 VSS.n3576 VSS.n3570 0.1805
R36528 VSS.n3688 VSS.n3572 0.1805
R36529 VSS.n3682 VSS.n3576 0.1805
R36530 VSS.n3683 VSS.n3571 0.1805
R36531 VSS.n3682 VSS.n3577 0.1805
R36532 VSS.n3683 VSS.n3575 0.1805
R36533 VSS.n3677 VSS.n3577 0.1805
R36534 VSS.n3676 VSS.n3575 0.1805
R36535 VSS.n3677 VSS.n3579 0.1805
R36536 VSS.n3676 VSS.n3580 0.1805
R36537 VSS.n3669 VSS.n3579 0.1805
R36538 VSS.n3670 VSS.n3580 0.1805
R36539 VSS.n3669 VSS.n3585 0.1805
R36540 VSS.n3670 VSS.n3584 0.1805
R36541 VSS.n3672 VSS.n3582 0.1805
R36542 VSS.n3665 VSS.n3585 0.1805
R36543 VSS.n3664 VSS.n3584 0.1805
R36544 VSS.n3663 VSS.n3583 0.1805
R36545 VSS.n3662 VSS.n3582 0.1805
R36546 VSS.n3661 VSS.n3591 0.1805
R36547 VSS.n3660 VSS.n3593 0.1805
R36548 VSS.n3659 VSS.n3595 0.1805
R36549 VSS.n3658 VSS.n3597 0.1805
R36550 VSS.n3657 VSS.n3599 0.1805
R36551 VSS.n3656 VSS.n3601 0.1805
R36552 VSS.n3655 VSS.n3603 0.1805
R36553 VSS.n3654 VSS.n3605 0.1805
R36554 VSS.n3653 VSS.n3607 0.1805
R36555 VSS.n3652 VSS.n3609 0.1805
R36556 VSS.n3651 VSS.n3611 0.1805
R36557 VSS.n3650 VSS.n3613 0.1805
R36558 VSS.n3649 VSS.n3615 0.1805
R36559 VSS.n3648 VSS.n3617 0.1805
R36560 VSS.n3647 VSS.n3619 0.1805
R36561 VSS.n3665 VSS.n3587 0.1805
R36562 VSS.n3664 VSS.n3588 0.1805
R36563 VSS.n3663 VSS.n3589 0.1805
R36564 VSS.n3662 VSS.n3590 0.1805
R36565 VSS.n3661 VSS.n3592 0.1805
R36566 VSS.n3660 VSS.n3594 0.1805
R36567 VSS.n3659 VSS.n3596 0.1805
R36568 VSS.n3658 VSS.n3598 0.1805
R36569 VSS.n3657 VSS.n3600 0.1805
R36570 VSS.n3656 VSS.n3602 0.1805
R36571 VSS.n3655 VSS.n3604 0.1805
R36572 VSS.n3654 VSS.n3606 0.1805
R36573 VSS.n3653 VSS.n3608 0.1805
R36574 VSS.n3652 VSS.n3610 0.1805
R36575 VSS.n3651 VSS.n3612 0.1805
R36576 VSS.n3650 VSS.n3614 0.1805
R36577 VSS.n3649 VSS.n3616 0.1805
R36578 VSS.n3648 VSS.n3618 0.1805
R36579 VSS.n3647 VSS.n3620 0.1805
R36580 VSS.n3642 VSS.n3621 0.1805
R36581 VSS.n3641 VSS.n3620 0.1805
R36582 VSS.n3640 VSS.n3618 0.1805
R36583 VSS.n3639 VSS.n3616 0.1805
R36584 VSS.n3638 VSS.n3614 0.1805
R36585 VSS.n3637 VSS.n3612 0.1805
R36586 VSS.n3636 VSS.n3610 0.1805
R36587 VSS.n3635 VSS.n3608 0.1805
R36588 VSS.n3634 VSS.n3606 0.1805
R36589 VSS.n3633 VSS.n3604 0.1805
R36590 VSS.n3632 VSS.n3602 0.1805
R36591 VSS.n3631 VSS.n3600 0.1805
R36592 VSS.n3630 VSS.n3598 0.1805
R36593 VSS.n3629 VSS.n3596 0.1805
R36594 VSS.n3628 VSS.n3594 0.1805
R36595 VSS.n3627 VSS.n3592 0.1805
R36596 VSS.n3626 VSS.n3590 0.1805
R36597 VSS.n3625 VSS.n3589 0.1805
R36598 VSS.n3624 VSS.n3588 0.1805
R36599 VSS.n3785 VSS.n3784 0.1805
R36600 VSS.n3776 VSS.n3694 0.1805
R36601 VSS.n3775 VSS.n3698 0.1805
R36602 VSS.n3774 VSS.n3700 0.1805
R36603 VSS.n3773 VSS.n3702 0.1805
R36604 VSS.n3772 VSS.n3704 0.1805
R36605 VSS.n3771 VSS.n3706 0.1805
R36606 VSS.n3770 VSS.n3708 0.1805
R36607 VSS.n3769 VSS.n3710 0.1805
R36608 VSS.n3768 VSS.n3712 0.1805
R36609 VSS.n3767 VSS.n3714 0.1805
R36610 VSS.n3766 VSS.n3716 0.1805
R36611 VSS.n3765 VSS.n3718 0.1805
R36612 VSS.n3764 VSS.n3720 0.1805
R36613 VSS.n4186 VSS.n450 0.1805
R36614 VSS.n4185 VSS.n451 0.1805
R36615 VSS.n4183 VSS.n455 0.1805
R36616 VSS.n1248 VSS.n1247 0.1805
R36617 VSS.n1249 VSS.n451 0.1805
R36618 VSS.n1249 VSS.n1244 0.1805
R36619 VSS.n1250 VSS.n454 0.1805
R36620 VSS.n1250 VSS.n1245 0.1805
R36621 VSS.n1251 VSS.n455 0.1805
R36622 VSS.n1252 VSS.n1251 0.1805
R36623 VSS.n1257 VSS.n1256 0.1805
R36624 VSS.n1255 VSS.n1244 0.1805
R36625 VSS.n1255 VSS.n1241 0.1805
R36626 VSS.n1254 VSS.n1245 0.1805
R36627 VSS.n1254 VSS.n1239 0.1805
R36628 VSS.n1253 VSS.n1252 0.1805
R36629 VSS.n1253 VSS.n1237 0.1805
R36630 VSS.n1297 VSS.n1296 0.1805
R36631 VSS.n1298 VSS.n1241 0.1805
R36632 VSS.n1298 VSS.n1242 0.1805
R36633 VSS.n1299 VSS.n1239 0.1805
R36634 VSS.n1299 VSS.n1240 0.1805
R36635 VSS.n1300 VSS.n1237 0.1805
R36636 VSS.n1300 VSS.n1238 0.1805
R36637 VSS.n1302 VSS.n1235 0.1805
R36638 VSS.n1303 VSS.n1234 0.1805
R36639 VSS.n1304 VSS.n1233 0.1805
R36640 VSS.n1305 VSS.n1232 0.1805
R36641 VSS.n1306 VSS.n1231 0.1805
R36642 VSS.n1307 VSS.n1230 0.1805
R36643 VSS.n1308 VSS.n1229 0.1805
R36644 VSS.n1309 VSS.n1228 0.1805
R36645 VSS.n1310 VSS.n1227 0.1805
R36646 VSS.n1311 VSS.n1226 0.1805
R36647 VSS.n1312 VSS.n1225 0.1805
R36648 VSS.n1313 VSS.n1224 0.1805
R36649 VSS.n1314 VSS.n1223 0.1805
R36650 VSS.n1315 VSS.n1222 0.1805
R36651 VSS.n1316 VSS.n1221 0.1805
R36652 VSS.n1317 VSS.n1220 0.1805
R36653 VSS.n1318 VSS.n1219 0.1805
R36654 VSS.n1319 VSS.n1218 0.1805
R36655 VSS.n1320 VSS.n1217 0.1805
R36656 VSS.n1321 VSS.n1216 0.1805
R36657 VSS.n1322 VSS.n1215 0.1805
R36658 VSS.n1323 VSS.n1214 0.1805
R36659 VSS.n1324 VSS.n1213 0.1805
R36660 VSS.n1325 VSS.n1212 0.1805
R36661 VSS.n1326 VSS.n1211 0.1805
R36662 VSS.n1327 VSS.n1210 0.1805
R36663 VSS.n1328 VSS.n1209 0.1805
R36664 VSS.n1329 VSS.n1208 0.1805
R36665 VSS.n1330 VSS.n1207 0.1805
R36666 VSS.n1331 VSS.n1206 0.1805
R36667 VSS.n1332 VSS.n1171 0.1805
R36668 VSS.n1333 VSS.n1169 0.1805
R36669 VSS.n1334 VSS.n1168 0.1805
R36670 VSS.n1301 VSS.n1236 0.1805
R36671 VSS.n3340 VSS.n1104 0.1805
R36672 VSS.n3341 VSS.n1102 0.1805
R36673 VSS.n3342 VSS.n1100 0.1805
R36674 VSS.n3343 VSS.n1098 0.1805
R36675 VSS.n3344 VSS.n1096 0.1805
R36676 VSS.n3345 VSS.n1094 0.1805
R36677 VSS.n3346 VSS.n1092 0.1805
R36678 VSS.n3347 VSS.n1090 0.1805
R36679 VSS.n3348 VSS.n1088 0.1805
R36680 VSS.n3349 VSS.n1086 0.1805
R36681 VSS.n3350 VSS.n1084 0.1805
R36682 VSS.n3351 VSS.n1082 0.1805
R36683 VSS.n3352 VSS.n1080 0.1805
R36684 VSS.n3353 VSS.n1078 0.1805
R36685 VSS.n3354 VSS.n1076 0.1805
R36686 VSS.n3355 VSS.n1074 0.1805
R36687 VSS.n3356 VSS.n1072 0.1805
R36688 VSS.n3357 VSS.n1070 0.1805
R36689 VSS.n3358 VSS.n1068 0.1805
R36690 VSS.n3359 VSS.n1066 0.1805
R36691 VSS.n3360 VSS.n1064 0.1805
R36692 VSS.n3361 VSS.n1062 0.1805
R36693 VSS.n3362 VSS.n1060 0.1805
R36694 VSS.n3363 VSS.n1058 0.1805
R36695 VSS.n3364 VSS.n1056 0.1805
R36696 VSS.n3365 VSS.n1054 0.1805
R36697 VSS.n3366 VSS.n1052 0.1805
R36698 VSS.n3367 VSS.n1050 0.1805
R36699 VSS.n3368 VSS.n1049 0.1805
R36700 VSS.n3339 VSS.n3338 0.1805
R36701 VSS.n3340 VSS.n1105 0.1805
R36702 VSS.n3341 VSS.n1103 0.1805
R36703 VSS.n3342 VSS.n1101 0.1805
R36704 VSS.n3343 VSS.n1099 0.1805
R36705 VSS.n3344 VSS.n1097 0.1805
R36706 VSS.n3345 VSS.n1095 0.1805
R36707 VSS.n3346 VSS.n1093 0.1805
R36708 VSS.n3347 VSS.n1091 0.1805
R36709 VSS.n3348 VSS.n1089 0.1805
R36710 VSS.n3349 VSS.n1087 0.1805
R36711 VSS.n3350 VSS.n1085 0.1805
R36712 VSS.n3351 VSS.n1083 0.1805
R36713 VSS.n3352 VSS.n1081 0.1805
R36714 VSS.n3353 VSS.n1079 0.1805
R36715 VSS.n3354 VSS.n1077 0.1805
R36716 VSS.n3355 VSS.n1075 0.1805
R36717 VSS.n3356 VSS.n1073 0.1805
R36718 VSS.n3357 VSS.n1071 0.1805
R36719 VSS.n3358 VSS.n1069 0.1805
R36720 VSS.n3359 VSS.n1067 0.1805
R36721 VSS.n3360 VSS.n1065 0.1805
R36722 VSS.n3361 VSS.n1063 0.1805
R36723 VSS.n3362 VSS.n1061 0.1805
R36724 VSS.n3363 VSS.n1059 0.1805
R36725 VSS.n3364 VSS.n1057 0.1805
R36726 VSS.n3365 VSS.n1055 0.1805
R36727 VSS.n3366 VSS.n1053 0.1805
R36728 VSS.n3367 VSS.n1051 0.1805
R36729 VSS.n3368 VSS.n1047 0.1805
R36730 VSS.n3338 VSS.n1107 0.1805
R36731 VSS.n3238 VSS.n1105 0.1805
R36732 VSS.n3239 VSS.n1103 0.1805
R36733 VSS.n3240 VSS.n1101 0.1805
R36734 VSS.n3241 VSS.n1099 0.1805
R36735 VSS.n3242 VSS.n1097 0.1805
R36736 VSS.n3243 VSS.n1095 0.1805
R36737 VSS.n3244 VSS.n1093 0.1805
R36738 VSS.n3245 VSS.n1091 0.1805
R36739 VSS.n3246 VSS.n1089 0.1805
R36740 VSS.n3248 VSS.n1087 0.1805
R36741 VSS.n3249 VSS.n1085 0.1805
R36742 VSS.n3250 VSS.n1083 0.1805
R36743 VSS.n3251 VSS.n1081 0.1805
R36744 VSS.n3252 VSS.n1079 0.1805
R36745 VSS.n3253 VSS.n1077 0.1805
R36746 VSS.n3254 VSS.n1075 0.1805
R36747 VSS.n3255 VSS.n1073 0.1805
R36748 VSS.n3256 VSS.n1071 0.1805
R36749 VSS.n3257 VSS.n1069 0.1805
R36750 VSS.n3258 VSS.n1067 0.1805
R36751 VSS.n3259 VSS.n1065 0.1805
R36752 VSS.n3260 VSS.n1063 0.1805
R36753 VSS.n3261 VSS.n1061 0.1805
R36754 VSS.n3262 VSS.n1059 0.1805
R36755 VSS.n3263 VSS.n1057 0.1805
R36756 VSS.n3264 VSS.n1055 0.1805
R36757 VSS.n3265 VSS.n1053 0.1805
R36758 VSS.n3266 VSS.n1051 0.1805
R36759 VSS.n3267 VSS.n1047 0.1805
R36760 VSS.n1108 VSS.n1107 0.1805
R36761 VSS.n3238 VSS.n3237 0.1805
R36762 VSS.n3239 VSS.n3235 0.1805
R36763 VSS.n3240 VSS.n3234 0.1805
R36764 VSS.n3241 VSS.n3233 0.1805
R36765 VSS.n3242 VSS.n3232 0.1805
R36766 VSS.n3243 VSS.n3230 0.1805
R36767 VSS.n3244 VSS.n3231 0.1805
R36768 VSS.n3289 VSS.n3245 0.1805
R36769 VSS.n3288 VSS.n3246 0.1805
R36770 VSS.n3287 VSS.n3248 0.1805
R36771 VSS.n3286 VSS.n3249 0.1805
R36772 VSS.n3285 VSS.n3250 0.1805
R36773 VSS.n3284 VSS.n3251 0.1805
R36774 VSS.n3283 VSS.n3252 0.1805
R36775 VSS.n3282 VSS.n3253 0.1805
R36776 VSS.n3281 VSS.n3254 0.1805
R36777 VSS.n3280 VSS.n3255 0.1805
R36778 VSS.n3279 VSS.n3256 0.1805
R36779 VSS.n3278 VSS.n3257 0.1805
R36780 VSS.n3277 VSS.n3258 0.1805
R36781 VSS.n3276 VSS.n3259 0.1805
R36782 VSS.n3275 VSS.n3260 0.1805
R36783 VSS.n3274 VSS.n3261 0.1805
R36784 VSS.n3273 VSS.n3262 0.1805
R36785 VSS.n3272 VSS.n3263 0.1805
R36786 VSS.n3271 VSS.n3264 0.1805
R36787 VSS.n3270 VSS.n3265 0.1805
R36788 VSS.n3269 VSS.n3266 0.1805
R36789 VSS.n3268 VSS.n3267 0.1805
R36790 VSS.n1109 VSS.n1108 0.1805
R36791 VSS.n3237 VSS.n3236 0.1805
R36792 VSS.n3235 VSS.n3226 0.1805
R36793 VSS.n3234 VSS.n3227 0.1805
R36794 VSS.n3233 VSS.n3228 0.1805
R36795 VSS.n3232 VSS.n3229 0.1805
R36796 VSS.n3292 VSS.n3230 0.1805
R36797 VSS.n3291 VSS.n3231 0.1805
R36798 VSS.n3290 VSS.n3289 0.1805
R36799 VSS.n3288 VSS.n3247 0.1805
R36800 VSS.n3287 VSS.n1017 0.1805
R36801 VSS.n3286 VSS.n1018 0.1805
R36802 VSS.n3285 VSS.n1019 0.1805
R36803 VSS.n3284 VSS.n1020 0.1805
R36804 VSS.n3283 VSS.n1021 0.1805
R36805 VSS.n3282 VSS.n1022 0.1805
R36806 VSS.n3281 VSS.n1023 0.1805
R36807 VSS.n3280 VSS.n1024 0.1805
R36808 VSS.n3279 VSS.n1025 0.1805
R36809 VSS.n3278 VSS.n1026 0.1805
R36810 VSS.n3277 VSS.n1027 0.1805
R36811 VSS.n3276 VSS.n1028 0.1805
R36812 VSS.n3275 VSS.n1029 0.1805
R36813 VSS.n3274 VSS.n1031 0.1805
R36814 VSS.n3273 VSS.n1032 0.1805
R36815 VSS.n3272 VSS.n1033 0.1805
R36816 VSS.n3271 VSS.n1034 0.1805
R36817 VSS.n3270 VSS.n1035 0.1805
R36818 VSS.n3269 VSS.n1036 0.1805
R36819 VSS.n3268 VSS.n1037 0.1805
R36820 VSS.n1110 VSS.n1109 0.1805
R36821 VSS.n3236 VSS.n3225 0.1805
R36822 VSS.n1111 VSS.n1110 0.1805
R36823 VSS.n1112 VSS.n1111 0.1805
R36824 VSS.n1113 VSS.n1112 0.1805
R36825 VSS.n1114 VSS.n1113 0.1805
R36826 VSS.n1115 VSS.n1114 0.1805
R36827 VSS.n1116 VSS.n1115 0.1805
R36828 VSS.n1117 VSS.n1116 0.1805
R36829 VSS.n1118 VSS.n1117 0.1805
R36830 VSS.n1119 VSS.n1118 0.1805
R36831 VSS.n1120 VSS.n1119 0.1805
R36832 VSS.n1121 VSS.n1120 0.1805
R36833 VSS.n1122 VSS.n1121 0.1805
R36834 VSS.n1123 VSS.n1122 0.1805
R36835 VSS.n3317 VSS.n1123 0.1805
R36836 VSS.n1149 VSS.n1138 0.1805
R36837 VSS.n1148 VSS.n1137 0.1805
R36838 VSS.n1147 VSS.n1136 0.1805
R36839 VSS.n1146 VSS.n1135 0.1805
R36840 VSS.n1145 VSS.n1134 0.1805
R36841 VSS.n1144 VSS.n1133 0.1805
R36842 VSS.n1143 VSS.n1132 0.1805
R36843 VSS.n1142 VSS.n1131 0.1805
R36844 VSS.n1141 VSS.n1130 0.1805
R36845 VSS.n1140 VSS.n1129 0.1805
R36846 VSS.n1128 VSS.n1124 0.1805
R36847 VSS.n3318 VSS.n1125 0.1805
R36848 VSS.n3317 VSS.n1126 0.1805
R36849 VSS.n1360 VSS.n1135 0.1805
R36850 VSS.n1359 VSS.n1136 0.1805
R36851 VSS.n1358 VSS.n1137 0.1805
R36852 VSS.n1357 VSS.n1138 0.1805
R36853 VSS.n1356 VSS.n1139 0.1805
R36854 VSS.n1182 VSS.n1178 0.1805
R36855 VSS.n1186 VSS.n1178 0.1805
R36856 VSS.n1187 VSS.n1186 0.1805
R36857 VSS.n1188 VSS.n1187 0.1805
R36858 VSS.n1188 VSS.n1176 0.1805
R36859 VSS.n1192 VSS.n1176 0.1805
R36860 VSS.n1193 VSS.n1192 0.1805
R36861 VSS.n1194 VSS.n1193 0.1805
R36862 VSS.n1194 VSS.n1174 0.1805
R36863 VSS.n1198 VSS.n1174 0.1805
R36864 VSS.n1199 VSS.n1198 0.1805
R36865 VSS.n1200 VSS.n1199 0.1805
R36866 VSS.n1200 VSS.n1172 0.1805
R36867 VSS.n1204 VSS.n1172 0.1805
R36868 VSS.n1333 VSS.n1170 0.1805
R36869 VSS.n1205 VSS.n1204 0.1805
R36870 VSS.n1332 VSS.n1205 0.1805
R36871 VSS.n1166 VSS.n1165 0.1805
R36872 VSS.n1334 VSS.n1166 0.1805
R36873 VSS.n1203 VSS.n1202 0.1805
R36874 VSS.n1203 VSS.n1170 0.1805
R36875 VSS.n1164 VSS.n1163 0.1805
R36876 VSS.n1165 VSS.n1164 0.1805
R36877 VSS.n1201 VSS.n1173 0.1805
R36878 VSS.n1202 VSS.n1201 0.1805
R36879 VSS.n1162 VSS.n1161 0.1805
R36880 VSS.n1163 VSS.n1162 0.1805
R36881 VSS.n1197 VSS.n1196 0.1805
R36882 VSS.n1197 VSS.n1173 0.1805
R36883 VSS.n1160 VSS.n1159 0.1805
R36884 VSS.n1161 VSS.n1160 0.1805
R36885 VSS.n1195 VSS.n1175 0.1805
R36886 VSS.n1196 VSS.n1195 0.1805
R36887 VSS.n1158 VSS.n1157 0.1805
R36888 VSS.n1159 VSS.n1158 0.1805
R36889 VSS.n1191 VSS.n1190 0.1805
R36890 VSS.n1191 VSS.n1175 0.1805
R36891 VSS.n1156 VSS.n1155 0.1805
R36892 VSS.n1157 VSS.n1156 0.1805
R36893 VSS.n1189 VSS.n1177 0.1805
R36894 VSS.n1190 VSS.n1189 0.1805
R36895 VSS.n1154 VSS.n1153 0.1805
R36896 VSS.n1155 VSS.n1154 0.1805
R36897 VSS.n1185 VSS.n1184 0.1805
R36898 VSS.n1185 VSS.n1177 0.1805
R36899 VSS.n1152 VSS.n1151 0.1805
R36900 VSS.n1153 VSS.n1152 0.1805
R36901 VSS.n1183 VSS.n1179 0.1805
R36902 VSS.n1184 VSS.n1183 0.1805
R36903 VSS.n1180 VSS.n1150 0.1805
R36904 VSS.n1151 VSS.n1150 0.1805
R36905 VSS.n1355 VSS.n1354 0.1805
R36906 VSS.n3212 VSS.n1372 0.1805
R36907 VSS.n3207 VSS.n1373 0.1805
R36908 VSS.n3211 VSS.n1373 0.1805
R36909 VSS.n3210 VSS.n1374 0.1805
R36910 VSS.n3215 VSS.n3214 0.1805
R36911 VSS.n1369 VSS.n1126 0.1805
R36912 VSS.n1368 VSS.n1125 0.1805
R36913 VSS.n1367 VSS.n1128 0.1805
R36914 VSS.n1366 VSS.n1129 0.1805
R36915 VSS.n1365 VSS.n1130 0.1805
R36916 VSS.n1364 VSS.n1131 0.1805
R36917 VSS.n1363 VSS.n1132 0.1805
R36918 VSS.n1362 VSS.n1133 0.1805
R36919 VSS.n1361 VSS.n1134 0.1805
R36920 VSS.n1370 VSS.n1127 0.1805
R36921 VSS.n3316 VSS.n1127 0.1805
R36922 VSS.n3216 VSS.n3215 0.1805
R36923 VSS.n3314 VSS.n3216 0.1805
R36924 VSS.n3316 VSS.n3315 0.1805
R36925 VSS.n3315 VSS.n3217 0.1805
R36926 VSS.n3314 VSS.n3313 0.1805
R36927 VSS.n3313 VSS.n3312 0.1805
R36928 VSS.n3218 VSS.n3217 0.1805
R36929 VSS.n3310 VSS.n3218 0.1805
R36930 VSS.n3312 VSS.n3311 0.1805
R36931 VSS.n3311 VSS.n3219 0.1805
R36932 VSS.n3310 VSS.n3309 0.1805
R36933 VSS.n3309 VSS.n3308 0.1805
R36934 VSS.n3220 VSS.n3219 0.1805
R36935 VSS.n3306 VSS.n3220 0.1805
R36936 VSS.n3308 VSS.n3307 0.1805
R36937 VSS.n3307 VSS.n3221 0.1805
R36938 VSS.n3306 VSS.n3305 0.1805
R36939 VSS.n3305 VSS.n3304 0.1805
R36940 VSS.n3222 VSS.n3221 0.1805
R36941 VSS.n3302 VSS.n3222 0.1805
R36942 VSS.n3304 VSS.n3303 0.1805
R36943 VSS.n3303 VSS.n3223 0.1805
R36944 VSS.n3302 VSS.n3301 0.1805
R36945 VSS.n3301 VSS.n3300 0.1805
R36946 VSS.n3224 VSS.n3223 0.1805
R36947 VSS.n3298 VSS.n3224 0.1805
R36948 VSS.n3300 VSS.n3299 0.1805
R36949 VSS.n3299 VSS.n3225 0.1805
R36950 VSS.n3298 VSS.n3297 0.1805
R36951 VSS.n3297 VSS.n3226 0.1805
R36952 VSS.n3296 VSS.n3227 0.1805
R36953 VSS.n3295 VSS.n3228 0.1805
R36954 VSS.n3294 VSS.n3229 0.1805
R36955 VSS.n3293 VSS.n3292 0.1805
R36956 VSS.n3291 VSS.n1015 0.1805
R36957 VSS.n3399 VSS.n1017 0.1805
R36958 VSS.n3398 VSS.n1018 0.1805
R36959 VSS.n3397 VSS.n1019 0.1805
R36960 VSS.n3396 VSS.n1020 0.1805
R36961 VSS.n3395 VSS.n1021 0.1805
R36962 VSS.n3394 VSS.n1022 0.1805
R36963 VSS.n3393 VSS.n1023 0.1805
R36964 VSS.n3392 VSS.n1024 0.1805
R36965 VSS.n3391 VSS.n1025 0.1805
R36966 VSS.n3390 VSS.n1026 0.1805
R36967 VSS.n3389 VSS.n1027 0.1805
R36968 VSS.n3385 VSS.n1031 0.1805
R36969 VSS.n3387 VSS.n1029 0.1805
R36970 VSS.n3388 VSS.n1028 0.1805
R36971 VSS.n3384 VSS.n1032 0.1805
R36972 VSS.n3383 VSS.n1033 0.1805
R36973 VSS.n3382 VSS.n1034 0.1805
R36974 VSS.n3381 VSS.n1035 0.1805
R36975 VSS.n3379 VSS.n1037 0.1805
R36976 VSS.n3379 VSS.n1038 0.1805
R36977 VSS.n3138 VSS.n1038 0.1805
R36978 VSS.n3150 VSS.n3138 0.1805
R36979 VSS.n3151 VSS.n3150 0.1805
R36980 VSS.n3152 VSS.n3151 0.1805
R36981 VSS.n3152 VSS.n3136 0.1805
R36982 VSS.n3136 VSS.n3135 0.1805
R36983 VSS.n3135 VSS.n3125 0.1805
R36984 VSS.n3162 VSS.n3125 0.1805
R36985 VSS.n3163 VSS.n3162 0.1805
R36986 VSS.n3164 VSS.n3163 0.1805
R36987 VSS.n3164 VSS.n3123 0.1805
R36988 VSS.n3168 VSS.n1380 0.1805
R36989 VSS.n3169 VSS.n1382 0.1805
R36990 VSS.n3171 VSS.n1384 0.1805
R36991 VSS.n3172 VSS.n1386 0.1805
R36992 VSS.n3173 VSS.n1388 0.1805
R36993 VSS.n3174 VSS.n1390 0.1805
R36994 VSS.n3175 VSS.n1392 0.1805
R36995 VSS.n3176 VSS.n1394 0.1805
R36996 VSS.n3177 VSS.n1396 0.1805
R36997 VSS.n3178 VSS.n1398 0.1805
R36998 VSS.n3179 VSS.n1400 0.1805
R36999 VSS.n3181 VSS.n1402 0.1805
R37000 VSS.n3075 VSS.n1444 0.1805
R37001 VSS.n3074 VSS.n1446 0.1805
R37002 VSS.n3073 VSS.n1448 0.1805
R37003 VSS.n3072 VSS.n1450 0.1805
R37004 VSS.n3071 VSS.n1452 0.1805
R37005 VSS.n3070 VSS.n1454 0.1805
R37006 VSS.n3069 VSS.n1456 0.1805
R37007 VSS.n3068 VSS.n1458 0.1805
R37008 VSS.n3067 VSS.n1460 0.1805
R37009 VSS.n3066 VSS.n1462 0.1805
R37010 VSS.n3065 VSS.n1464 0.1805
R37011 VSS.n3064 VSS.n1466 0.1805
R37012 VSS.n3063 VSS.n1468 0.1805
R37013 VSS.n3062 VSS.n1470 0.1805
R37014 VSS.n3061 VSS.n1472 0.1805
R37015 VSS.n3060 VSS.n1474 0.1805
R37016 VSS.n3059 VSS.n1476 0.1805
R37017 VSS.n3076 VSS.n1443 0.1805
R37018 VSS.n3075 VSS.n1445 0.1805
R37019 VSS.n3074 VSS.n1447 0.1805
R37020 VSS.n3073 VSS.n1449 0.1805
R37021 VSS.n3072 VSS.n1451 0.1805
R37022 VSS.n3071 VSS.n1453 0.1805
R37023 VSS.n3070 VSS.n1455 0.1805
R37024 VSS.n3069 VSS.n1457 0.1805
R37025 VSS.n3068 VSS.n1459 0.1805
R37026 VSS.n3067 VSS.n1461 0.1805
R37027 VSS.n3066 VSS.n1463 0.1805
R37028 VSS.n3065 VSS.n1465 0.1805
R37029 VSS.n3064 VSS.n1467 0.1805
R37030 VSS.n3063 VSS.n1469 0.1805
R37031 VSS.n3062 VSS.n1471 0.1805
R37032 VSS.n3061 VSS.n1473 0.1805
R37033 VSS.n3060 VSS.n1475 0.1805
R37034 VSS.n3059 VSS.n1477 0.1805
R37035 VSS.n1443 VSS.n1442 0.1805
R37036 VSS.n1529 VSS.n1445 0.1805
R37037 VSS.n1530 VSS.n1447 0.1805
R37038 VSS.n1442 VSS.n1441 0.1805
R37039 VSS.n1529 VSS.n1528 0.1805
R37040 VSS.n1441 VSS.n1438 0.1805
R37041 VSS.n1528 VSS.n1437 0.1805
R37042 VSS.n3087 VSS.n1434 0.1805
R37043 VSS.n3083 VSS.n1438 0.1805
R37044 VSS.n3084 VSS.n1437 0.1805
R37045 VSS.n3086 VSS.n1431 0.1805
R37046 VSS.n1439 VSS.n1429 0.1805
R37047 VSS.n3083 VSS.n1439 0.1805
R37048 VSS.n1435 VSS.n1430 0.1805
R37049 VSS.n3084 VSS.n1435 0.1805
R37050 VSS.n3086 VSS.n3085 0.1805
R37051 VSS.n3085 VSS.n1436 0.1805
R37052 VSS.n1525 VSS.n1434 0.1805
R37053 VSS.n1526 VSS.n1525 0.1805
R37054 VSS.n1527 VSS.n1436 0.1805
R37055 VSS.n1530 VSS.n1527 0.1805
R37056 VSS.n1531 VSS.n1526 0.1805
R37057 VSS.n1531 VSS.n1449 0.1805
R37058 VSS.n1533 VSS.n1453 0.1805
R37059 VSS.n1534 VSS.n1455 0.1805
R37060 VSS.n1535 VSS.n1457 0.1805
R37061 VSS.n1536 VSS.n1459 0.1805
R37062 VSS.n1537 VSS.n1461 0.1805
R37063 VSS.n1538 VSS.n1463 0.1805
R37064 VSS.n1539 VSS.n1465 0.1805
R37065 VSS.n1540 VSS.n1467 0.1805
R37066 VSS.n1541 VSS.n1469 0.1805
R37067 VSS.n1542 VSS.n1471 0.1805
R37068 VSS.n1543 VSS.n1473 0.1805
R37069 VSS.n1544 VSS.n1475 0.1805
R37070 VSS.n1545 VSS.n1477 0.1805
R37071 VSS.n1545 VSS.n1524 0.1805
R37072 VSS.n1553 VSS.n1524 0.1805
R37073 VSS.n1554 VSS.n1553 0.1805
R37074 VSS.n1555 VSS.n1554 0.1805
R37075 VSS.n1555 VSS.n1521 0.1805
R37076 VSS.n1559 VSS.n1521 0.1805
R37077 VSS.n1560 VSS.n1559 0.1805
R37078 VSS.n1561 VSS.n1560 0.1805
R37079 VSS.n1561 VSS.n1519 0.1805
R37080 VSS.n1565 VSS.n1519 0.1805
R37081 VSS.n1566 VSS.n1565 0.1805
R37082 VSS.n1567 VSS.n1566 0.1805
R37083 VSS.n1567 VSS.n1517 0.1805
R37084 VSS.n1571 VSS.n1517 0.1805
R37085 VSS.n1572 VSS.n1571 0.1805
R37086 VSS.n1573 VSS.n1572 0.1805
R37087 VSS.n1573 VSS.n1515 0.1805
R37088 VSS.n1577 VSS.n1515 0.1805
R37089 VSS.n1578 VSS.n1577 0.1805
R37090 VSS.n1579 VSS.n1578 0.1805
R37091 VSS.n1579 VSS.n1513 0.1805
R37092 VSS.n1583 VSS.n1513 0.1805
R37093 VSS.n1584 VSS.n1583 0.1805
R37094 VSS.n1585 VSS.n1584 0.1805
R37095 VSS.n1585 VSS.n1511 0.1805
R37096 VSS.n1589 VSS.n1511 0.1805
R37097 VSS.n1590 VSS.n1589 0.1805
R37098 VSS.n2258 VSS.n1590 0.1805
R37099 VSS.n2260 VSS.n1508 0.1805
R37100 VSS.n2245 VSS.n1603 0.1805
R37101 VSS.n1616 VSS.n1602 0.1805
R37102 VSS.n2246 VSS.n1602 0.1805
R37103 VSS.n1615 VSS.n1601 0.1805
R37104 VSS.n2247 VSS.n1601 0.1805
R37105 VSS.n1614 VSS.n1600 0.1805
R37106 VSS.n2248 VSS.n1600 0.1805
R37107 VSS.n1613 VSS.n1599 0.1805
R37108 VSS.n2249 VSS.n1599 0.1805
R37109 VSS.n1612 VSS.n1598 0.1805
R37110 VSS.n2250 VSS.n1598 0.1805
R37111 VSS.n1611 VSS.n1597 0.1805
R37112 VSS.n2251 VSS.n1597 0.1805
R37113 VSS.n1610 VSS.n1596 0.1805
R37114 VSS.n2252 VSS.n1596 0.1805
R37115 VSS.n1609 VSS.n1595 0.1805
R37116 VSS.n2253 VSS.n1595 0.1805
R37117 VSS.n1608 VSS.n1594 0.1805
R37118 VSS.n2254 VSS.n1594 0.1805
R37119 VSS.n1607 VSS.n1593 0.1805
R37120 VSS.n2255 VSS.n1593 0.1805
R37121 VSS.n1606 VSS.n1592 0.1805
R37122 VSS.n2256 VSS.n1592 0.1805
R37123 VSS.n1605 VSS.n1591 0.1805
R37124 VSS.n2257 VSS.n1591 0.1805
R37125 VSS.n1604 VSS.n1509 0.1805
R37126 VSS.n2258 VSS.n1509 0.1805
R37127 VSS.n2261 VSS.n1507 0.1805
R37128 VSS.n2260 VSS.n2259 0.1805
R37129 VSS.n2259 VSS.n1510 0.1805
R37130 VSS.n1507 VSS.n1506 0.1805
R37131 VSS.n1506 VSS.n1505 0.1805
R37132 VSS.n1588 VSS.n1510 0.1805
R37133 VSS.n1588 VSS.n1587 0.1805
R37134 VSS.n1505 VSS.n1504 0.1805
R37135 VSS.n1504 VSS.n1503 0.1805
R37136 VSS.n1587 VSS.n1586 0.1805
R37137 VSS.n1586 VSS.n1512 0.1805
R37138 VSS.n1503 VSS.n1502 0.1805
R37139 VSS.n1502 VSS.n1501 0.1805
R37140 VSS.n1582 VSS.n1512 0.1805
R37141 VSS.n1582 VSS.n1581 0.1805
R37142 VSS.n1501 VSS.n1500 0.1805
R37143 VSS.n1500 VSS.n1499 0.1805
R37144 VSS.n1581 VSS.n1580 0.1805
R37145 VSS.n1580 VSS.n1514 0.1805
R37146 VSS.n1499 VSS.n1498 0.1805
R37147 VSS.n1498 VSS.n1497 0.1805
R37148 VSS.n1576 VSS.n1514 0.1805
R37149 VSS.n1576 VSS.n1575 0.1805
R37150 VSS.n1497 VSS.n1496 0.1805
R37151 VSS.n1496 VSS.n1495 0.1805
R37152 VSS.n1575 VSS.n1574 0.1805
R37153 VSS.n1574 VSS.n1516 0.1805
R37154 VSS.n1495 VSS.n1494 0.1805
R37155 VSS.n1494 VSS.n1493 0.1805
R37156 VSS.n1570 VSS.n1516 0.1805
R37157 VSS.n1570 VSS.n1569 0.1805
R37158 VSS.n1493 VSS.n1492 0.1805
R37159 VSS.n1492 VSS.n1491 0.1805
R37160 VSS.n1569 VSS.n1568 0.1805
R37161 VSS.n1568 VSS.n1518 0.1805
R37162 VSS.n1491 VSS.n1490 0.1805
R37163 VSS.n1490 VSS.n1489 0.1805
R37164 VSS.n1564 VSS.n1518 0.1805
R37165 VSS.n1564 VSS.n1563 0.1805
R37166 VSS.n1489 VSS.n1488 0.1805
R37167 VSS.n1488 VSS.n1487 0.1805
R37168 VSS.n1563 VSS.n1562 0.1805
R37169 VSS.n1562 VSS.n1520 0.1805
R37170 VSS.n1487 VSS.n1486 0.1805
R37171 VSS.n1486 VSS.n1485 0.1805
R37172 VSS.n1558 VSS.n1520 0.1805
R37173 VSS.n1558 VSS.n1557 0.1805
R37174 VSS.n1485 VSS.n1484 0.1805
R37175 VSS.n1484 VSS.n1481 0.1805
R37176 VSS.n1557 VSS.n1556 0.1805
R37177 VSS.n1556 VSS.n1523 0.1805
R37178 VSS.n1522 VSS.n1481 0.1805
R37179 VSS.n1552 VSS.n1523 0.1805
R37180 VSS.n1552 VSS.n1549 0.1805
R37181 VSS.n1551 VSS.n1550 0.1805
R37182 VSS.n1549 VSS.n1548 0.1805
R37183 VSS.n1548 VSS.n1478 0.1805
R37184 VSS.n1532 VSS.n1451 0.1805
R37185 VSS.n1547 VSS.n1546 0.1805
R37186 VSS.n3058 VSS.n1478 0.1805
R37187 VSS.n3058 VSS.n1479 0.1805
R37188 VSS.n3057 VSS.n3056 0.1805
R37189 VSS.n3122 VSS.n1377 0.1805
R37190 VSS.n3123 VSS.n3122 0.1805
R37191 VSS.n3120 VSS.n1378 0.1805
R37192 VSS.n3166 VSS.n3120 0.1805
R37193 VSS.n3168 VSS.n3167 0.1805
R37194 VSS.n3167 VSS.n3121 0.1805
R37195 VSS.n3166 VSS.n3165 0.1805
R37196 VSS.n3165 VSS.n3124 0.1805
R37197 VSS.n3127 VSS.n3121 0.1805
R37198 VSS.n3160 VSS.n3127 0.1805
R37199 VSS.n3161 VSS.n3124 0.1805
R37200 VSS.n3161 VSS.n3126 0.1805
R37201 VSS.n3160 VSS.n3159 0.1805
R37202 VSS.n3159 VSS.n3131 0.1805
R37203 VSS.n3134 VSS.n3126 0.1805
R37204 VSS.n3154 VSS.n3134 0.1805
R37205 VSS.n3155 VSS.n3131 0.1805
R37206 VSS.n3155 VSS.n3133 0.1805
R37207 VSS.n3154 VSS.n3153 0.1805
R37208 VSS.n3153 VSS.n3137 0.1805
R37209 VSS.n3140 VSS.n3133 0.1805
R37210 VSS.n3148 VSS.n3140 0.1805
R37211 VSS.n3149 VSS.n3137 0.1805
R37212 VSS.n3149 VSS.n3139 0.1805
R37213 VSS.n3148 VSS.n3147 0.1805
R37214 VSS.n3147 VSS.n3143 0.1805
R37215 VSS.n3139 VSS.n1039 0.1805
R37216 VSS.n3378 VSS.n1039 0.1805
R37217 VSS.n3143 VSS.n1040 0.1805
R37218 VSS.n3376 VSS.n1040 0.1805
R37219 VSS.n3380 VSS.n1036 0.1805
R37220 VSS.n3378 VSS.n3377 0.1805
R37221 VSS.n3377 VSS.n1041 0.1805
R37222 VSS.n3376 VSS.n3375 0.1805
R37223 VSS.n3375 VSS.n1043 0.1805
R37224 VSS.n1046 VSS.n1041 0.1805
R37225 VSS.n3370 VSS.n1046 0.1805
R37226 VSS.n3371 VSS.n1043 0.1805
R37227 VSS.n3371 VSS.n1045 0.1805
R37228 VSS.n3370 VSS.n3369 0.1805
R37229 VSS.n3369 VSS.n1048 0.1805
R37230 VSS.n1294 VSS.n1242 0.1805
R37231 VSS.n1293 VSS.n1240 0.1805
R37232 VSS.n1292 VSS.n1238 0.1805
R37233 VSS.n1291 VSS.n1236 0.1805
R37234 VSS.n1290 VSS.n1235 0.1805
R37235 VSS.n1289 VSS.n1234 0.1805
R37236 VSS.n1288 VSS.n1233 0.1805
R37237 VSS.n1287 VSS.n1232 0.1805
R37238 VSS.n1286 VSS.n1231 0.1805
R37239 VSS.n1285 VSS.n1230 0.1805
R37240 VSS.n1284 VSS.n1229 0.1805
R37241 VSS.n1283 VSS.n1228 0.1805
R37242 VSS.n1282 VSS.n1227 0.1805
R37243 VSS.n1281 VSS.n1226 0.1805
R37244 VSS.n1280 VSS.n1225 0.1805
R37245 VSS.n1279 VSS.n1224 0.1805
R37246 VSS.n1278 VSS.n1223 0.1805
R37247 VSS.n1277 VSS.n1222 0.1805
R37248 VSS.n1276 VSS.n1221 0.1805
R37249 VSS.n1275 VSS.n1220 0.1805
R37250 VSS.n1274 VSS.n1219 0.1805
R37251 VSS.n1273 VSS.n1218 0.1805
R37252 VSS.n1272 VSS.n1217 0.1805
R37253 VSS.n1271 VSS.n1216 0.1805
R37254 VSS.n1270 VSS.n1215 0.1805
R37255 VSS.n1269 VSS.n1214 0.1805
R37256 VSS.n1268 VSS.n1213 0.1805
R37257 VSS.n1267 VSS.n1212 0.1805
R37258 VSS.n1266 VSS.n1211 0.1805
R37259 VSS.n1265 VSS.n1210 0.1805
R37260 VSS.n1264 VSS.n1209 0.1805
R37261 VSS.n1263 VSS.n1208 0.1805
R37262 VSS.n1262 VSS.n1207 0.1805
R37263 VSS.n1261 VSS.n1206 0.1805
R37264 VSS.n1260 VSS.n1171 0.1805
R37265 VSS.n1259 VSS.n1169 0.1805
R37266 VSS.n3645 VSS.n3623 0.1805
R37267 VSS.n3646 VSS.n3621 0.1805
R37268 VSS.n3646 VSS.n3622 0.1805
R37269 VSS.n3671 VSS.n3583 0.1805
R37270 VSS.n3671 VSS.n3581 0.1805
R37271 VSS.n3673 VSS.n3672 0.1805
R37272 VSS.n3674 VSS.n3673 0.1805
R37273 VSS.n3675 VSS.n3581 0.1805
R37274 VSS.n3675 VSS.n3574 0.1805
R37275 VSS.n3674 VSS.n3573 0.1805
R37276 VSS.n3685 VSS.n3573 0.1805
R37277 VSS.n3684 VSS.n3574 0.1805
R37278 VSS.n3684 VSS.n3572 0.1805
R37279 VSS.n3686 VSS.n3685 0.1805
R37280 VSS.n3689 VSS.n3571 0.1805
R37281 VSS.n3690 VSS.n3689 0.1805
R37282 VSS.n3688 VSS.n3563 0.1805
R37283 VSS.n3791 VSS.n3563 0.1805
R37284 VSS.n3690 VSS.n3564 0.1805
R37285 VSS.n3789 VSS.n3564 0.1805
R37286 VSS.n3791 VSS.n3790 0.1805
R37287 VSS.n3790 VSS.n3565 0.1805
R37288 VSS.n3779 VSS.n3562 0.1805
R37289 VSS.n3781 VSS.n3565 0.1805
R37290 VSS.n3757 VSS.n3717 0.1805
R37291 VSS.n3757 VSS.n3725 0.1805
R37292 VSS.n3756 VSS.n3755 0.1805
R37293 VSS.n3755 VSS.n3754 0.1805
R37294 VSS.n3726 VSS.n3725 0.1805
R37295 VSS.n3752 VSS.n3726 0.1805
R37296 VSS.n3754 VSS.n3753 0.1805
R37297 VSS.n3753 VSS.n3727 0.1805
R37298 VSS.n3752 VSS.n3751 0.1805
R37299 VSS.n3751 VSS.n3729 0.1805
R37300 VSS.n3740 VSS.n3727 0.1805
R37301 VSS.n3744 VSS.n3730 0.1805
R37302 VSS.n3744 VSS.n3739 0.1805
R37303 VSS.n3743 VSS.n3742 0.1805
R37304 VSS.n3742 VSS.n453 0.1805
R37305 VSS.n3739 VSS.n452 0.1805
R37306 VSS.n4185 VSS.n452 0.1805
R37307 VSS.n4184 VSS.n453 0.1805
R37308 VSS.n4184 VSS.n454 0.1805
R37309 VSS.n3088 VSS.n3087 0.1805
R37310 VSS.n3091 VSS.n1426 0.1805
R37311 VSS.n3091 VSS.n1430 0.1805
R37312 VSS.n3098 VSS.n1425 0.1805
R37313 VSS.n3090 VSS.n1425 0.1805
R37314 VSS.n3097 VSS.n1422 0.1805
R37315 VSS.n3097 VSS.n1426 0.1805
R37316 VSS.n3102 VSS.n1423 0.1805
R37317 VSS.n3098 VSS.n1423 0.1805
R37318 VSS.n3101 VSS.n1416 0.1805
R37319 VSS.n3101 VSS.n3100 0.1805
R37320 VSS.n3110 VSS.n1417 0.1805
R37321 VSS.n3102 VSS.n1417 0.1805
R37322 VSS.n3112 VSS.n3111 0.1805
R37323 VSS.n3111 VSS.n1416 0.1805
R37324 VSS.n3114 VSS.n1415 0.1805
R37325 VSS.n3110 VSS.n1415 0.1805
R37326 VSS.n3113 VSS.n1408 0.1805
R37327 VSS.n3113 VSS.n3112 0.1805
R37328 VSS.n3184 VSS.n1409 0.1805
R37329 VSS.n3114 VSS.n1409 0.1805
R37330 VSS.n3186 VSS.n3185 0.1805
R37331 VSS.n3185 VSS.n1408 0.1805
R37332 VSS.n3188 VSS.n1407 0.1805
R37333 VSS.n3184 VSS.n1407 0.1805
R37334 VSS.n1759 VSS.n1697 0.179316
R37335 VSS.n4014 VSS.n4013 0.17825
R37336 VSS.n4015 VSS.n3877 0.17825
R37337 VSS.n4017 VSS.n4016 0.17825
R37338 VSS.n4018 VSS.n711 0.17825
R37339 VSS.n4024 VSS.n712 0.17825
R37340 VSS.n4023 VSS.n4022 0.17825
R37341 VSS.n2003 VSS.n1945 0.17825
R37342 VSS.n2002 VSS.n2001 0.17825
R37343 VSS.n2000 VSS.n1996 0.17825
R37344 VSS.n2130 VSS.n2129 0.17825
R37345 VSS.n1999 VSS.n1998 0.17825
R37346 VSS.n2021 VSS.n2020 0.17825
R37347 VSS.n2023 VSS.n2022 0.17825
R37348 VSS.n2010 VSS.n2008 0.17825
R37349 VSS.n2123 VSS.n2122 0.17825
R37350 VSS.n2009 VSS.n2007 0.17825
R37351 VSS.n2102 VSS.n2101 0.17825
R37352 VSS.n2104 VSS.n2103 0.17825
R37353 VSS.n2105 VSS.n2034 0.17825
R37354 VSS.n2037 VSS.n2036 0.17825
R37355 VSS.n2041 VSS.n2039 0.17825
R37356 VSS.n2096 VSS.n2095 0.17825
R37357 VSS.n2040 VSS.n2038 0.17825
R37358 VSS.n2079 VSS.n2078 0.17825
R37359 VSS.n2081 VSS.n2080 0.17825
R37360 VSS.n2082 VSS.n2055 0.17825
R37361 VSS.n2084 VSS.n2083 0.17825
R37362 VSS.n2076 VSS.n2057 0.17825
R37363 VSS.n2075 VSS.n2074 0.17825
R37364 VSS.n2059 VSS.n2058 0.17825
R37365 VSS.n2065 VSS.n2064 0.17825
R37366 VSS.n3856 VSS.n714 0.17825
R37367 VSS.n3858 VSS.n3857 0.17825
R37368 VSS.n2064 VSS.n1630 0.178132
R37369 VSS.n2128 VSS.n2000 0.176947
R37370 VSS.n1915 VSS.n1867 0.176947
R37371 VSS.n3504 VSS.n3503 0.175763
R37372 VSS.n1295 VSS.n1294 0.17513
R37373 VSS.n703 VSS.n688 0.173395
R37374 VSS.n3511 VSS.n769 0.173395
R37375 VSS.n3998 VSS.n3997 0.172211
R37376 VSS.n3862 VSS.n3861 0.1715
R37377 VSS.n3557 VSS.n3556 0.1715
R37378 VSS.n3807 VSS.n3804 0.1715
R37379 VSS.n3850 VSS.n3849 0.1715
R37380 VSS.n3806 VSS.n3805 0.1715
R37381 VSS.n3833 VSS.n3832 0.1715
R37382 VSS.n3835 VSS.n3834 0.1715
R37383 VSS.n3836 VSS.n3821 0.1715
R37384 VSS.n3838 VSS.n3837 0.1715
R37385 VSS.n3830 VSS.n3828 0.1715
R37386 VSS.n3829 VSS.n603 0.1715
R37387 VSS.n4035 VSS.n4034 0.1715
R37388 VSS.n4174 VSS.n4172 0.16925
R37389 VSS.n4178 VSS.n4176 0.1685
R37390 VSS.n4176 VSS.n4174 0.1685
R37391 VSS.n4170 VSS.n4168 0.1685
R37392 VSS.n4168 VSS.n4166 0.1685
R37393 VSS.n4166 VSS.n4164 0.1685
R37394 VSS.n4164 VSS.n4162 0.1685
R37395 VSS.n4172 VSS.n4170 0.16775
R37396 VSS.n2188 VSS.n1651 0.167474
R37397 VSS.n4021 VSS.n3875 0.161875
R37398 VSS.n3829 VSS.n604 0.156816
R37399 VSS.n675 VSS.n674 0.156816
R37400 VSS.n2109 VSS.n2105 0.156816
R37401 VSS.n1888 VSS.n1659 0.156816
R37402 VSS.n892 VSS.n757 0.155632
R37403 VSS.n2241 VSS.n2240 0.154584
R37404 VSS.n3415 VSS.n3414 0.153263
R37405 VSS.n1751 VSS.n801 0.147342
R37406 VSS.n4125 VSS.n468 0.146158
R37407 VSS.n3856 VSS.n713 0.146158
R37408 VSS.n1739 VSS.n1738 0.146158
R37409 VSS.n945 VSS.n944 0.146158
R37410 VSS.n2110 VSS.n2100 0.144974
R37411 VSS.n2183 VSS.n2182 0.144974
R37412 VSS.n3997 VSS.n471 0.144944
R37413 VSS.n3560 VSS.n471 0.144944
R37414 VSS.n4149 VSS.n4148 0.140237
R37415 VSS.n3857 VSS.n3855 0.140237
R37416 VSS.n1752 VSS.n1704 0.140237
R37417 VSS.n3420 VSS.n898 0.140237
R37418 VSS.n2183 VSS.n1658 0.140237
R37419 VSS.n4009 VSS.n3880 0.1355
R37420 VSS.n4010 VSS.n4009 0.1355
R37421 VSS.n4012 VSS.n4010 0.1355
R37422 VSS.n4012 VSS.n4011 0.1355
R37423 VSS.n4011 VSS.n3876 0.1355
R37424 VSS.n4019 VSS.n3876 0.1355
R37425 VSS.n4020 VSS.n4019 0.1355
R37426 VSS.n1762 VSS.n768 0.1355
R37427 VSS.n2068 VSS.n1636 0.1355
R37428 VSS.n2069 VSS.n2068 0.1355
R37429 VSS.n2070 VSS.n2069 0.1355
R37430 VSS.n2070 VSS.n2063 0.1355
R37431 VSS.n2063 VSS.n2062 0.1355
R37432 VSS.n2062 VSS.n2052 0.1355
R37433 VSS.n2088 VSS.n2052 0.1355
R37434 VSS.n2089 VSS.n2088 0.1355
R37435 VSS.n2090 VSS.n2089 0.1355
R37436 VSS.n2090 VSS.n2050 0.1355
R37437 VSS.n2050 VSS.n2049 0.1355
R37438 VSS.n2049 VSS.n2048 0.1355
R37439 VSS.n2048 VSS.n2045 0.1355
R37440 VSS.n2045 VSS.n2031 0.1355
R37441 VSS.n2115 VSS.n2031 0.1355
R37442 VSS.n2116 VSS.n2115 0.1355
R37443 VSS.n2117 VSS.n2116 0.1355
R37444 VSS.n2117 VSS.n2029 0.1355
R37445 VSS.n2029 VSS.n2028 0.1355
R37446 VSS.n2028 VSS.n2027 0.1355
R37447 VSS.n2027 VSS.n2014 0.1355
R37448 VSS.n2017 VSS.n2014 0.1355
R37449 VSS.n2017 VSS.n2016 0.1355
R37450 VSS.n2016 VSS.n1993 0.1355
R37451 VSS.n2134 VSS.n1993 0.1355
R37452 VSS.n2135 VSS.n2134 0.1355
R37453 VSS.n2136 VSS.n2135 0.1355
R37454 VSS.n2136 VSS.n1991 0.1355
R37455 VSS.n1991 VSS.n1990 0.1355
R37456 VSS.n1718 VSS.n1678 0.1355
R37457 VSS.n1719 VSS.n1718 0.1355
R37458 VSS.n1719 VSS.n1717 0.1355
R37459 VSS.n1730 VSS.n1717 0.1355
R37460 VSS.n1731 VSS.n1730 0.1355
R37461 VSS.n1732 VSS.n1731 0.1355
R37462 VSS.n1732 VSS.n1709 0.1355
R37463 VSS.n1743 VSS.n1709 0.1355
R37464 VSS.n1744 VSS.n1743 0.1355
R37465 VSS.n1747 VSS.n1744 0.1355
R37466 VSS.n1747 VSS.n1746 0.1355
R37467 VSS.n1746 VSS.n1745 0.1355
R37468 VSS.n1745 VSS.n808 0.1355
R37469 VSS.n3484 VSS.n808 0.1355
R37470 VSS.n3484 VSS.n3483 0.1355
R37471 VSS.n3483 VSS.n3482 0.1355
R37472 VSS.n1833 VSS.n1832 0.1355
R37473 VSS.n1834 VSS.n1833 0.1355
R37474 VSS.n1835 VSS.n1834 0.1355
R37475 VSS.n1836 VSS.n1835 0.1355
R37476 VSS.n1837 VSS.n1836 0.1355
R37477 VSS.n1838 VSS.n1837 0.1355
R37478 VSS.n1839 VSS.n1838 0.1355
R37479 VSS.n1840 VSS.n1839 0.1355
R37480 VSS.n2173 VSS.n2172 0.1355
R37481 VSS.n2172 VSS.n2171 0.1355
R37482 VSS.n2171 VSS.n2170 0.1355
R37483 VSS.n2170 VSS.n2169 0.1355
R37484 VSS.n2169 VSS.n2168 0.1355
R37485 VSS.n2168 VSS.n2167 0.1355
R37486 VSS.n2167 VSS.n2166 0.1355
R37487 VSS.n2166 VSS.n2165 0.1355
R37488 VSS.n2165 VSS.n2164 0.1355
R37489 VSS.n2164 VSS.n2163 0.1355
R37490 VSS.n2163 VSS.n2162 0.1355
R37491 VSS.n2162 VSS.n2161 0.1355
R37492 VSS.n2161 VSS.n2160 0.1355
R37493 VSS.n2160 VSS.n2159 0.1355
R37494 VSS.n2159 VSS.n2158 0.1355
R37495 VSS.n2158 VSS.n1855 0.1355
R37496 VSS.n1967 VSS.n1966 0.1355
R37497 VSS.n1966 VSS.n1965 0.1355
R37498 VSS.n1965 VSS.n1964 0.1355
R37499 VSS.n1964 VSS.n1963 0.1355
R37500 VSS.n1963 VSS.n1962 0.1355
R37501 VSS.n1962 VSS.n1961 0.1355
R37502 VSS.n1961 VSS.n1960 0.1355
R37503 VSS.n1960 VSS.n1959 0.1355
R37504 VSS.n1959 VSS.n1958 0.1355
R37505 VSS.n1958 VSS.n1957 0.1355
R37506 VSS.n1957 VSS.n1956 0.1355
R37507 VSS.n1956 VSS.n1955 0.1355
R37508 VSS.n1955 VSS.n1954 0.1355
R37509 VSS.n1954 VSS.n1953 0.1355
R37510 VSS.n1953 VSS.n1952 0.1355
R37511 VSS.n1952 VSS.n1951 0.1355
R37512 VSS.n1951 VSS.n1950 0.1355
R37513 VSS.n2111 VSS.n2110 0.1355
R37514 VSS.n2215 VSS.n2214 0.1355
R37515 VSS.n2216 VSS.n2215 0.1355
R37516 VSS.n2217 VSS.n2216 0.1355
R37517 VSS.n2218 VSS.n2217 0.1355
R37518 VSS.n2219 VSS.n2218 0.1355
R37519 VSS.n2220 VSS.n2219 0.1355
R37520 VSS.n2221 VSS.n2220 0.1355
R37521 VSS.n2222 VSS.n2221 0.1355
R37522 VSS.n2223 VSS.n2222 0.1355
R37523 VSS.n2224 VSS.n2223 0.1355
R37524 VSS.n2225 VSS.n2224 0.1355
R37525 VSS.n2226 VSS.n2225 0.1355
R37526 VSS.n2227 VSS.n2226 0.1355
R37527 VSS.n1648 VSS.n1647 0.1355
R37528 VSS.n1649 VSS.n1648 0.1355
R37529 VSS.n1650 VSS.n1649 0.1355
R37530 VSS.n1792 VSS.n1650 0.1355
R37531 VSS.n1793 VSS.n1792 0.1355
R37532 VSS.n1793 VSS.n1791 0.1355
R37533 VSS.n1784 VSS.n1783 0.1355
R37534 VSS.n1785 VSS.n1784 0.1355
R37535 VSS.n1786 VSS.n1785 0.1355
R37536 VSS.n1787 VSS.n1786 0.1355
R37537 VSS.n1788 VSS.n1787 0.1355
R37538 VSS.n870 VSS.n868 0.1355
R37539 VSS.n868 VSS.n866 0.1355
R37540 VSS.n866 VSS.n864 0.1355
R37541 VSS.n864 VSS.n862 0.1355
R37542 VSS.n862 VSS.n860 0.1355
R37543 VSS.n860 VSS.n858 0.1355
R37544 VSS.n858 VSS.n856 0.1355
R37545 VSS.n856 VSS.n854 0.1355
R37546 VSS.n854 VSS.n852 0.1355
R37547 VSS.n852 VSS.n850 0.1355
R37548 VSS.n850 VSS.n848 0.1355
R37549 VSS.n848 VSS.n846 0.1355
R37550 VSS.n846 VSS.n844 0.1355
R37551 VSS.n844 VSS.n842 0.1355
R37552 VSS.n842 VSS.n840 0.1355
R37553 VSS.n840 VSS.n838 0.1355
R37554 VSS.n838 VSS.n836 0.1355
R37555 VSS.n836 VSS.n834 0.1355
R37556 VSS.n834 VSS.n832 0.1355
R37557 VSS.n832 VSS.n830 0.1355
R37558 VSS.n830 VSS.n828 0.1355
R37559 VSS.n828 VSS.n826 0.1355
R37560 VSS.n826 VSS.n824 0.1355
R37561 VSS.n824 VSS.n822 0.1355
R37562 VSS.n822 VSS.n820 0.1355
R37563 VSS.n820 VSS.n818 0.1355
R37564 VSS.n818 VSS.n816 0.1355
R37565 VSS.n816 VSS.n815 0.1355
R37566 VSS.n815 VSS.n814 0.1355
R37567 VSS.n3431 VSS.n729 0.1355
R37568 VSS.n3432 VSS.n3431 0.1355
R37569 VSS.n3433 VSS.n3432 0.1355
R37570 VSS.n3434 VSS.n3433 0.1355
R37571 VSS.n3435 VSS.n3434 0.1355
R37572 VSS.n3436 VSS.n3435 0.1355
R37573 VSS.n3437 VSS.n3436 0.1355
R37574 VSS.n3438 VSS.n3437 0.1355
R37575 VSS.n3439 VSS.n3438 0.1355
R37576 VSS.n3440 VSS.n3439 0.1355
R37577 VSS.n3441 VSS.n3440 0.1355
R37578 VSS.n3442 VSS.n3441 0.1355
R37579 VSS.n3443 VSS.n3442 0.1355
R37580 VSS.n3444 VSS.n3443 0.1355
R37581 VSS.n3445 VSS.n3444 0.1355
R37582 VSS.n3446 VSS.n3445 0.1355
R37583 VSS.n3447 VSS.n3446 0.1355
R37584 VSS.n3868 VSS.n3549 0.1355
R37585 VSS.n3868 VSS.n3867 0.1355
R37586 VSS.n3867 VSS.n3866 0.1355
R37587 VSS.n3866 VSS.n3551 0.1355
R37588 VSS.n3811 VSS.n3551 0.1355
R37589 VSS.n3814 VSS.n3811 0.1355
R37590 VSS.n3815 VSS.n3814 0.1355
R37591 VSS.n3816 VSS.n3815 0.1355
R37592 VSS.n3844 VSS.n3816 0.1355
R37593 VSS.n3844 VSS.n3843 0.1355
R37594 VSS.n3843 VSS.n3842 0.1355
R37595 VSS.n3842 VSS.n3818 0.1355
R37596 VSS.n3823 VSS.n3818 0.1355
R37597 VSS.n3824 VSS.n3823 0.1355
R37598 VSS.n3824 VSS.n600 0.1355
R37599 VSS.n4039 VSS.n600 0.1355
R37600 VSS.n4040 VSS.n4039 0.1355
R37601 VSS.n3547 VSS.n3546 0.1355
R37602 VSS.n3546 VSS.n3545 0.1355
R37603 VSS.n3545 VSS.n3544 0.1355
R37604 VSS.n3544 VSS.n3543 0.1355
R37605 VSS.n3543 VSS.n3542 0.1355
R37606 VSS.n3542 VSS.n3541 0.1355
R37607 VSS.n3541 VSS.n3540 0.1355
R37608 VSS.n3540 VSS.n3539 0.1355
R37609 VSS.n3539 VSS.n3538 0.1355
R37610 VSS.n3538 VSS.n3537 0.1355
R37611 VSS.n741 VSS.n740 0.1355
R37612 VSS.n742 VSS.n741 0.1355
R37613 VSS.n743 VSS.n742 0.1355
R37614 VSS.n3873 VSS.n3872 0.1355
R37615 VSS.n3872 VSS.n715 0.1355
R37616 VSS.n529 VSS.n527 0.1355
R37617 VSS.n531 VSS.n529 0.1355
R37618 VSS.n533 VSS.n531 0.1355
R37619 VSS.n535 VSS.n533 0.1355
R37620 VSS.n537 VSS.n535 0.1355
R37621 VSS.n539 VSS.n537 0.1355
R37622 VSS.n541 VSS.n539 0.1355
R37623 VSS.n543 VSS.n541 0.1355
R37624 VSS.n545 VSS.n543 0.1355
R37625 VSS.n547 VSS.n545 0.1355
R37626 VSS.n549 VSS.n547 0.1355
R37627 VSS.n551 VSS.n549 0.1355
R37628 VSS.n553 VSS.n551 0.1355
R37629 VSS.n555 VSS.n553 0.1355
R37630 VSS.n557 VSS.n555 0.1355
R37631 VSS.n559 VSS.n557 0.1355
R37632 VSS.n561 VSS.n559 0.1355
R37633 VSS.n563 VSS.n561 0.1355
R37634 VSS.n565 VSS.n563 0.1355
R37635 VSS.n567 VSS.n565 0.1355
R37636 VSS.n569 VSS.n567 0.1355
R37637 VSS.n571 VSS.n569 0.1355
R37638 VSS.n573 VSS.n571 0.1355
R37639 VSS.n575 VSS.n573 0.1355
R37640 VSS.n577 VSS.n575 0.1355
R37641 VSS.n579 VSS.n577 0.1355
R37642 VSS.n581 VSS.n579 0.1355
R37643 VSS.n583 VSS.n581 0.1355
R37644 VSS.n585 VSS.n583 0.1355
R37645 VSS.n587 VSS.n585 0.1355
R37646 VSS.n589 VSS.n587 0.1355
R37647 VSS.n591 VSS.n589 0.1355
R37648 VSS.n593 VSS.n591 0.1355
R37649 VSS.n595 VSS.n593 0.1355
R37650 VSS.n598 VSS.n595 0.1355
R37651 VSS.n4097 VSS.n4096 0.1355
R37652 VSS.n4096 VSS.n4095 0.1355
R37653 VSS.n4095 VSS.n4094 0.1355
R37654 VSS.n4094 VSS.n4093 0.1355
R37655 VSS.n4093 VSS.n4092 0.1355
R37656 VSS.n4092 VSS.n4091 0.1355
R37657 VSS.n4091 VSS.n4090 0.1355
R37658 VSS.n4090 VSS.n4089 0.1355
R37659 VSS.n4089 VSS.n4088 0.1355
R37660 VSS.n4088 VSS.n4087 0.1355
R37661 VSS.n4087 VSS.n4086 0.1355
R37662 VSS.n4086 VSS.n4085 0.1355
R37663 VSS.n4085 VSS.n4084 0.1355
R37664 VSS.n4084 VSS.n4083 0.1355
R37665 VSS.n4083 VSS.n4082 0.1355
R37666 VSS.n4082 VSS.n4081 0.1355
R37667 VSS.n508 VSS.n506 0.1355
R37668 VSS.n506 VSS.n504 0.1355
R37669 VSS.n504 VSS.n502 0.1355
R37670 VSS.n502 VSS.n500 0.1355
R37671 VSS.n500 VSS.n498 0.1355
R37672 VSS.n498 VSS.n496 0.1355
R37673 VSS.n496 VSS.n494 0.1355
R37674 VSS.n494 VSS.n492 0.1355
R37675 VSS.n492 VSS.n490 0.1355
R37676 VSS.n490 VSS.n488 0.1355
R37677 VSS.n488 VSS.n486 0.1355
R37678 VSS.n486 VSS.n485 0.1355
R37679 VSS.n3976 VSS.n3915 0.1355
R37680 VSS.n3977 VSS.n3976 0.1355
R37681 VSS.n3978 VSS.n3977 0.1355
R37682 VSS.n3984 VSS.n3978 0.1355
R37683 VSS.n3984 VSS.n3983 0.1355
R37684 VSS.n3983 VSS.n3982 0.1355
R37685 VSS.n3982 VSS.n482 0.1355
R37686 VSS.n4136 VSS.n482 0.1355
R37687 VSS.n4136 VSS.n4135 0.1355
R37688 VSS.n4135 VSS.n4134 0.1355
R37689 VSS.n4134 VSS.n4133 0.1355
R37690 VSS.n3934 VSS.n3933 0.1355
R37691 VSS.n3935 VSS.n3934 0.1355
R37692 VSS.n3936 VSS.n3935 0.1355
R37693 VSS.n3937 VSS.n3936 0.1355
R37694 VSS.n3938 VSS.n3937 0.1355
R37695 VSS.n3939 VSS.n3938 0.1355
R37696 VSS.n3940 VSS.n3939 0.1355
R37697 VSS.n3941 VSS.n3940 0.1355
R37698 VSS.n3942 VSS.n3941 0.1355
R37699 VSS.n3943 VSS.n3942 0.1355
R37700 VSS.n3944 VSS.n3943 0.1355
R37701 VSS.n3945 VSS.n3944 0.1355
R37702 VSS.n3946 VSS.n3945 0.1355
R37703 VSS.n3947 VSS.n3946 0.1355
R37704 VSS.n3948 VSS.n3947 0.1355
R37705 VSS.n3949 VSS.n3948 0.1355
R37706 VSS.n3950 VSS.n3949 0.1355
R37707 VSS.n3951 VSS.n3950 0.1355
R37708 VSS.n1358 VSS.n1357 0.1355
R37709 VSS.n1359 VSS.n1358 0.1355
R37710 VSS.n1360 VSS.n1359 0.1355
R37711 VSS.n1446 VSS.n1444 0.1355
R37712 VSS.n1448 VSS.n1446 0.1355
R37713 VSS.n1450 VSS.n1448 0.1355
R37714 VSS.n1452 VSS.n1450 0.1355
R37715 VSS.n1454 VSS.n1452 0.1355
R37716 VSS.n1456 VSS.n1454 0.1355
R37717 VSS.n1458 VSS.n1456 0.1355
R37718 VSS.n1460 VSS.n1458 0.1355
R37719 VSS.n1462 VSS.n1460 0.1355
R37720 VSS.n1464 VSS.n1462 0.1355
R37721 VSS.n1466 VSS.n1464 0.1355
R37722 VSS.n1468 VSS.n1466 0.1355
R37723 VSS.n1470 VSS.n1468 0.1355
R37724 VSS.n1472 VSS.n1470 0.1355
R37725 VSS.n1474 VSS.n1472 0.1355
R37726 VSS.n1476 VSS.n1474 0.1355
R37727 VSS.n1479 VSS.n1476 0.1355
R37728 VSS.n3056 VSS.n1479 0.1355
R37729 VSS.n3118 VSS.n3117 0.1355
R37730 VSS.n3117 VSS.n1412 0.1355
R37731 VSS.n3107 VSS.n1412 0.1355
R37732 VSS.n3107 VSS.n3106 0.1355
R37733 VSS.n3106 VSS.n3105 0.1355
R37734 VSS.n3105 VSS.n1420 0.1355
R37735 VSS.n3095 VSS.n1420 0.1355
R37736 VSS.n3095 VSS.n3094 0.1355
R37737 VSS.n3094 VSS.n3093 0.1355
R37738 VSS.n3093 VSS.n1428 0.1355
R37739 VSS.n1440 VSS.n1428 0.1355
R37740 VSS.n3082 VSS.n1440 0.1355
R37741 VSS.n3082 VSS.n3081 0.1355
R37742 VSS.n3081 VSS.n3080 0.1355
R37743 VSS.n3080 VSS.n3079 0.1355
R37744 VSS.n3079 VSS.n3078 0.1355
R37745 VSS.n3128 VSS.n3119 0.1355
R37746 VSS.n3129 VSS.n3128 0.1355
R37747 VSS.n3130 VSS.n3129 0.1355
R37748 VSS.n3158 VSS.n3130 0.1355
R37749 VSS.n3158 VSS.n3157 0.1355
R37750 VSS.n3157 VSS.n3156 0.1355
R37751 VSS.n3156 VSS.n3132 0.1355
R37752 VSS.n3141 VSS.n3132 0.1355
R37753 VSS.n3142 VSS.n3141 0.1355
R37754 VSS.n3146 VSS.n3142 0.1355
R37755 VSS.n3146 VSS.n3145 0.1355
R37756 VSS.n3145 VSS.n3144 0.1355
R37757 VSS.n3144 VSS.n1042 0.1355
R37758 VSS.n3374 VSS.n1042 0.1355
R37759 VSS.n3374 VSS.n3373 0.1355
R37760 VSS.n3373 VSS.n3372 0.1355
R37761 VSS.n3172 VSS.n3171 0.1355
R37762 VSS.n3173 VSS.n3172 0.1355
R37763 VSS.n3174 VSS.n3173 0.1355
R37764 VSS.n3175 VSS.n3174 0.1355
R37765 VSS.n3176 VSS.n3175 0.1355
R37766 VSS.n3177 VSS.n3176 0.1355
R37767 VSS.n3178 VSS.n3177 0.1355
R37768 VSS.n3179 VSS.n3178 0.1355
R37769 VSS.n1104 VSS.n1102 0.1355
R37770 VSS.n1102 VSS.n1100 0.1355
R37771 VSS.n1100 VSS.n1098 0.1355
R37772 VSS.n1098 VSS.n1096 0.1355
R37773 VSS.n1096 VSS.n1094 0.1355
R37774 VSS.n1094 VSS.n1092 0.1355
R37775 VSS.n1092 VSS.n1090 0.1355
R37776 VSS.n1090 VSS.n1088 0.1355
R37777 VSS.n1088 VSS.n1086 0.1355
R37778 VSS.n1086 VSS.n1084 0.1355
R37779 VSS.n1084 VSS.n1082 0.1355
R37780 VSS.n1082 VSS.n1080 0.1355
R37781 VSS.n1080 VSS.n1078 0.1355
R37782 VSS.n1078 VSS.n1076 0.1355
R37783 VSS.n1076 VSS.n1074 0.1355
R37784 VSS.n1074 VSS.n1072 0.1355
R37785 VSS.n1072 VSS.n1070 0.1355
R37786 VSS.n1070 VSS.n1068 0.1355
R37787 VSS.n1068 VSS.n1066 0.1355
R37788 VSS.n1066 VSS.n1064 0.1355
R37789 VSS.n1064 VSS.n1062 0.1355
R37790 VSS.n1062 VSS.n1060 0.1355
R37791 VSS.n1060 VSS.n1058 0.1355
R37792 VSS.n1058 VSS.n1056 0.1355
R37793 VSS.n1056 VSS.n1054 0.1355
R37794 VSS.n1054 VSS.n1052 0.1355
R37795 VSS.n1052 VSS.n1050 0.1355
R37796 VSS.n1050 VSS.n1049 0.1355
R37797 VSS.n1049 VSS.n1048 0.1355
R37798 VSS.n3321 VSS.n3320 0.1355
R37799 VSS.n3322 VSS.n3321 0.1355
R37800 VSS.n3323 VSS.n3322 0.1355
R37801 VSS.n3324 VSS.n3323 0.1355
R37802 VSS.n3325 VSS.n3324 0.1355
R37803 VSS.n3326 VSS.n3325 0.1355
R37804 VSS.n3327 VSS.n3326 0.1355
R37805 VSS.n3328 VSS.n3327 0.1355
R37806 VSS.n3329 VSS.n3328 0.1355
R37807 VSS.n3330 VSS.n3329 0.1355
R37808 VSS.n3331 VSS.n3330 0.1355
R37809 VSS.n3332 VSS.n3331 0.1355
R37810 VSS.n3333 VSS.n3332 0.1355
R37811 VSS.n3334 VSS.n3333 0.1355
R37812 VSS.n3335 VSS.n3334 0.1355
R37813 VSS.n3336 VSS.n3335 0.1355
R37814 VSS.n3337 VSS.n3336 0.1355
R37815 VSS.n1149 VSS.n1148 0.1355
R37816 VSS.n1148 VSS.n1147 0.1355
R37817 VSS.n1147 VSS.n1146 0.1355
R37818 VSS.n1146 VSS.n1145 0.1355
R37819 VSS.n1145 VSS.n1144 0.1355
R37820 VSS.n1144 VSS.n1143 0.1355
R37821 VSS.n1143 VSS.n1142 0.1355
R37822 VSS.n1142 VSS.n1141 0.1355
R37823 VSS.n1141 VSS.n1140 0.1355
R37824 VSS.n1140 VSS.n1124 0.1355
R37825 VSS.n1352 VSS.n1351 0.1355
R37826 VSS.n1351 VSS.n1350 0.1355
R37827 VSS.n1350 VSS.n1349 0.1355
R37828 VSS.n1349 VSS.n1348 0.1355
R37829 VSS.n1348 VSS.n1347 0.1355
R37830 VSS.n1347 VSS.n1346 0.1355
R37831 VSS.n1346 VSS.n1345 0.1355
R37832 VSS.n1345 VSS.n1344 0.1355
R37833 VSS.n1344 VSS.n1343 0.1355
R37834 VSS.n1343 VSS.n1342 0.1355
R37835 VSS.n1342 VSS.n1341 0.1355
R37836 VSS.n1341 VSS.n1340 0.1355
R37837 VSS.n1340 VSS.n1339 0.1355
R37838 VSS.n1339 VSS.n1338 0.1355
R37839 VSS.n1338 VSS.n1337 0.1355
R37840 VSS.n1337 VSS.n1336 0.1355
R37841 VSS.n1336 VSS.n1335 0.1355
R37842 VSS.n1294 VSS.n1293 0.1355
R37843 VSS.n1293 VSS.n1292 0.1355
R37844 VSS.n1292 VSS.n1291 0.1355
R37845 VSS.n1291 VSS.n1290 0.1355
R37846 VSS.n1290 VSS.n1289 0.1355
R37847 VSS.n1289 VSS.n1288 0.1355
R37848 VSS.n1288 VSS.n1287 0.1355
R37849 VSS.n1287 VSS.n1286 0.1355
R37850 VSS.n1286 VSS.n1285 0.1355
R37851 VSS.n1285 VSS.n1284 0.1355
R37852 VSS.n1284 VSS.n1283 0.1355
R37853 VSS.n1283 VSS.n1282 0.1355
R37854 VSS.n1282 VSS.n1281 0.1355
R37855 VSS.n1281 VSS.n1280 0.1355
R37856 VSS.n1280 VSS.n1279 0.1355
R37857 VSS.n1279 VSS.n1278 0.1355
R37858 VSS.n1278 VSS.n1277 0.1355
R37859 VSS.n1277 VSS.n1276 0.1355
R37860 VSS.n1276 VSS.n1275 0.1355
R37861 VSS.n1275 VSS.n1274 0.1355
R37862 VSS.n1274 VSS.n1273 0.1355
R37863 VSS.n1273 VSS.n1272 0.1355
R37864 VSS.n1272 VSS.n1271 0.1355
R37865 VSS.n1271 VSS.n1270 0.1355
R37866 VSS.n1270 VSS.n1269 0.1355
R37867 VSS.n1269 VSS.n1268 0.1355
R37868 VSS.n1268 VSS.n1267 0.1355
R37869 VSS.n1267 VSS.n1266 0.1355
R37870 VSS.n1266 VSS.n1265 0.1355
R37871 VSS.n1265 VSS.n1264 0.1355
R37872 VSS.n1264 VSS.n1263 0.1355
R37873 VSS.n1263 VSS.n1262 0.1355
R37874 VSS.n1262 VSS.n1261 0.1355
R37875 VSS.n1261 VSS.n1260 0.1355
R37876 VSS.n1260 VSS.n1259 0.1355
R37877 VSS.n3761 VSS.n3760 0.1355
R37878 VSS.n3760 VSS.n3722 0.1355
R37879 VSS.n3735 VSS.n3722 0.1355
R37880 VSS.n3736 VSS.n3735 0.1355
R37881 VSS.n3748 VSS.n3736 0.1355
R37882 VSS.n3748 VSS.n3747 0.1355
R37883 VSS.n3747 VSS.n3746 0.1355
R37884 VSS.n3746 VSS.n3737 0.1355
R37885 VSS.n3737 VSS.n448 0.1355
R37886 VSS.n4187 VSS.n448 0.1355
R37887 VSS.n3720 VSS.n3718 0.1355
R37888 VSS.n3718 VSS.n3716 0.1355
R37889 VSS.n3716 VSS.n3714 0.1355
R37890 VSS.n3714 VSS.n3712 0.1355
R37891 VSS.n3712 VSS.n3710 0.1355
R37892 VSS.n3710 VSS.n3708 0.1355
R37893 VSS.n3708 VSS.n3706 0.1355
R37894 VSS.n3706 VSS.n3704 0.1355
R37895 VSS.n3704 VSS.n3702 0.1355
R37896 VSS.n3702 VSS.n3700 0.1355
R37897 VSS.n3700 VSS.n3698 0.1355
R37898 VSS.n3698 VSS.n3694 0.1355
R37899 VSS.n3667 VSS.n3666 0.1355
R37900 VSS.n3668 VSS.n3667 0.1355
R37901 VSS.n3668 VSS.n3578 0.1355
R37902 VSS.n3678 VSS.n3578 0.1355
R37903 VSS.n3679 VSS.n3678 0.1355
R37904 VSS.n3681 VSS.n3679 0.1355
R37905 VSS.n3681 VSS.n3680 0.1355
R37906 VSS.n3680 VSS.n3569 0.1355
R37907 VSS.n3692 VSS.n3569 0.1355
R37908 VSS.n3693 VSS.n3692 0.1355
R37909 VSS.n3787 VSS.n3693 0.1355
R37910 VSS.n3625 VSS.n3624 0.1355
R37911 VSS.n3626 VSS.n3625 0.1355
R37912 VSS.n3627 VSS.n3626 0.1355
R37913 VSS.n3628 VSS.n3627 0.1355
R37914 VSS.n3629 VSS.n3628 0.1355
R37915 VSS.n3630 VSS.n3629 0.1355
R37916 VSS.n3631 VSS.n3630 0.1355
R37917 VSS.n3632 VSS.n3631 0.1355
R37918 VSS.n3633 VSS.n3632 0.1355
R37919 VSS.n3634 VSS.n3633 0.1355
R37920 VSS.n3635 VSS.n3634 0.1355
R37921 VSS.n3636 VSS.n3635 0.1355
R37922 VSS.n3637 VSS.n3636 0.1355
R37923 VSS.n3638 VSS.n3637 0.1355
R37924 VSS.n3639 VSS.n3638 0.1355
R37925 VSS.n3640 VSS.n3639 0.1355
R37926 VSS.n3641 VSS.n3640 0.1355
R37927 VSS.n3642 VSS.n3641 0.1355
R37928 VSS.n1616 VSS.n1615 0.1355
R37929 VSS.n1615 VSS.n1614 0.1355
R37930 VSS.n1614 VSS.n1613 0.1355
R37931 VSS.n1613 VSS.n1612 0.1355
R37932 VSS.n1612 VSS.n1611 0.1355
R37933 VSS.n1611 VSS.n1610 0.1355
R37934 VSS.n1610 VSS.n1609 0.1355
R37935 VSS.n1609 VSS.n1608 0.1355
R37936 VSS.n1608 VSS.n1607 0.1355
R37937 VSS.n1607 VSS.n1606 0.1355
R37938 VSS.n1606 VSS.n1605 0.1355
R37939 VSS.n1605 VSS.n1604 0.1355
R37940 VSS.n1604 VSS.n1508 0.1355
R37941 VSS.n2264 VSS.n2263 0.1355
R37942 VSS.n2265 VSS.n2264 0.1355
R37943 VSS.n2266 VSS.n2265 0.1355
R37944 VSS.n2267 VSS.n2266 0.1355
R37945 VSS.n2268 VSS.n2267 0.1355
R37946 VSS.n2269 VSS.n2268 0.1355
R37947 VSS.n2270 VSS.n2269 0.1355
R37948 VSS.n2271 VSS.n2270 0.1355
R37949 VSS.n2272 VSS.n2271 0.1355
R37950 VSS.n2273 VSS.n2272 0.1355
R37951 VSS.n2274 VSS.n2273 0.1355
R37952 VSS.n2275 VSS.n2274 0.1355
R37953 VSS.n2276 VSS.n2275 0.1355
R37954 VSS.n2277 VSS.n2276 0.1355
R37955 VSS.n2278 VSS.n2277 0.1355
R37956 VSS.n2279 VSS.n2278 0.1355
R37957 VSS.n2280 VSS.n2279 0.1355
R37958 VSS.n2281 VSS.n2280 0.1355
R37959 VSS.n2282 VSS.n2281 0.1355
R37960 VSS.n2283 VSS.n2282 0.1355
R37961 VSS.n2284 VSS.n2283 0.1355
R37962 VSS.n2285 VSS.n2284 0.1355
R37963 VSS.n2286 VSS.n2285 0.1355
R37964 VSS.n3851 VSS.n3804 0.134316
R37965 VSS.n628 VSS.n627 0.134316
R37966 VSS.n1940 VSS.n1939 0.134316
R37967 VSS.n2237 VSS.n2236 0.134316
R37968 VSS.n2141 VSS.n1944 0.13325
R37969 VSS.n2142 VSS.n1942 0.13325
R37970 VSS.n2143 VSS.n1940 0.13325
R37971 VSS.n2144 VSS.n1937 0.13325
R37972 VSS.n2145 VSS.n1935 0.13325
R37973 VSS.n2146 VSS.n1933 0.13325
R37974 VSS.n2147 VSS.n1931 0.13325
R37975 VSS.n2148 VSS.n1929 0.13325
R37976 VSS.n2149 VSS.n1927 0.13325
R37977 VSS.n2150 VSS.n1923 0.13325
R37978 VSS.n2151 VSS.n1921 0.13325
R37979 VSS.n2152 VSS.n1919 0.13325
R37980 VSS.n4014 VSS.n3878 0.130763
R37981 VSS.n4158 VSS.n4157 0.1305
R37982 VSS.n4159 VSS.n4158 0.1305
R37983 VSS.n3831 VSS.n3830 0.129579
R37984 VSS.n617 VSS.n608 0.129579
R37985 VSS.n1926 VSS.n1923 0.128395
R37986 VSS.n2197 VSS.n2196 0.128395
R37987 VSS.n2083 VSS.n2077 0.120105
R37988 VSS.n1393 VSS.n1375 0.119
R37989 VSS.n4143 VSS.n472 0.117737
R37990 VSS.n4025 VSS.n711 0.117737
R37991 VSS.n1824 VSS.n1686 0.117737
R37992 VSS.n3426 VSS.n3425 0.117737
R37993 VSS.n2189 VSS.n2188 0.117737
R37994 VSS.n754 VSS.n736 0.11329
R37995 VSS.n1832 VSS.n1831 0.113
R37996 VSS.n2174 VSS.n1840 0.113
R37997 VSS.n1790 VSS.n1788 0.113
R37998 VSS.n3548 VSS.n3547 0.113
R37999 VSS.n3537 VSS.n3536 0.113
R38000 VSS.n4132 VSS.n485 0.113
R38001 VSS.n3056 VSS.n3055 0.113
R38002 VSS.n3171 VSS.n3170 0.113
R38003 VSS.n3180 VSS.n3179 0.113
R38004 VSS.n1353 VSS.n1149 0.113
R38005 VSS.n3319 VSS.n1124 0.113
R38006 VSS.n3786 VSS.n3694 0.113
R38007 VSS.n4031 VSS.n4030 0.110632
R38008 VSS.n4034 VSS.n4033 0.109447
R38009 VSS.n3407 VSS.n1014 0.109447
R38010 VSS.n2004 VSS.n2002 0.109447
R38011 VSS.n1917 VSS.n1916 0.109447
R38012 VSS.n3403 VSS.n764 0.107079
R38013 VSS.n2124 VSS.n2123 0.103526
R38014 VSS.n1881 VSS.n1879 0.103526
R38015 VSS.n4157 VSS.n460 0.102342
R38016 VSS.n2100 VSS.n2037 0.0928684
R38017 VSS.n738 VSS.n715 0.0905
R38018 VSS.n1180 VSS.n1139 0.0905
R38019 VSS.n3874 VSS.n3873 0.089375
R38020 VSS.n4157 VSS.n4156 0.0881316
R38021 VSS.n1772 VSS.n1688 0.0876667
R38022 VSS.n2124 VSS.n2007 0.0869474
R38023 VSS.n1891 VSS.n1881 0.0869474
R38024 VSS.n3206 VSS.n3205 0.0864511
R38025 VSS.n705 VSS.n703 0.0857459
R38026 VSS.n705 VSS.n704 0.0857459
R38027 VSS.n3403 VSS.n763 0.0833947
R38028 VSS.n3055 VSS.n1482 0.0813572
R38029 VSS.n3055 VSS.n1483 0.0813572
R38030 VSS.n3055 VSS.n1480 0.0813572
R38031 VSS.n1258 VSS.n447 0.0813572
R38032 VSS.n1243 VSS.n447 0.0813572
R38033 VSS.n1246 VSS.n447 0.0813572
R38034 VSS.n3408 VSS.n3407 0.0810263
R38035 VSS.n2004 VSS.n2003 0.0810263
R38036 VSS.n1918 VSS.n1917 0.0810263
R38037 VSS.n2110 VSS.n2109 0.0810263
R38038 VSS.n2182 VSS.n1659 0.0810263
R38039 VSS.n3205 VSS.n3204 0.0808261
R38040 VSS.n4030 VSS.n605 0.0798421
R38041 VSS.n1296 VSS.n1295 0.0792609
R38042 VSS.n3290 VSS.n1016 0.0781429
R38043 VSS.n3247 VSS.n1016 0.0781429
R38044 VSS.n3687 VSS.n3561 0.0749828
R38045 VSS.n4143 VSS.n4142 0.0727368
R38046 VSS.n4025 VSS.n4024 0.0727368
R38047 VSS.n1724 VSS.n1686 0.0727368
R38048 VSS.n3425 VSS.n891 0.0727368
R38049 VSS.n2077 VSS.n2076 0.0703684
R38050 VSS.n3741 VSS.n456 0.0697308
R38051 VSS.n3793 VSS.n3792 0.0693966
R38052 VSS.n1831 VSS.n1678 0.068
R38053 VSS.n2174 VSS.n2173 0.068
R38054 VSS.n1791 VSS.n1790 0.068
R38055 VSS.n3536 VSS.n729 0.068
R38056 VSS.n3549 VSS.n3548 0.068
R38057 VSS.n4133 VSS.n4132 0.068
R38058 VSS.n3180 VSS.n3118 0.068
R38059 VSS.n3170 VSS.n3119 0.068
R38060 VSS.n3320 VSS.n3319 0.068
R38061 VSS.n1353 VSS.n1352 0.068
R38062 VSS.n3787 VSS.n3786 0.068
R38063 VSS.n3419 VSS.n3418 0.067693
R38064 VSS.n1248 VSS.n1246 0.0652857
R38065 VSS.n1256 VSS.n1243 0.0652857
R38066 VSS.n1297 VSS.n1258 0.0652857
R38067 VSS.n1522 VSS.n1482 0.0652857
R38068 VSS.n1551 VSS.n1482 0.0652857
R38069 VSS.n1550 VSS.n1483 0.0652857
R38070 VSS.n1547 VSS.n1483 0.0652857
R38071 VSS.n1546 VSS.n1480 0.0652857
R38072 VSS.n3057 VSS.n1480 0.0652857
R38073 VSS.n1246 VSS.n450 0.0652857
R38074 VSS.n1247 VSS.n1243 0.0652857
R38075 VSS.n1258 VSS.n1257 0.0652857
R38076 VSS.n1181 VSS.n1179 0.0645294
R38077 VSS.n3512 VSS.n3511 0.0644474
R38078 VSS.n3400 VSS.n1016 0.0636786
R38079 VSS.n3504 VSS.n777 0.0620789
R38080 VSS.n1927 VSS.n1926 0.0620789
R38081 VSS.n2198 VSS.n2197 0.0620789
R38082 VSS.n4080 VSS.n4079 0.061
R38083 VSS.n4099 VSS.n510 0.061
R38084 VSS.n4022 VSS.n4021 0.061
R38085 VSS.n3449 VSS.n872 0.061
R38086 VSS.n3516 VSS.n3515 0.061
R38087 VSS.n3518 VSS.n766 0.061
R38088 VSS.n1969 VSS.n1968 0.061
R38089 VSS.n1989 VSS.n1988 0.061
R38090 VSS.n2213 VSS.n2212 0.061
R38091 VSS.n2229 VSS.n2228 0.061
R38092 VSS.n811 VSS.n810 0.061
R38093 VSS.n4042 VSS.n4041 0.061
R38094 VSS.n3932 VSS.n3931 0.061
R38095 VSS.n3953 VSS.n3952 0.061
R38096 VSS.n3339 VSS.n1106 0.061
R38097 VSS.n1372 VSS.n1371 0.061
R38098 VSS.n3208 VSS.n1374 0.061
R38099 VSS.n3077 VSS.n3076 0.061
R38100 VSS.n1617 VSS.n1603 0.061
R38101 VSS.n2262 VSS.n2261 0.061
R38102 VSS.n1045 VSS.n1044 0.061
R38103 VSS.n1168 VSS.n1167 0.061
R38104 VSS.n3587 VSS.n3586 0.061
R38105 VSS.n3643 VSS.n3623 0.061
R38106 VSS.n3763 VSS.n3762 0.061
R38107 VSS.n3837 VSS.n3831 0.0608947
R38108 VSS.n618 VSS.n617 0.0608947
R38109 VSS.n4182 VSS.n4181 0.0602115
R38110 VSS.n3645 VSS.n3644 0.0594563
R38111 VSS.n3388 VSS.n3387 0.058254
R38112 VSS.n3851 VSS.n3850 0.0561579
R38113 VSS.n627 VSS.n620 0.0561579
R38114 VSS.n1939 VSS.n1937 0.0561579
R38115 VSS.n2237 VSS.n1624 0.0561579
R38116 VSS.n3781 VSS.n3780 0.055
R38117 VSS.n2003 VSS.n1944 0.0549737
R38118 VSS.n1433 VSS.n1432 0.0544256
R38119 VSS.n3386 VSS.n3385 0.0541631
R38120 VSS.n3099 VSS.n1424 0.0536818
R38121 VSS.n3860 VSS.n3554 0.0508731
R38122 VSS.n3855 VSS.n3558 0.0502368
R38123 VSS.n1752 VSS.n1751 0.0502368
R38124 VSS.n3420 VSS.n3419 0.0502368
R38125 VSS.n3188 VSS.n3187 0.0500909
R38126 VSS.n1295 VSS.n447 0.049913
R38127 VSS.n739 VSS.n737 0.0455
R38128 VSS.n1356 VSS.n1355 0.0455
R38129 VSS.n4126 VSS.n4125 0.0443158
R38130 VSS.n3874 VSS.n713 0.0443158
R38131 VSS.n1738 VSS.n1737 0.0443158
R38132 VSS.n944 VSS.n943 0.0443158
R38133 VSS.n1800 VSS.n1799 0.0443158
R38134 VSS.n3860 VSS.n3558 0.0406613
R38135 VSS.n3548 VSS.n717 0.038
R38136 VSS.n1354 VSS.n1353 0.038
R38137 VSS.n3414 VSS.n3413 0.0372105
R38138 VSS.n3051 VSS.n3050 0.0369787
R38139 VSS.n3860 VSS.n3859 0.0367903
R38140 VSS.n1432 VSS.n1424 0.0365744
R38141 VSS.n4414 VSS.n4413 0.0362313
R38142 VSS.n4504 VSS.n384 0.0362313
R38143 VSS.n2860 VSS.n2859 0.0362313
R38144 VSS.n3089 VSS.n1433 0.0358306
R38145 VSS.n4412 VSS.n4411 0.0353837
R38146 VSS.n4410 VSS.n4253 0.0353837
R38147 VSS.n4409 VSS.n4254 0.0353837
R38148 VSS.n4408 VSS.n4255 0.0353837
R38149 VSS.n4407 VSS.n4256 0.0353837
R38150 VSS.n4406 VSS.n4257 0.0353837
R38151 VSS.n4405 VSS.n4258 0.0353837
R38152 VSS.n4404 VSS.n4259 0.0353837
R38153 VSS.n4403 VSS.n4260 0.0353837
R38154 VSS.n4402 VSS.n4261 0.0353837
R38155 VSS.n4401 VSS.n4262 0.0353837
R38156 VSS.n4400 VSS.n4263 0.0353837
R38157 VSS.n4399 VSS.n4264 0.0353837
R38158 VSS.n4398 VSS.n4265 0.0353837
R38159 VSS.n4397 VSS.n4266 0.0353837
R38160 VSS.n4396 VSS.n4267 0.0353837
R38161 VSS.n4395 VSS.n4268 0.0353837
R38162 VSS.n4394 VSS.n4269 0.0353837
R38163 VSS.n4393 VSS.n4270 0.0353837
R38164 VSS.n4392 VSS.n4271 0.0353837
R38165 VSS.n4391 VSS.n4272 0.0353837
R38166 VSS.n4390 VSS.n4273 0.0353837
R38167 VSS.n4389 VSS.n4274 0.0353837
R38168 VSS.n4388 VSS.n4275 0.0353837
R38169 VSS.n4387 VSS.n4276 0.0353837
R38170 VSS.n4386 VSS.n4277 0.0353837
R38171 VSS.n4385 VSS.n4278 0.0353837
R38172 VSS.n4384 VSS.n4279 0.0353837
R38173 VSS.n4383 VSS.n4280 0.0353837
R38174 VSS.n4382 VSS.n4281 0.0353837
R38175 VSS.n4381 VSS.n4282 0.0353837
R38176 VSS.n4380 VSS.n4283 0.0353837
R38177 VSS.n4379 VSS.n4284 0.0353837
R38178 VSS.n4378 VSS.n4285 0.0353837
R38179 VSS.n4377 VSS.n4286 0.0353837
R38180 VSS.n4376 VSS.n4287 0.0353837
R38181 VSS.n4375 VSS.n4288 0.0353837
R38182 VSS.n4374 VSS.n4289 0.0353837
R38183 VSS.n4373 VSS.n4290 0.0353837
R38184 VSS.n4372 VSS.n4291 0.0353837
R38185 VSS.n4371 VSS.n4292 0.0353837
R38186 VSS.n4370 VSS.n4293 0.0353837
R38187 VSS.n4369 VSS.n4294 0.0353837
R38188 VSS.n4368 VSS.n4295 0.0353837
R38189 VSS.n4367 VSS.n4296 0.0353837
R38190 VSS.n4366 VSS.n4297 0.0353837
R38191 VSS.n4365 VSS.n4298 0.0353837
R38192 VSS.n4364 VSS.n4299 0.0353837
R38193 VSS.n4363 VSS.n4300 0.0353837
R38194 VSS.n4362 VSS.n4301 0.0353837
R38195 VSS.n4361 VSS.n4302 0.0353837
R38196 VSS.n4360 VSS.n4303 0.0353837
R38197 VSS.n4359 VSS.n4304 0.0353837
R38198 VSS.n4358 VSS.n4305 0.0353837
R38199 VSS.n4357 VSS.n4306 0.0353837
R38200 VSS.n4356 VSS.n4307 0.0353837
R38201 VSS.n4355 VSS.n4308 0.0353837
R38202 VSS.n4354 VSS.n4309 0.0353837
R38203 VSS.n4353 VSS.n4310 0.0353837
R38204 VSS.n4352 VSS.n4311 0.0353837
R38205 VSS.n4351 VSS.n4312 0.0353837
R38206 VSS.n4350 VSS.n4313 0.0353837
R38207 VSS.n4349 VSS.n4314 0.0353837
R38208 VSS.n4348 VSS.n4315 0.0353837
R38209 VSS.n4347 VSS.n4316 0.0353837
R38210 VSS.n4346 VSS.n4317 0.0353837
R38211 VSS.n4345 VSS.n4318 0.0353837
R38212 VSS.n4344 VSS.n4319 0.0353837
R38213 VSS.n4343 VSS.n4320 0.0353837
R38214 VSS.n4342 VSS.n4321 0.0353837
R38215 VSS.n4341 VSS.n4322 0.0353837
R38216 VSS.n4340 VSS.n4323 0.0353837
R38217 VSS.n4339 VSS.n4324 0.0353837
R38218 VSS.n4338 VSS.n4325 0.0353837
R38219 VSS.n4337 VSS.n4326 0.0353837
R38220 VSS.n4336 VSS.n4327 0.0353837
R38221 VSS.n4335 VSS.n4328 0.0353837
R38222 VSS.n4334 VSS.n4329 0.0353837
R38223 VSS.n4333 VSS.n4330 0.0353837
R38224 VSS.n4332 VSS.n4331 0.0353837
R38225 VSS.n2 VSS.n0 0.0353837
R38226 VSS.n4508 VSS.n4507 0.0353837
R38227 VSS.n3 VSS.n1 0.0353837
R38228 VSS.n4438 VSS.n4437 0.0353837
R38229 VSS.n4440 VSS.n4439 0.0353837
R38230 VSS.n4441 VSS.n4436 0.0353837
R38231 VSS.n4443 VSS.n4442 0.0353837
R38232 VSS.n4444 VSS.n4435 0.0353837
R38233 VSS.n4446 VSS.n4445 0.0353837
R38234 VSS.n4447 VSS.n4434 0.0353837
R38235 VSS.n4449 VSS.n4448 0.0353837
R38236 VSS.n4450 VSS.n4433 0.0353837
R38237 VSS.n4452 VSS.n4451 0.0353837
R38238 VSS.n4453 VSS.n4432 0.0353837
R38239 VSS.n4455 VSS.n4454 0.0353837
R38240 VSS.n4456 VSS.n4431 0.0353837
R38241 VSS.n4458 VSS.n4457 0.0353837
R38242 VSS.n4459 VSS.n4430 0.0353837
R38243 VSS.n4461 VSS.n4460 0.0353837
R38244 VSS.n4462 VSS.n4429 0.0353837
R38245 VSS.n4464 VSS.n4463 0.0353837
R38246 VSS.n4465 VSS.n4428 0.0353837
R38247 VSS.n4467 VSS.n4466 0.0353837
R38248 VSS.n4468 VSS.n4427 0.0353837
R38249 VSS.n4470 VSS.n4469 0.0353837
R38250 VSS.n4471 VSS.n4426 0.0353837
R38251 VSS.n4473 VSS.n4472 0.0353837
R38252 VSS.n4474 VSS.n4425 0.0353837
R38253 VSS.n4476 VSS.n4475 0.0353837
R38254 VSS.n4477 VSS.n4424 0.0353837
R38255 VSS.n4479 VSS.n4478 0.0353837
R38256 VSS.n4480 VSS.n4423 0.0353837
R38257 VSS.n4482 VSS.n4481 0.0353837
R38258 VSS.n4483 VSS.n4422 0.0353837
R38259 VSS.n4485 VSS.n4484 0.0353837
R38260 VSS.n4486 VSS.n4421 0.0353837
R38261 VSS.n4488 VSS.n4487 0.0353837
R38262 VSS.n4489 VSS.n4420 0.0353837
R38263 VSS.n4491 VSS.n4490 0.0353837
R38264 VSS.n4492 VSS.n4419 0.0353837
R38265 VSS.n4494 VSS.n4493 0.0353837
R38266 VSS.n4495 VSS.n4418 0.0353837
R38267 VSS.n4497 VSS.n4496 0.0353837
R38268 VSS.n4498 VSS.n4417 0.0353837
R38269 VSS.n4501 VSS.n4499 0.0353837
R38270 VSS.n4252 VSS.n193 0.0353837
R38271 VSS.n4411 VSS.n195 0.0353837
R38272 VSS.n4410 VSS.n192 0.0353837
R38273 VSS.n4409 VSS.n196 0.0353837
R38274 VSS.n4408 VSS.n191 0.0353837
R38275 VSS.n4407 VSS.n197 0.0353837
R38276 VSS.n4406 VSS.n190 0.0353837
R38277 VSS.n4405 VSS.n198 0.0353837
R38278 VSS.n4404 VSS.n189 0.0353837
R38279 VSS.n4403 VSS.n199 0.0353837
R38280 VSS.n4402 VSS.n188 0.0353837
R38281 VSS.n4401 VSS.n200 0.0353837
R38282 VSS.n4400 VSS.n187 0.0353837
R38283 VSS.n4399 VSS.n201 0.0353837
R38284 VSS.n4398 VSS.n186 0.0353837
R38285 VSS.n4397 VSS.n202 0.0353837
R38286 VSS.n4396 VSS.n185 0.0353837
R38287 VSS.n4395 VSS.n203 0.0353837
R38288 VSS.n4394 VSS.n184 0.0353837
R38289 VSS.n4393 VSS.n204 0.0353837
R38290 VSS.n4392 VSS.n183 0.0353837
R38291 VSS.n4391 VSS.n205 0.0353837
R38292 VSS.n4390 VSS.n182 0.0353837
R38293 VSS.n4389 VSS.n206 0.0353837
R38294 VSS.n4388 VSS.n181 0.0353837
R38295 VSS.n4387 VSS.n207 0.0353837
R38296 VSS.n4386 VSS.n180 0.0353837
R38297 VSS.n4385 VSS.n208 0.0353837
R38298 VSS.n4384 VSS.n179 0.0353837
R38299 VSS.n4383 VSS.n209 0.0353837
R38300 VSS.n4382 VSS.n178 0.0353837
R38301 VSS.n4381 VSS.n210 0.0353837
R38302 VSS.n4380 VSS.n177 0.0353837
R38303 VSS.n4379 VSS.n211 0.0353837
R38304 VSS.n4378 VSS.n176 0.0353837
R38305 VSS.n4377 VSS.n212 0.0353837
R38306 VSS.n4376 VSS.n175 0.0353837
R38307 VSS.n4375 VSS.n213 0.0353837
R38308 VSS.n4374 VSS.n174 0.0353837
R38309 VSS.n4373 VSS.n214 0.0353837
R38310 VSS.n4372 VSS.n173 0.0353837
R38311 VSS.n4371 VSS.n215 0.0353837
R38312 VSS.n4370 VSS.n172 0.0353837
R38313 VSS.n4369 VSS.n216 0.0353837
R38314 VSS.n4368 VSS.n171 0.0353837
R38315 VSS.n4367 VSS.n217 0.0353837
R38316 VSS.n4366 VSS.n170 0.0353837
R38317 VSS.n4365 VSS.n218 0.0353837
R38318 VSS.n4364 VSS.n169 0.0353837
R38319 VSS.n4363 VSS.n219 0.0353837
R38320 VSS.n4362 VSS.n168 0.0353837
R38321 VSS.n4361 VSS.n220 0.0353837
R38322 VSS.n4360 VSS.n167 0.0353837
R38323 VSS.n4359 VSS.n221 0.0353837
R38324 VSS.n4358 VSS.n166 0.0353837
R38325 VSS.n4357 VSS.n222 0.0353837
R38326 VSS.n4356 VSS.n165 0.0353837
R38327 VSS.n4355 VSS.n223 0.0353837
R38328 VSS.n4354 VSS.n164 0.0353837
R38329 VSS.n4353 VSS.n224 0.0353837
R38330 VSS.n4352 VSS.n163 0.0353837
R38331 VSS.n4351 VSS.n225 0.0353837
R38332 VSS.n4350 VSS.n162 0.0353837
R38333 VSS.n4349 VSS.n226 0.0353837
R38334 VSS.n4348 VSS.n161 0.0353837
R38335 VSS.n4347 VSS.n227 0.0353837
R38336 VSS.n4346 VSS.n160 0.0353837
R38337 VSS.n4345 VSS.n228 0.0353837
R38338 VSS.n4344 VSS.n159 0.0353837
R38339 VSS.n4343 VSS.n229 0.0353837
R38340 VSS.n4342 VSS.n158 0.0353837
R38341 VSS.n4341 VSS.n230 0.0353837
R38342 VSS.n4340 VSS.n157 0.0353837
R38343 VSS.n4339 VSS.n231 0.0353837
R38344 VSS.n4338 VSS.n156 0.0353837
R38345 VSS.n4337 VSS.n232 0.0353837
R38346 VSS.n4336 VSS.n155 0.0353837
R38347 VSS.n4335 VSS.n233 0.0353837
R38348 VSS.n4334 VSS.n154 0.0353837
R38349 VSS.n4333 VSS.n234 0.0353837
R38350 VSS.n4332 VSS.n153 0.0353837
R38351 VSS.n235 VSS.n2 0.0353837
R38352 VSS.n4507 VSS.n4506 0.0353837
R38353 VSS.n236 VSS.n3 0.0353837
R38354 VSS.n4437 VSS.n152 0.0353837
R38355 VSS.n4440 VSS.n237 0.0353837
R38356 VSS.n4441 VSS.n151 0.0353837
R38357 VSS.n4442 VSS.n238 0.0353837
R38358 VSS.n4435 VSS.n150 0.0353837
R38359 VSS.n4446 VSS.n239 0.0353837
R38360 VSS.n4447 VSS.n149 0.0353837
R38361 VSS.n4448 VSS.n240 0.0353837
R38362 VSS.n4433 VSS.n148 0.0353837
R38363 VSS.n4452 VSS.n241 0.0353837
R38364 VSS.n4453 VSS.n147 0.0353837
R38365 VSS.n4454 VSS.n242 0.0353837
R38366 VSS.n4431 VSS.n146 0.0353837
R38367 VSS.n4458 VSS.n243 0.0353837
R38368 VSS.n4459 VSS.n145 0.0353837
R38369 VSS.n4460 VSS.n244 0.0353837
R38370 VSS.n4429 VSS.n144 0.0353837
R38371 VSS.n4464 VSS.n245 0.0353837
R38372 VSS.n4465 VSS.n143 0.0353837
R38373 VSS.n4466 VSS.n246 0.0353837
R38374 VSS.n4427 VSS.n142 0.0353837
R38375 VSS.n4470 VSS.n247 0.0353837
R38376 VSS.n4471 VSS.n141 0.0353837
R38377 VSS.n4472 VSS.n248 0.0353837
R38378 VSS.n4425 VSS.n140 0.0353837
R38379 VSS.n4476 VSS.n249 0.0353837
R38380 VSS.n4477 VSS.n139 0.0353837
R38381 VSS.n4478 VSS.n250 0.0353837
R38382 VSS.n4423 VSS.n138 0.0353837
R38383 VSS.n4482 VSS.n251 0.0353837
R38384 VSS.n4483 VSS.n137 0.0353837
R38385 VSS.n4484 VSS.n252 0.0353837
R38386 VSS.n4421 VSS.n136 0.0353837
R38387 VSS.n4488 VSS.n253 0.0353837
R38388 VSS.n4489 VSS.n135 0.0353837
R38389 VSS.n4490 VSS.n254 0.0353837
R38390 VSS.n4419 VSS.n134 0.0353837
R38391 VSS.n4494 VSS.n255 0.0353837
R38392 VSS.n4495 VSS.n133 0.0353837
R38393 VSS.n4496 VSS.n256 0.0353837
R38394 VSS.n4417 VSS.n132 0.0353837
R38395 VSS.n4502 VSS.n4501 0.0353837
R38396 VSS.n4500 VSS.n321 0.0353837
R38397 VSS.n2480 VSS.n2351 0.0353837
R38398 VSS.n3048 VSS.n2483 0.0353837
R38399 VSS.n3047 VSS.n2484 0.0353837
R38400 VSS.n3046 VSS.n2486 0.0353837
R38401 VSS.n2489 VSS.n2487 0.0353837
R38402 VSS.n3042 VSS.n2491 0.0353837
R38403 VSS.n3041 VSS.n2492 0.0353837
R38404 VSS.n3040 VSS.n2494 0.0353837
R38405 VSS.n2497 VSS.n2495 0.0353837
R38406 VSS.n3036 VSS.n2499 0.0353837
R38407 VSS.n3035 VSS.n2500 0.0353837
R38408 VSS.n3034 VSS.n2502 0.0353837
R38409 VSS.n2505 VSS.n2503 0.0353837
R38410 VSS.n3030 VSS.n2507 0.0353837
R38411 VSS.n3029 VSS.n2508 0.0353837
R38412 VSS.n3028 VSS.n2510 0.0353837
R38413 VSS.n2513 VSS.n2511 0.0353837
R38414 VSS.n3024 VSS.n2515 0.0353837
R38415 VSS.n3023 VSS.n2516 0.0353837
R38416 VSS.n3022 VSS.n2518 0.0353837
R38417 VSS.n2521 VSS.n2519 0.0353837
R38418 VSS.n3018 VSS.n2523 0.0353837
R38419 VSS.n3017 VSS.n2524 0.0353837
R38420 VSS.n3016 VSS.n2526 0.0353837
R38421 VSS.n2529 VSS.n2527 0.0353837
R38422 VSS.n3012 VSS.n2531 0.0353837
R38423 VSS.n3011 VSS.n2532 0.0353837
R38424 VSS.n3010 VSS.n2534 0.0353837
R38425 VSS.n2537 VSS.n2535 0.0353837
R38426 VSS.n3006 VSS.n2539 0.0353837
R38427 VSS.n3005 VSS.n2540 0.0353837
R38428 VSS.n3004 VSS.n2542 0.0353837
R38429 VSS.n2545 VSS.n2543 0.0353837
R38430 VSS.n3000 VSS.n2547 0.0353837
R38431 VSS.n2999 VSS.n2548 0.0353837
R38432 VSS.n2998 VSS.n2550 0.0353837
R38433 VSS.n2553 VSS.n2551 0.0353837
R38434 VSS.n2994 VSS.n2555 0.0353837
R38435 VSS.n2993 VSS.n2556 0.0353837
R38436 VSS.n2992 VSS.n2558 0.0353837
R38437 VSS.n2561 VSS.n2559 0.0353837
R38438 VSS.n2988 VSS.n2563 0.0353837
R38439 VSS.n2987 VSS.n2564 0.0353837
R38440 VSS.n2986 VSS.n2566 0.0353837
R38441 VSS.n2569 VSS.n2567 0.0353837
R38442 VSS.n2982 VSS.n2571 0.0353837
R38443 VSS.n2981 VSS.n2572 0.0353837
R38444 VSS.n2980 VSS.n2574 0.0353837
R38445 VSS.n2577 VSS.n2575 0.0353837
R38446 VSS.n2976 VSS.n2579 0.0353837
R38447 VSS.n2975 VSS.n2580 0.0353837
R38448 VSS.n2974 VSS.n2582 0.0353837
R38449 VSS.n2585 VSS.n2583 0.0353837
R38450 VSS.n2970 VSS.n2587 0.0353837
R38451 VSS.n2969 VSS.n2588 0.0353837
R38452 VSS.n2968 VSS.n2590 0.0353837
R38453 VSS.n2593 VSS.n2591 0.0353837
R38454 VSS.n2964 VSS.n2595 0.0353837
R38455 VSS.n2963 VSS.n2596 0.0353837
R38456 VSS.n2962 VSS.n2598 0.0353837
R38457 VSS.n2601 VSS.n2599 0.0353837
R38458 VSS.n2958 VSS.n2603 0.0353837
R38459 VSS.n2957 VSS.n2604 0.0353837
R38460 VSS.n2956 VSS.n2606 0.0353837
R38461 VSS.n2609 VSS.n2607 0.0353837
R38462 VSS.n2952 VSS.n2611 0.0353837
R38463 VSS.n2951 VSS.n2612 0.0353837
R38464 VSS.n2950 VSS.n2614 0.0353837
R38465 VSS.n2617 VSS.n2615 0.0353837
R38466 VSS.n2946 VSS.n2619 0.0353837
R38467 VSS.n2945 VSS.n2620 0.0353837
R38468 VSS.n2944 VSS.n2622 0.0353837
R38469 VSS.n2625 VSS.n2623 0.0353837
R38470 VSS.n2940 VSS.n2627 0.0353837
R38471 VSS.n2939 VSS.n2628 0.0353837
R38472 VSS.n2938 VSS.n2630 0.0353837
R38473 VSS.n2633 VSS.n2631 0.0353837
R38474 VSS.n2934 VSS.n2635 0.0353837
R38475 VSS.n2933 VSS.n2636 0.0353837
R38476 VSS.n2932 VSS.n2638 0.0353837
R38477 VSS.n2640 VSS.n2639 0.0353837
R38478 VSS.n2928 VSS.n2642 0.0353837
R38479 VSS.n2927 VSS.n2643 0.0353837
R38480 VSS.n2646 VSS.n2645 0.0353837
R38481 VSS.n2923 VSS.n2648 0.0353837
R38482 VSS.n2922 VSS.n2650 0.0353837
R38483 VSS.n2921 VSS.n2651 0.0353837
R38484 VSS.n2654 VSS.n2653 0.0353837
R38485 VSS.n2917 VSS.n2656 0.0353837
R38486 VSS.n2916 VSS.n2658 0.0353837
R38487 VSS.n2915 VSS.n2659 0.0353837
R38488 VSS.n2662 VSS.n2661 0.0353837
R38489 VSS.n2911 VSS.n2664 0.0353837
R38490 VSS.n2910 VSS.n2666 0.0353837
R38491 VSS.n2909 VSS.n2667 0.0353837
R38492 VSS.n2670 VSS.n2669 0.0353837
R38493 VSS.n2905 VSS.n2672 0.0353837
R38494 VSS.n2904 VSS.n2674 0.0353837
R38495 VSS.n2903 VSS.n2675 0.0353837
R38496 VSS.n2678 VSS.n2677 0.0353837
R38497 VSS.n2899 VSS.n2680 0.0353837
R38498 VSS.n2898 VSS.n2682 0.0353837
R38499 VSS.n2897 VSS.n2683 0.0353837
R38500 VSS.n2686 VSS.n2685 0.0353837
R38501 VSS.n2893 VSS.n2688 0.0353837
R38502 VSS.n2892 VSS.n2690 0.0353837
R38503 VSS.n2891 VSS.n2691 0.0353837
R38504 VSS.n2694 VSS.n2693 0.0353837
R38505 VSS.n2887 VSS.n2696 0.0353837
R38506 VSS.n2886 VSS.n2698 0.0353837
R38507 VSS.n2885 VSS.n2699 0.0353837
R38508 VSS.n2702 VSS.n2701 0.0353837
R38509 VSS.n2881 VSS.n2704 0.0353837
R38510 VSS.n2880 VSS.n2706 0.0353837
R38511 VSS.n2879 VSS.n2707 0.0353837
R38512 VSS.n2710 VSS.n2709 0.0353837
R38513 VSS.n2875 VSS.n2712 0.0353837
R38514 VSS.n2874 VSS.n2714 0.0353837
R38515 VSS.n2873 VSS.n2715 0.0353837
R38516 VSS.n2718 VSS.n2717 0.0353837
R38517 VSS.n2869 VSS.n2720 0.0353837
R38518 VSS.n2868 VSS.n2722 0.0353837
R38519 VSS.n2867 VSS.n2723 0.0353837
R38520 VSS.n2726 VSS.n2725 0.0353837
R38521 VSS.n2863 VSS.n2791 0.0353837
R38522 VSS.n2862 VSS.n2793 0.0353837
R38523 VSS.n2861 VSS.n2858 0.0353837
R38524 VSS.n3049 VSS.n3048 0.0353837
R38525 VSS.n3047 VSS.n2481 0.0353837
R38526 VSS.n3046 VSS.n3045 0.0353837
R38527 VSS.n3044 VSS.n2487 0.0353837
R38528 VSS.n3043 VSS.n3042 0.0353837
R38529 VSS.n3041 VSS.n2488 0.0353837
R38530 VSS.n3040 VSS.n3039 0.0353837
R38531 VSS.n3038 VSS.n2495 0.0353837
R38532 VSS.n3037 VSS.n3036 0.0353837
R38533 VSS.n3035 VSS.n2496 0.0353837
R38534 VSS.n3034 VSS.n3033 0.0353837
R38535 VSS.n3032 VSS.n2503 0.0353837
R38536 VSS.n3031 VSS.n3030 0.0353837
R38537 VSS.n3029 VSS.n2504 0.0353837
R38538 VSS.n3028 VSS.n3027 0.0353837
R38539 VSS.n3026 VSS.n2511 0.0353837
R38540 VSS.n3025 VSS.n3024 0.0353837
R38541 VSS.n3023 VSS.n2512 0.0353837
R38542 VSS.n3022 VSS.n3021 0.0353837
R38543 VSS.n3020 VSS.n2519 0.0353837
R38544 VSS.n3019 VSS.n3018 0.0353837
R38545 VSS.n3017 VSS.n2520 0.0353837
R38546 VSS.n3016 VSS.n3015 0.0353837
R38547 VSS.n3014 VSS.n2527 0.0353837
R38548 VSS.n3013 VSS.n3012 0.0353837
R38549 VSS.n3011 VSS.n2528 0.0353837
R38550 VSS.n3010 VSS.n3009 0.0353837
R38551 VSS.n3008 VSS.n2535 0.0353837
R38552 VSS.n3007 VSS.n3006 0.0353837
R38553 VSS.n3005 VSS.n2536 0.0353837
R38554 VSS.n3004 VSS.n3003 0.0353837
R38555 VSS.n3002 VSS.n2543 0.0353837
R38556 VSS.n3001 VSS.n3000 0.0353837
R38557 VSS.n2999 VSS.n2544 0.0353837
R38558 VSS.n2998 VSS.n2997 0.0353837
R38559 VSS.n2996 VSS.n2551 0.0353837
R38560 VSS.n2995 VSS.n2994 0.0353837
R38561 VSS.n2993 VSS.n2552 0.0353837
R38562 VSS.n2992 VSS.n2991 0.0353837
R38563 VSS.n2990 VSS.n2559 0.0353837
R38564 VSS.n2989 VSS.n2988 0.0353837
R38565 VSS.n2987 VSS.n2560 0.0353837
R38566 VSS.n2986 VSS.n2985 0.0353837
R38567 VSS.n2984 VSS.n2567 0.0353837
R38568 VSS.n2983 VSS.n2982 0.0353837
R38569 VSS.n2981 VSS.n2568 0.0353837
R38570 VSS.n2980 VSS.n2979 0.0353837
R38571 VSS.n2978 VSS.n2575 0.0353837
R38572 VSS.n2977 VSS.n2976 0.0353837
R38573 VSS.n2975 VSS.n2576 0.0353837
R38574 VSS.n2974 VSS.n2973 0.0353837
R38575 VSS.n2972 VSS.n2583 0.0353837
R38576 VSS.n2971 VSS.n2970 0.0353837
R38577 VSS.n2969 VSS.n2584 0.0353837
R38578 VSS.n2968 VSS.n2967 0.0353837
R38579 VSS.n2966 VSS.n2591 0.0353837
R38580 VSS.n2965 VSS.n2964 0.0353837
R38581 VSS.n2963 VSS.n2592 0.0353837
R38582 VSS.n2962 VSS.n2961 0.0353837
R38583 VSS.n2960 VSS.n2599 0.0353837
R38584 VSS.n2959 VSS.n2958 0.0353837
R38585 VSS.n2957 VSS.n2600 0.0353837
R38586 VSS.n2956 VSS.n2955 0.0353837
R38587 VSS.n2954 VSS.n2607 0.0353837
R38588 VSS.n2953 VSS.n2952 0.0353837
R38589 VSS.n2951 VSS.n2608 0.0353837
R38590 VSS.n2950 VSS.n2949 0.0353837
R38591 VSS.n2948 VSS.n2615 0.0353837
R38592 VSS.n2947 VSS.n2946 0.0353837
R38593 VSS.n2945 VSS.n2616 0.0353837
R38594 VSS.n2944 VSS.n2943 0.0353837
R38595 VSS.n2942 VSS.n2623 0.0353837
R38596 VSS.n2941 VSS.n2940 0.0353837
R38597 VSS.n2939 VSS.n2624 0.0353837
R38598 VSS.n2938 VSS.n2937 0.0353837
R38599 VSS.n2936 VSS.n2631 0.0353837
R38600 VSS.n2935 VSS.n2934 0.0353837
R38601 VSS.n2933 VSS.n2632 0.0353837
R38602 VSS.n2932 VSS.n2931 0.0353837
R38603 VSS.n2930 VSS.n2639 0.0353837
R38604 VSS.n2929 VSS.n2928 0.0353837
R38605 VSS.n2927 VSS.n2926 0.0353837
R38606 VSS.n2925 VSS.n2646 0.0353837
R38607 VSS.n2924 VSS.n2923 0.0353837
R38608 VSS.n2922 VSS.n2647 0.0353837
R38609 VSS.n2921 VSS.n2920 0.0353837
R38610 VSS.n2919 VSS.n2654 0.0353837
R38611 VSS.n2918 VSS.n2917 0.0353837
R38612 VSS.n2916 VSS.n2655 0.0353837
R38613 VSS.n2915 VSS.n2914 0.0353837
R38614 VSS.n2913 VSS.n2662 0.0353837
R38615 VSS.n2912 VSS.n2911 0.0353837
R38616 VSS.n2910 VSS.n2663 0.0353837
R38617 VSS.n2909 VSS.n2908 0.0353837
R38618 VSS.n2907 VSS.n2670 0.0353837
R38619 VSS.n2906 VSS.n2905 0.0353837
R38620 VSS.n2904 VSS.n2671 0.0353837
R38621 VSS.n2903 VSS.n2902 0.0353837
R38622 VSS.n2901 VSS.n2678 0.0353837
R38623 VSS.n2900 VSS.n2899 0.0353837
R38624 VSS.n2898 VSS.n2679 0.0353837
R38625 VSS.n2897 VSS.n2896 0.0353837
R38626 VSS.n2895 VSS.n2686 0.0353837
R38627 VSS.n2894 VSS.n2893 0.0353837
R38628 VSS.n2892 VSS.n2687 0.0353837
R38629 VSS.n2891 VSS.n2890 0.0353837
R38630 VSS.n2889 VSS.n2694 0.0353837
R38631 VSS.n2888 VSS.n2887 0.0353837
R38632 VSS.n2886 VSS.n2695 0.0353837
R38633 VSS.n2885 VSS.n2884 0.0353837
R38634 VSS.n2883 VSS.n2702 0.0353837
R38635 VSS.n2882 VSS.n2881 0.0353837
R38636 VSS.n2880 VSS.n2703 0.0353837
R38637 VSS.n2879 VSS.n2878 0.0353837
R38638 VSS.n2877 VSS.n2710 0.0353837
R38639 VSS.n2876 VSS.n2875 0.0353837
R38640 VSS.n2874 VSS.n2711 0.0353837
R38641 VSS.n2873 VSS.n2872 0.0353837
R38642 VSS.n2871 VSS.n2718 0.0353837
R38643 VSS.n2870 VSS.n2869 0.0353837
R38644 VSS.n2868 VSS.n2719 0.0353837
R38645 VSS.n2867 VSS.n2866 0.0353837
R38646 VSS.n2865 VSS.n2726 0.0353837
R38647 VSS.n2864 VSS.n2863 0.0353837
R38648 VSS.n2862 VSS.n2727 0.0353837
R38649 VSS.n892 VSS.n758 0.0348421
R38650 VSS.n4034 VSS.n604 0.0336579
R38651 VSS.n676 VSS.n675 0.0336579
R38652 VSS.n4027 VSS.n709 0.0283884
R38653 VSS.n3802 VSS.n708 0.0283884
R38654 VSS.n3508 VSS.n3507 0.0283884
R38655 VSS.n1755 VSS.n1754 0.0283884
R38656 VSS.n2098 VSS.n1620 0.0283884
R38657 VSS.n4180 VSS.n4179 0.0267963
R38658 VSS.n1831 VSS.n1830 0.023
R38659 VSS.n2175 VSS.n2174 0.023
R38660 VSS.n1790 VSS.n1789 0.023
R38661 VSS.n3536 VSS.n3535 0.023
R38662 VSS.n738 VSS.n717 0.023
R38663 VSS.n4132 VSS.n4131 0.023
R38664 VSS.n1354 VSS.n1139 0.023
R38665 VSS.n3170 VSS.n3169 0.023
R38666 VSS.n3181 VSS.n3180 0.023
R38667 VSS.n3319 VSS.n3318 0.023
R38668 VSS.n4188 VSS.n4187 0.023
R38669 VSS.n3786 VSS.n3785 0.023
R38670 VSS.n3054 VSS.n2286 0.023
R38671 VSS.n3050 VSS.n3049 0.0188524
R38672 VSS.n4413 VSS.n4412 0.0188497
R38673 VSS.n4499 VSS.n384 0.0188497
R38674 VSS.n2860 VSS.n2727 0.0188497
R38675 VSS.n3997 VSS.n3896 0.0182632
R38676 VSS.n703 VSS.n702 0.0170789
R38677 VSS.n2129 VSS.n2128 0.0135263
R38678 VSS.n1912 VSS.n1867 0.0135263
R38679 VSS.n1761 VSS.n1759 0.0111579
R38680 VSS.n4181 VSS.n456 0.0100192
R38681 VSS.n1700 VSS.n783 0.00878947
R38682 VSS.n3793 VSS.n3561 0.00608621
R38683 VSS.n3387 VSS.n3386 0.00459091
R38684 VSS.n4188 VSS.n447 0.0041
R38685 VSS.n3055 VSS.n3054 0.0041
R38686 VSS.n2185 VSS.n1655 0.00223758
R38687 VSS.n2126 VSS.n1620 0.00223758
R38688 VSS.n4146 VSS.n4145 0.00223758
R38689 VSS.n615 VSS.n457 0.00223758
R38690 VSS.n3423 VSS.n3422 0.00223758
R38691 VSS.n2186 VSS.n2185 0.00223758
R38692 VSS.n3050 VSS.n2480 0.00158269
R38693 VSS.n4415 VSS.n4414 0.00134872
R38694 VSS.n382 VSS.n193 0.00134872
R38695 VSS.n446 VSS.n192 0.00134872
R38696 VSS.n381 VSS.n192 0.00134872
R38697 VSS.n445 VSS.n191 0.00134872
R38698 VSS.n380 VSS.n191 0.00134872
R38699 VSS.n444 VSS.n190 0.00134872
R38700 VSS.n379 VSS.n190 0.00134872
R38701 VSS.n443 VSS.n189 0.00134872
R38702 VSS.n378 VSS.n189 0.00134872
R38703 VSS.n442 VSS.n188 0.00134872
R38704 VSS.n377 VSS.n188 0.00134872
R38705 VSS.n441 VSS.n187 0.00134872
R38706 VSS.n376 VSS.n187 0.00134872
R38707 VSS.n440 VSS.n186 0.00134872
R38708 VSS.n375 VSS.n186 0.00134872
R38709 VSS.n439 VSS.n185 0.00134872
R38710 VSS.n374 VSS.n185 0.00134872
R38711 VSS.n438 VSS.n184 0.00134872
R38712 VSS.n373 VSS.n184 0.00134872
R38713 VSS.n437 VSS.n183 0.00134872
R38714 VSS.n372 VSS.n183 0.00134872
R38715 VSS.n436 VSS.n182 0.00134872
R38716 VSS.n371 VSS.n182 0.00134872
R38717 VSS.n435 VSS.n181 0.00134872
R38718 VSS.n370 VSS.n181 0.00134872
R38719 VSS.n434 VSS.n180 0.00134872
R38720 VSS.n369 VSS.n180 0.00134872
R38721 VSS.n433 VSS.n179 0.00134872
R38722 VSS.n368 VSS.n179 0.00134872
R38723 VSS.n432 VSS.n178 0.00134872
R38724 VSS.n367 VSS.n178 0.00134872
R38725 VSS.n431 VSS.n177 0.00134872
R38726 VSS.n366 VSS.n177 0.00134872
R38727 VSS.n430 VSS.n176 0.00134872
R38728 VSS.n365 VSS.n176 0.00134872
R38729 VSS.n429 VSS.n175 0.00134872
R38730 VSS.n364 VSS.n175 0.00134872
R38731 VSS.n428 VSS.n174 0.00134872
R38732 VSS.n363 VSS.n174 0.00134872
R38733 VSS.n427 VSS.n173 0.00134872
R38734 VSS.n362 VSS.n173 0.00134872
R38735 VSS.n426 VSS.n172 0.00134872
R38736 VSS.n361 VSS.n172 0.00134872
R38737 VSS.n425 VSS.n171 0.00134872
R38738 VSS.n360 VSS.n171 0.00134872
R38739 VSS.n424 VSS.n170 0.00134872
R38740 VSS.n359 VSS.n170 0.00134872
R38741 VSS.n423 VSS.n169 0.00134872
R38742 VSS.n358 VSS.n169 0.00134872
R38743 VSS.n422 VSS.n168 0.00134872
R38744 VSS.n357 VSS.n168 0.00134872
R38745 VSS.n421 VSS.n167 0.00134872
R38746 VSS.n356 VSS.n167 0.00134872
R38747 VSS.n420 VSS.n166 0.00134872
R38748 VSS.n355 VSS.n166 0.00134872
R38749 VSS.n419 VSS.n165 0.00134872
R38750 VSS.n354 VSS.n165 0.00134872
R38751 VSS.n418 VSS.n164 0.00134872
R38752 VSS.n353 VSS.n164 0.00134872
R38753 VSS.n417 VSS.n163 0.00134872
R38754 VSS.n352 VSS.n163 0.00134872
R38755 VSS.n416 VSS.n162 0.00134872
R38756 VSS.n351 VSS.n162 0.00134872
R38757 VSS.n415 VSS.n161 0.00134872
R38758 VSS.n350 VSS.n161 0.00134872
R38759 VSS.n414 VSS.n160 0.00134872
R38760 VSS.n349 VSS.n160 0.00134872
R38761 VSS.n413 VSS.n159 0.00134872
R38762 VSS.n348 VSS.n159 0.00134872
R38763 VSS.n412 VSS.n158 0.00134872
R38764 VSS.n347 VSS.n158 0.00134872
R38765 VSS.n411 VSS.n157 0.00134872
R38766 VSS.n346 VSS.n157 0.00134872
R38767 VSS.n410 VSS.n156 0.00134872
R38768 VSS.n345 VSS.n156 0.00134872
R38769 VSS.n409 VSS.n155 0.00134872
R38770 VSS.n344 VSS.n155 0.00134872
R38771 VSS.n408 VSS.n154 0.00134872
R38772 VSS.n343 VSS.n154 0.00134872
R38773 VSS.n407 VSS.n153 0.00134872
R38774 VSS.n342 VSS.n153 0.00134872
R38775 VSS.n4506 VSS.n4 0.00134872
R38776 VSS.n4506 VSS.n68 0.00134872
R38777 VSS.n406 VSS.n152 0.00134872
R38778 VSS.n341 VSS.n152 0.00134872
R38779 VSS.n405 VSS.n151 0.00134872
R38780 VSS.n340 VSS.n151 0.00134872
R38781 VSS.n404 VSS.n150 0.00134872
R38782 VSS.n339 VSS.n150 0.00134872
R38783 VSS.n403 VSS.n149 0.00134872
R38784 VSS.n338 VSS.n149 0.00134872
R38785 VSS.n402 VSS.n148 0.00134872
R38786 VSS.n337 VSS.n148 0.00134872
R38787 VSS.n401 VSS.n147 0.00134872
R38788 VSS.n336 VSS.n147 0.00134872
R38789 VSS.n400 VSS.n146 0.00134872
R38790 VSS.n335 VSS.n146 0.00134872
R38791 VSS.n399 VSS.n145 0.00134872
R38792 VSS.n334 VSS.n145 0.00134872
R38793 VSS.n398 VSS.n144 0.00134872
R38794 VSS.n333 VSS.n144 0.00134872
R38795 VSS.n397 VSS.n143 0.00134872
R38796 VSS.n332 VSS.n143 0.00134872
R38797 VSS.n396 VSS.n142 0.00134872
R38798 VSS.n331 VSS.n142 0.00134872
R38799 VSS.n395 VSS.n141 0.00134872
R38800 VSS.n330 VSS.n141 0.00134872
R38801 VSS.n394 VSS.n140 0.00134872
R38802 VSS.n329 VSS.n140 0.00134872
R38803 VSS.n393 VSS.n139 0.00134872
R38804 VSS.n328 VSS.n139 0.00134872
R38805 VSS.n392 VSS.n138 0.00134872
R38806 VSS.n327 VSS.n138 0.00134872
R38807 VSS.n391 VSS.n137 0.00134872
R38808 VSS.n326 VSS.n137 0.00134872
R38809 VSS.n390 VSS.n136 0.00134872
R38810 VSS.n325 VSS.n136 0.00134872
R38811 VSS.n389 VSS.n135 0.00134872
R38812 VSS.n324 VSS.n135 0.00134872
R38813 VSS.n388 VSS.n134 0.00134872
R38814 VSS.n323 VSS.n134 0.00134872
R38815 VSS.n387 VSS.n133 0.00134872
R38816 VSS.n322 VSS.n133 0.00134872
R38817 VSS.n386 VSS.n132 0.00134872
R38818 VSS.n4416 VSS.n132 0.00134872
R38819 VSS.n4502 VSS.n257 0.00134872
R38820 VSS.n4505 VSS.n194 0.00134872
R38821 VSS.n320 VSS.n131 0.00134872
R38822 VSS.n4189 VSS.n131 0.00134872
R38823 VSS.n319 VSS.n130 0.00134872
R38824 VSS.n4190 VSS.n130 0.00134872
R38825 VSS.n318 VSS.n129 0.00134872
R38826 VSS.n4191 VSS.n129 0.00134872
R38827 VSS.n317 VSS.n128 0.00134872
R38828 VSS.n4192 VSS.n128 0.00134872
R38829 VSS.n316 VSS.n127 0.00134872
R38830 VSS.n4193 VSS.n127 0.00134872
R38831 VSS.n315 VSS.n126 0.00134872
R38832 VSS.n4194 VSS.n126 0.00134872
R38833 VSS.n314 VSS.n125 0.00134872
R38834 VSS.n4195 VSS.n125 0.00134872
R38835 VSS.n313 VSS.n124 0.00134872
R38836 VSS.n4196 VSS.n124 0.00134872
R38837 VSS.n312 VSS.n123 0.00134872
R38838 VSS.n4197 VSS.n123 0.00134872
R38839 VSS.n311 VSS.n122 0.00134872
R38840 VSS.n4198 VSS.n122 0.00134872
R38841 VSS.n310 VSS.n121 0.00134872
R38842 VSS.n4199 VSS.n121 0.00134872
R38843 VSS.n309 VSS.n120 0.00134872
R38844 VSS.n4200 VSS.n120 0.00134872
R38845 VSS.n308 VSS.n119 0.00134872
R38846 VSS.n4201 VSS.n119 0.00134872
R38847 VSS.n307 VSS.n118 0.00134872
R38848 VSS.n4202 VSS.n118 0.00134872
R38849 VSS.n306 VSS.n117 0.00134872
R38850 VSS.n4203 VSS.n117 0.00134872
R38851 VSS.n305 VSS.n116 0.00134872
R38852 VSS.n4204 VSS.n116 0.00134872
R38853 VSS.n304 VSS.n115 0.00134872
R38854 VSS.n4205 VSS.n115 0.00134872
R38855 VSS.n303 VSS.n114 0.00134872
R38856 VSS.n4206 VSS.n114 0.00134872
R38857 VSS.n302 VSS.n113 0.00134872
R38858 VSS.n4207 VSS.n113 0.00134872
R38859 VSS.n301 VSS.n112 0.00134872
R38860 VSS.n4208 VSS.n112 0.00134872
R38861 VSS.n300 VSS.n111 0.00134872
R38862 VSS.n4209 VSS.n111 0.00134872
R38863 VSS.n299 VSS.n110 0.00134872
R38864 VSS.n4210 VSS.n110 0.00134872
R38865 VSS.n298 VSS.n109 0.00134872
R38866 VSS.n4211 VSS.n109 0.00134872
R38867 VSS.n297 VSS.n108 0.00134872
R38868 VSS.n4212 VSS.n108 0.00134872
R38869 VSS.n296 VSS.n107 0.00134872
R38870 VSS.n4213 VSS.n107 0.00134872
R38871 VSS.n295 VSS.n106 0.00134872
R38872 VSS.n4214 VSS.n106 0.00134872
R38873 VSS.n294 VSS.n105 0.00134872
R38874 VSS.n4215 VSS.n105 0.00134872
R38875 VSS.n293 VSS.n104 0.00134872
R38876 VSS.n4216 VSS.n104 0.00134872
R38877 VSS.n292 VSS.n103 0.00134872
R38878 VSS.n4217 VSS.n103 0.00134872
R38879 VSS.n291 VSS.n102 0.00134872
R38880 VSS.n4218 VSS.n102 0.00134872
R38881 VSS.n290 VSS.n101 0.00134872
R38882 VSS.n4219 VSS.n101 0.00134872
R38883 VSS.n289 VSS.n100 0.00134872
R38884 VSS.n4220 VSS.n100 0.00134872
R38885 VSS.n288 VSS.n99 0.00134872
R38886 VSS.n4221 VSS.n99 0.00134872
R38887 VSS.n287 VSS.n98 0.00134872
R38888 VSS.n4222 VSS.n98 0.00134872
R38889 VSS.n286 VSS.n97 0.00134872
R38890 VSS.n4223 VSS.n97 0.00134872
R38891 VSS.n285 VSS.n96 0.00134872
R38892 VSS.n4224 VSS.n96 0.00134872
R38893 VSS.n284 VSS.n95 0.00134872
R38894 VSS.n4225 VSS.n95 0.00134872
R38895 VSS.n283 VSS.n94 0.00134872
R38896 VSS.n4226 VSS.n94 0.00134872
R38897 VSS.n282 VSS.n93 0.00134872
R38898 VSS.n4227 VSS.n93 0.00134872
R38899 VSS.n281 VSS.n92 0.00134872
R38900 VSS.n4228 VSS.n92 0.00134872
R38901 VSS.n280 VSS.n91 0.00134872
R38902 VSS.n4229 VSS.n91 0.00134872
R38903 VSS.n279 VSS.n90 0.00134872
R38904 VSS.n4230 VSS.n90 0.00134872
R38905 VSS.n278 VSS.n89 0.00134872
R38906 VSS.n4231 VSS.n89 0.00134872
R38907 VSS.n277 VSS.n88 0.00134872
R38908 VSS.n4232 VSS.n88 0.00134872
R38909 VSS.n276 VSS.n87 0.00134872
R38910 VSS.n4233 VSS.n87 0.00134872
R38911 VSS.n275 VSS.n86 0.00134872
R38912 VSS.n4234 VSS.n86 0.00134872
R38913 VSS.n274 VSS.n85 0.00134872
R38914 VSS.n4235 VSS.n85 0.00134872
R38915 VSS.n273 VSS.n84 0.00134872
R38916 VSS.n4236 VSS.n84 0.00134872
R38917 VSS.n272 VSS.n83 0.00134872
R38918 VSS.n4237 VSS.n83 0.00134872
R38919 VSS.n271 VSS.n82 0.00134872
R38920 VSS.n4238 VSS.n82 0.00134872
R38921 VSS.n270 VSS.n81 0.00134872
R38922 VSS.n4239 VSS.n81 0.00134872
R38923 VSS.n269 VSS.n80 0.00134872
R38924 VSS.n4240 VSS.n80 0.00134872
R38925 VSS.n268 VSS.n79 0.00134872
R38926 VSS.n4241 VSS.n79 0.00134872
R38927 VSS.n267 VSS.n78 0.00134872
R38928 VSS.n4242 VSS.n78 0.00134872
R38929 VSS.n266 VSS.n77 0.00134872
R38930 VSS.n4243 VSS.n77 0.00134872
R38931 VSS.n265 VSS.n76 0.00134872
R38932 VSS.n4244 VSS.n76 0.00134872
R38933 VSS.n264 VSS.n75 0.00134872
R38934 VSS.n4245 VSS.n75 0.00134872
R38935 VSS.n263 VSS.n74 0.00134872
R38936 VSS.n4246 VSS.n74 0.00134872
R38937 VSS.n262 VSS.n73 0.00134872
R38938 VSS.n4247 VSS.n73 0.00134872
R38939 VSS.n261 VSS.n72 0.00134872
R38940 VSS.n4248 VSS.n72 0.00134872
R38941 VSS.n260 VSS.n71 0.00134872
R38942 VSS.n4249 VSS.n71 0.00134872
R38943 VSS.n259 VSS.n70 0.00134872
R38944 VSS.n4250 VSS.n70 0.00134872
R38945 VSS.n258 VSS.n69 0.00134872
R38946 VSS.n4251 VSS.n69 0.00134872
R38947 VSS.n4503 VSS.n385 0.00134872
R38948 VSS.n4415 VSS.n193 0.00134872
R38949 VSS.n446 VSS.n195 0.00134872
R38950 VSS.n445 VSS.n196 0.00134872
R38951 VSS.n444 VSS.n197 0.00134872
R38952 VSS.n443 VSS.n198 0.00134872
R38953 VSS.n442 VSS.n199 0.00134872
R38954 VSS.n441 VSS.n200 0.00134872
R38955 VSS.n440 VSS.n201 0.00134872
R38956 VSS.n439 VSS.n202 0.00134872
R38957 VSS.n438 VSS.n203 0.00134872
R38958 VSS.n437 VSS.n204 0.00134872
R38959 VSS.n436 VSS.n205 0.00134872
R38960 VSS.n435 VSS.n206 0.00134872
R38961 VSS.n434 VSS.n207 0.00134872
R38962 VSS.n433 VSS.n208 0.00134872
R38963 VSS.n432 VSS.n209 0.00134872
R38964 VSS.n431 VSS.n210 0.00134872
R38965 VSS.n430 VSS.n211 0.00134872
R38966 VSS.n429 VSS.n212 0.00134872
R38967 VSS.n428 VSS.n213 0.00134872
R38968 VSS.n427 VSS.n214 0.00134872
R38969 VSS.n426 VSS.n215 0.00134872
R38970 VSS.n425 VSS.n216 0.00134872
R38971 VSS.n424 VSS.n217 0.00134872
R38972 VSS.n423 VSS.n218 0.00134872
R38973 VSS.n422 VSS.n219 0.00134872
R38974 VSS.n421 VSS.n220 0.00134872
R38975 VSS.n420 VSS.n221 0.00134872
R38976 VSS.n419 VSS.n222 0.00134872
R38977 VSS.n418 VSS.n223 0.00134872
R38978 VSS.n417 VSS.n224 0.00134872
R38979 VSS.n416 VSS.n225 0.00134872
R38980 VSS.n415 VSS.n226 0.00134872
R38981 VSS.n414 VSS.n227 0.00134872
R38982 VSS.n413 VSS.n228 0.00134872
R38983 VSS.n412 VSS.n229 0.00134872
R38984 VSS.n411 VSS.n230 0.00134872
R38985 VSS.n410 VSS.n231 0.00134872
R38986 VSS.n409 VSS.n232 0.00134872
R38987 VSS.n408 VSS.n233 0.00134872
R38988 VSS.n407 VSS.n234 0.00134872
R38989 VSS.n235 VSS.n4 0.00134872
R38990 VSS.n406 VSS.n236 0.00134872
R38991 VSS.n405 VSS.n237 0.00134872
R38992 VSS.n404 VSS.n238 0.00134872
R38993 VSS.n403 VSS.n239 0.00134872
R38994 VSS.n402 VSS.n240 0.00134872
R38995 VSS.n401 VSS.n241 0.00134872
R38996 VSS.n400 VSS.n242 0.00134872
R38997 VSS.n399 VSS.n243 0.00134872
R38998 VSS.n398 VSS.n244 0.00134872
R38999 VSS.n397 VSS.n245 0.00134872
R39000 VSS.n396 VSS.n246 0.00134872
R39001 VSS.n395 VSS.n247 0.00134872
R39002 VSS.n394 VSS.n248 0.00134872
R39003 VSS.n393 VSS.n249 0.00134872
R39004 VSS.n392 VSS.n250 0.00134872
R39005 VSS.n391 VSS.n251 0.00134872
R39006 VSS.n390 VSS.n252 0.00134872
R39007 VSS.n389 VSS.n253 0.00134872
R39008 VSS.n388 VSS.n254 0.00134872
R39009 VSS.n387 VSS.n255 0.00134872
R39010 VSS.n386 VSS.n256 0.00134872
R39011 VSS.n4251 VSS.n383 0.00134872
R39012 VSS.n382 VSS.n195 0.00134872
R39013 VSS.n381 VSS.n196 0.00134872
R39014 VSS.n380 VSS.n197 0.00134872
R39015 VSS.n379 VSS.n198 0.00134872
R39016 VSS.n378 VSS.n199 0.00134872
R39017 VSS.n377 VSS.n200 0.00134872
R39018 VSS.n376 VSS.n201 0.00134872
R39019 VSS.n375 VSS.n202 0.00134872
R39020 VSS.n374 VSS.n203 0.00134872
R39021 VSS.n373 VSS.n204 0.00134872
R39022 VSS.n372 VSS.n205 0.00134872
R39023 VSS.n371 VSS.n206 0.00134872
R39024 VSS.n370 VSS.n207 0.00134872
R39025 VSS.n369 VSS.n208 0.00134872
R39026 VSS.n368 VSS.n209 0.00134872
R39027 VSS.n367 VSS.n210 0.00134872
R39028 VSS.n366 VSS.n211 0.00134872
R39029 VSS.n365 VSS.n212 0.00134872
R39030 VSS.n364 VSS.n213 0.00134872
R39031 VSS.n363 VSS.n214 0.00134872
R39032 VSS.n362 VSS.n215 0.00134872
R39033 VSS.n361 VSS.n216 0.00134872
R39034 VSS.n360 VSS.n217 0.00134872
R39035 VSS.n359 VSS.n218 0.00134872
R39036 VSS.n358 VSS.n219 0.00134872
R39037 VSS.n357 VSS.n220 0.00134872
R39038 VSS.n356 VSS.n221 0.00134872
R39039 VSS.n355 VSS.n222 0.00134872
R39040 VSS.n354 VSS.n223 0.00134872
R39041 VSS.n353 VSS.n224 0.00134872
R39042 VSS.n352 VSS.n225 0.00134872
R39043 VSS.n351 VSS.n226 0.00134872
R39044 VSS.n350 VSS.n227 0.00134872
R39045 VSS.n349 VSS.n228 0.00134872
R39046 VSS.n348 VSS.n229 0.00134872
R39047 VSS.n347 VSS.n230 0.00134872
R39048 VSS.n346 VSS.n231 0.00134872
R39049 VSS.n345 VSS.n232 0.00134872
R39050 VSS.n344 VSS.n233 0.00134872
R39051 VSS.n343 VSS.n234 0.00134872
R39052 VSS.n342 VSS.n235 0.00134872
R39053 VSS.n236 VSS.n68 0.00134872
R39054 VSS.n341 VSS.n237 0.00134872
R39055 VSS.n340 VSS.n238 0.00134872
R39056 VSS.n339 VSS.n239 0.00134872
R39057 VSS.n338 VSS.n240 0.00134872
R39058 VSS.n337 VSS.n241 0.00134872
R39059 VSS.n336 VSS.n242 0.00134872
R39060 VSS.n335 VSS.n243 0.00134872
R39061 VSS.n334 VSS.n244 0.00134872
R39062 VSS.n333 VSS.n245 0.00134872
R39063 VSS.n332 VSS.n246 0.00134872
R39064 VSS.n331 VSS.n247 0.00134872
R39065 VSS.n330 VSS.n248 0.00134872
R39066 VSS.n329 VSS.n249 0.00134872
R39067 VSS.n328 VSS.n250 0.00134872
R39068 VSS.n327 VSS.n251 0.00134872
R39069 VSS.n326 VSS.n252 0.00134872
R39070 VSS.n325 VSS.n253 0.00134872
R39071 VSS.n324 VSS.n254 0.00134872
R39072 VSS.n323 VSS.n255 0.00134872
R39073 VSS.n322 VSS.n256 0.00134872
R39074 VSS.n4502 VSS.n4416 0.00134872
R39075 VSS.n385 VSS.n383 0.00134872
R39076 VSS.n4250 VSS.n67 0.00134872
R39077 VSS.n258 VSS.n67 0.00134872
R39078 VSS.n4249 VSS.n66 0.00134872
R39079 VSS.n259 VSS.n66 0.00134872
R39080 VSS.n4248 VSS.n65 0.00134872
R39081 VSS.n260 VSS.n65 0.00134872
R39082 VSS.n4247 VSS.n64 0.00134872
R39083 VSS.n261 VSS.n64 0.00134872
R39084 VSS.n4246 VSS.n63 0.00134872
R39085 VSS.n262 VSS.n63 0.00134872
R39086 VSS.n4245 VSS.n62 0.00134872
R39087 VSS.n263 VSS.n62 0.00134872
R39088 VSS.n4244 VSS.n61 0.00134872
R39089 VSS.n264 VSS.n61 0.00134872
R39090 VSS.n4243 VSS.n60 0.00134872
R39091 VSS.n265 VSS.n60 0.00134872
R39092 VSS.n4242 VSS.n59 0.00134872
R39093 VSS.n266 VSS.n59 0.00134872
R39094 VSS.n4241 VSS.n58 0.00134872
R39095 VSS.n267 VSS.n58 0.00134872
R39096 VSS.n4240 VSS.n57 0.00134872
R39097 VSS.n268 VSS.n57 0.00134872
R39098 VSS.n4239 VSS.n56 0.00134872
R39099 VSS.n269 VSS.n56 0.00134872
R39100 VSS.n4238 VSS.n55 0.00134872
R39101 VSS.n270 VSS.n55 0.00134872
R39102 VSS.n4237 VSS.n54 0.00134872
R39103 VSS.n271 VSS.n54 0.00134872
R39104 VSS.n4236 VSS.n53 0.00134872
R39105 VSS.n272 VSS.n53 0.00134872
R39106 VSS.n4235 VSS.n52 0.00134872
R39107 VSS.n273 VSS.n52 0.00134872
R39108 VSS.n4234 VSS.n51 0.00134872
R39109 VSS.n274 VSS.n51 0.00134872
R39110 VSS.n4233 VSS.n50 0.00134872
R39111 VSS.n275 VSS.n50 0.00134872
R39112 VSS.n4232 VSS.n49 0.00134872
R39113 VSS.n276 VSS.n49 0.00134872
R39114 VSS.n4231 VSS.n48 0.00134872
R39115 VSS.n277 VSS.n48 0.00134872
R39116 VSS.n4230 VSS.n47 0.00134872
R39117 VSS.n278 VSS.n47 0.00134872
R39118 VSS.n4229 VSS.n46 0.00134872
R39119 VSS.n279 VSS.n46 0.00134872
R39120 VSS.n4228 VSS.n45 0.00134872
R39121 VSS.n280 VSS.n45 0.00134872
R39122 VSS.n4227 VSS.n44 0.00134872
R39123 VSS.n281 VSS.n44 0.00134872
R39124 VSS.n4226 VSS.n43 0.00134872
R39125 VSS.n282 VSS.n43 0.00134872
R39126 VSS.n4225 VSS.n42 0.00134872
R39127 VSS.n283 VSS.n42 0.00134872
R39128 VSS.n4224 VSS.n41 0.00134872
R39129 VSS.n284 VSS.n41 0.00134872
R39130 VSS.n4223 VSS.n40 0.00134872
R39131 VSS.n285 VSS.n40 0.00134872
R39132 VSS.n4222 VSS.n39 0.00134872
R39133 VSS.n286 VSS.n39 0.00134872
R39134 VSS.n4221 VSS.n38 0.00134872
R39135 VSS.n287 VSS.n38 0.00134872
R39136 VSS.n4220 VSS.n37 0.00134872
R39137 VSS.n288 VSS.n37 0.00134872
R39138 VSS.n4219 VSS.n36 0.00134872
R39139 VSS.n289 VSS.n36 0.00134872
R39140 VSS.n4218 VSS.n35 0.00134872
R39141 VSS.n290 VSS.n35 0.00134872
R39142 VSS.n4217 VSS.n34 0.00134872
R39143 VSS.n291 VSS.n34 0.00134872
R39144 VSS.n4216 VSS.n33 0.00134872
R39145 VSS.n292 VSS.n33 0.00134872
R39146 VSS.n4215 VSS.n32 0.00134872
R39147 VSS.n293 VSS.n32 0.00134872
R39148 VSS.n4214 VSS.n31 0.00134872
R39149 VSS.n294 VSS.n31 0.00134872
R39150 VSS.n4213 VSS.n30 0.00134872
R39151 VSS.n295 VSS.n30 0.00134872
R39152 VSS.n4212 VSS.n29 0.00134872
R39153 VSS.n296 VSS.n29 0.00134872
R39154 VSS.n4211 VSS.n28 0.00134872
R39155 VSS.n297 VSS.n28 0.00134872
R39156 VSS.n4210 VSS.n27 0.00134872
R39157 VSS.n298 VSS.n27 0.00134872
R39158 VSS.n4209 VSS.n26 0.00134872
R39159 VSS.n299 VSS.n26 0.00134872
R39160 VSS.n4208 VSS.n25 0.00134872
R39161 VSS.n300 VSS.n25 0.00134872
R39162 VSS.n4207 VSS.n24 0.00134872
R39163 VSS.n301 VSS.n24 0.00134872
R39164 VSS.n4206 VSS.n23 0.00134872
R39165 VSS.n302 VSS.n23 0.00134872
R39166 VSS.n4205 VSS.n22 0.00134872
R39167 VSS.n303 VSS.n22 0.00134872
R39168 VSS.n4204 VSS.n21 0.00134872
R39169 VSS.n304 VSS.n21 0.00134872
R39170 VSS.n4203 VSS.n20 0.00134872
R39171 VSS.n305 VSS.n20 0.00134872
R39172 VSS.n4202 VSS.n19 0.00134872
R39173 VSS.n306 VSS.n19 0.00134872
R39174 VSS.n4201 VSS.n18 0.00134872
R39175 VSS.n307 VSS.n18 0.00134872
R39176 VSS.n4200 VSS.n17 0.00134872
R39177 VSS.n308 VSS.n17 0.00134872
R39178 VSS.n4199 VSS.n16 0.00134872
R39179 VSS.n309 VSS.n16 0.00134872
R39180 VSS.n4198 VSS.n15 0.00134872
R39181 VSS.n310 VSS.n15 0.00134872
R39182 VSS.n4197 VSS.n14 0.00134872
R39183 VSS.n311 VSS.n14 0.00134872
R39184 VSS.n4196 VSS.n13 0.00134872
R39185 VSS.n312 VSS.n13 0.00134872
R39186 VSS.n4195 VSS.n12 0.00134872
R39187 VSS.n313 VSS.n12 0.00134872
R39188 VSS.n4194 VSS.n11 0.00134872
R39189 VSS.n314 VSS.n11 0.00134872
R39190 VSS.n4193 VSS.n10 0.00134872
R39191 VSS.n315 VSS.n10 0.00134872
R39192 VSS.n4192 VSS.n9 0.00134872
R39193 VSS.n316 VSS.n9 0.00134872
R39194 VSS.n4191 VSS.n8 0.00134872
R39195 VSS.n317 VSS.n8 0.00134872
R39196 VSS.n4190 VSS.n7 0.00134872
R39197 VSS.n318 VSS.n7 0.00134872
R39198 VSS.n4189 VSS.n6 0.00134872
R39199 VSS.n319 VSS.n6 0.00134872
R39200 VSS.n194 VSS.n5 0.00134872
R39201 VSS.n320 VSS.n5 0.00134872
R39202 VSS.n321 VSS.n257 0.00134872
R39203 VSS.n2857 VSS.n2479 0.00134872
R39204 VSS.n2728 VSS.n2353 0.00134872
R39205 VSS.n2856 VSS.n2478 0.00134872
R39206 VSS.n2729 VSS.n2354 0.00134872
R39207 VSS.n2855 VSS.n2477 0.00134872
R39208 VSS.n2730 VSS.n2355 0.00134872
R39209 VSS.n2854 VSS.n2476 0.00134872
R39210 VSS.n2731 VSS.n2356 0.00134872
R39211 VSS.n2853 VSS.n2475 0.00134872
R39212 VSS.n2732 VSS.n2357 0.00134872
R39213 VSS.n2852 VSS.n2474 0.00134872
R39214 VSS.n2733 VSS.n2358 0.00134872
R39215 VSS.n2851 VSS.n2473 0.00134872
R39216 VSS.n2734 VSS.n2359 0.00134872
R39217 VSS.n2850 VSS.n2472 0.00134872
R39218 VSS.n2735 VSS.n2360 0.00134872
R39219 VSS.n2849 VSS.n2471 0.00134872
R39220 VSS.n2736 VSS.n2361 0.00134872
R39221 VSS.n2848 VSS.n2470 0.00134872
R39222 VSS.n2737 VSS.n2362 0.00134872
R39223 VSS.n2847 VSS.n2469 0.00134872
R39224 VSS.n2738 VSS.n2363 0.00134872
R39225 VSS.n2846 VSS.n2468 0.00134872
R39226 VSS.n2739 VSS.n2364 0.00134872
R39227 VSS.n2845 VSS.n2467 0.00134872
R39228 VSS.n2740 VSS.n2365 0.00134872
R39229 VSS.n2844 VSS.n2466 0.00134872
R39230 VSS.n2741 VSS.n2366 0.00134872
R39231 VSS.n2843 VSS.n2465 0.00134872
R39232 VSS.n2742 VSS.n2367 0.00134872
R39233 VSS.n2842 VSS.n2464 0.00134872
R39234 VSS.n2743 VSS.n2368 0.00134872
R39235 VSS.n2841 VSS.n2463 0.00134872
R39236 VSS.n2744 VSS.n2369 0.00134872
R39237 VSS.n2840 VSS.n2462 0.00134872
R39238 VSS.n2745 VSS.n2370 0.00134872
R39239 VSS.n2839 VSS.n2461 0.00134872
R39240 VSS.n2746 VSS.n2371 0.00134872
R39241 VSS.n2838 VSS.n2460 0.00134872
R39242 VSS.n2747 VSS.n2372 0.00134872
R39243 VSS.n2837 VSS.n2459 0.00134872
R39244 VSS.n2748 VSS.n2373 0.00134872
R39245 VSS.n2836 VSS.n2458 0.00134872
R39246 VSS.n2749 VSS.n2374 0.00134872
R39247 VSS.n2835 VSS.n2457 0.00134872
R39248 VSS.n2750 VSS.n2375 0.00134872
R39249 VSS.n2834 VSS.n2456 0.00134872
R39250 VSS.n2751 VSS.n2376 0.00134872
R39251 VSS.n2833 VSS.n2455 0.00134872
R39252 VSS.n2752 VSS.n2377 0.00134872
R39253 VSS.n2832 VSS.n2454 0.00134872
R39254 VSS.n2753 VSS.n2378 0.00134872
R39255 VSS.n2831 VSS.n2453 0.00134872
R39256 VSS.n2754 VSS.n2379 0.00134872
R39257 VSS.n2830 VSS.n2452 0.00134872
R39258 VSS.n2755 VSS.n2380 0.00134872
R39259 VSS.n2829 VSS.n2451 0.00134872
R39260 VSS.n2756 VSS.n2381 0.00134872
R39261 VSS.n2828 VSS.n2450 0.00134872
R39262 VSS.n2757 VSS.n2382 0.00134872
R39263 VSS.n2827 VSS.n2449 0.00134872
R39264 VSS.n2758 VSS.n2383 0.00134872
R39265 VSS.n2826 VSS.n2448 0.00134872
R39266 VSS.n2759 VSS.n2384 0.00134872
R39267 VSS.n2825 VSS.n2447 0.00134872
R39268 VSS.n2760 VSS.n2385 0.00134872
R39269 VSS.n2824 VSS.n2446 0.00134872
R39270 VSS.n2761 VSS.n2386 0.00134872
R39271 VSS.n2823 VSS.n2445 0.00134872
R39272 VSS.n2762 VSS.n2387 0.00134872
R39273 VSS.n2822 VSS.n2444 0.00134872
R39274 VSS.n2763 VSS.n2388 0.00134872
R39275 VSS.n2821 VSS.n2443 0.00134872
R39276 VSS.n2764 VSS.n2389 0.00134872
R39277 VSS.n2820 VSS.n2442 0.00134872
R39278 VSS.n2765 VSS.n2390 0.00134872
R39279 VSS.n2819 VSS.n2441 0.00134872
R39280 VSS.n2766 VSS.n2391 0.00134872
R39281 VSS.n2818 VSS.n2440 0.00134872
R39282 VSS.n2767 VSS.n2392 0.00134872
R39283 VSS.n2817 VSS.n2439 0.00134872
R39284 VSS.n2768 VSS.n2393 0.00134872
R39285 VSS.n2816 VSS.n2438 0.00134872
R39286 VSS.n2769 VSS.n2394 0.00134872
R39287 VSS.n2815 VSS.n2437 0.00134872
R39288 VSS.n2770 VSS.n2395 0.00134872
R39289 VSS.n2814 VSS.n2436 0.00134872
R39290 VSS.n2771 VSS.n2396 0.00134872
R39291 VSS.n2813 VSS.n2435 0.00134872
R39292 VSS.n2772 VSS.n2397 0.00134872
R39293 VSS.n2812 VSS.n2434 0.00134872
R39294 VSS.n2773 VSS.n2398 0.00134872
R39295 VSS.n2811 VSS.n2433 0.00134872
R39296 VSS.n2774 VSS.n2399 0.00134872
R39297 VSS.n2810 VSS.n2432 0.00134872
R39298 VSS.n2775 VSS.n2400 0.00134872
R39299 VSS.n2809 VSS.n2431 0.00134872
R39300 VSS.n2776 VSS.n2401 0.00134872
R39301 VSS.n2808 VSS.n2430 0.00134872
R39302 VSS.n2777 VSS.n2402 0.00134872
R39303 VSS.n2807 VSS.n2429 0.00134872
R39304 VSS.n2778 VSS.n2403 0.00134872
R39305 VSS.n2806 VSS.n2428 0.00134872
R39306 VSS.n2779 VSS.n2404 0.00134872
R39307 VSS.n2805 VSS.n2427 0.00134872
R39308 VSS.n2780 VSS.n2405 0.00134872
R39309 VSS.n2804 VSS.n2426 0.00134872
R39310 VSS.n2781 VSS.n2406 0.00134872
R39311 VSS.n2803 VSS.n2425 0.00134872
R39312 VSS.n2782 VSS.n2407 0.00134872
R39313 VSS.n2802 VSS.n2424 0.00134872
R39314 VSS.n2783 VSS.n2408 0.00134872
R39315 VSS.n2801 VSS.n2423 0.00134872
R39316 VSS.n2784 VSS.n2409 0.00134872
R39317 VSS.n2800 VSS.n2422 0.00134872
R39318 VSS.n2785 VSS.n2410 0.00134872
R39319 VSS.n2799 VSS.n2421 0.00134872
R39320 VSS.n2786 VSS.n2411 0.00134872
R39321 VSS.n2798 VSS.n2420 0.00134872
R39322 VSS.n2787 VSS.n2412 0.00134872
R39323 VSS.n2797 VSS.n2419 0.00134872
R39324 VSS.n2788 VSS.n2413 0.00134872
R39325 VSS.n2796 VSS.n2418 0.00134872
R39326 VSS.n2789 VSS.n2414 0.00134872
R39327 VSS.n2795 VSS.n2417 0.00134872
R39328 VSS.n2790 VSS.n2415 0.00134872
R39329 VSS.n2794 VSS.n2416 0.00134872
R39330 VSS.n3053 VSS.n2287 0.00134872
R39331 VSS.n3052 VSS.n2351 0.00134872
R39332 VSS.n2482 VSS.n2351 0.00134872
R39333 VSS.n2484 VSS.n2350 0.00134872
R39334 VSS.n2485 VSS.n2484 0.00134872
R39335 VSS.n2489 VSS.n2349 0.00134872
R39336 VSS.n2490 VSS.n2489 0.00134872
R39337 VSS.n2492 VSS.n2348 0.00134872
R39338 VSS.n2493 VSS.n2492 0.00134872
R39339 VSS.n2497 VSS.n2347 0.00134872
R39340 VSS.n2498 VSS.n2497 0.00134872
R39341 VSS.n2500 VSS.n2346 0.00134872
R39342 VSS.n2501 VSS.n2500 0.00134872
R39343 VSS.n2505 VSS.n2345 0.00134872
R39344 VSS.n2506 VSS.n2505 0.00134872
R39345 VSS.n2508 VSS.n2344 0.00134872
R39346 VSS.n2509 VSS.n2508 0.00134872
R39347 VSS.n2513 VSS.n2343 0.00134872
R39348 VSS.n2514 VSS.n2513 0.00134872
R39349 VSS.n2516 VSS.n2342 0.00134872
R39350 VSS.n2517 VSS.n2516 0.00134872
R39351 VSS.n2521 VSS.n2341 0.00134872
R39352 VSS.n2522 VSS.n2521 0.00134872
R39353 VSS.n2524 VSS.n2340 0.00134872
R39354 VSS.n2525 VSS.n2524 0.00134872
R39355 VSS.n2529 VSS.n2339 0.00134872
R39356 VSS.n2530 VSS.n2529 0.00134872
R39357 VSS.n2532 VSS.n2338 0.00134872
R39358 VSS.n2533 VSS.n2532 0.00134872
R39359 VSS.n2537 VSS.n2337 0.00134872
R39360 VSS.n2538 VSS.n2537 0.00134872
R39361 VSS.n2540 VSS.n2336 0.00134872
R39362 VSS.n2541 VSS.n2540 0.00134872
R39363 VSS.n2545 VSS.n2335 0.00134872
R39364 VSS.n2546 VSS.n2545 0.00134872
R39365 VSS.n2548 VSS.n2334 0.00134872
R39366 VSS.n2549 VSS.n2548 0.00134872
R39367 VSS.n2553 VSS.n2333 0.00134872
R39368 VSS.n2554 VSS.n2553 0.00134872
R39369 VSS.n2556 VSS.n2332 0.00134872
R39370 VSS.n2557 VSS.n2556 0.00134872
R39371 VSS.n2561 VSS.n2331 0.00134872
R39372 VSS.n2562 VSS.n2561 0.00134872
R39373 VSS.n2564 VSS.n2330 0.00134872
R39374 VSS.n2565 VSS.n2564 0.00134872
R39375 VSS.n2569 VSS.n2329 0.00134872
R39376 VSS.n2570 VSS.n2569 0.00134872
R39377 VSS.n2572 VSS.n2328 0.00134872
R39378 VSS.n2573 VSS.n2572 0.00134872
R39379 VSS.n2577 VSS.n2327 0.00134872
R39380 VSS.n2578 VSS.n2577 0.00134872
R39381 VSS.n2580 VSS.n2326 0.00134872
R39382 VSS.n2581 VSS.n2580 0.00134872
R39383 VSS.n2585 VSS.n2325 0.00134872
R39384 VSS.n2586 VSS.n2585 0.00134872
R39385 VSS.n2588 VSS.n2324 0.00134872
R39386 VSS.n2589 VSS.n2588 0.00134872
R39387 VSS.n2593 VSS.n2323 0.00134872
R39388 VSS.n2594 VSS.n2593 0.00134872
R39389 VSS.n2596 VSS.n2322 0.00134872
R39390 VSS.n2597 VSS.n2596 0.00134872
R39391 VSS.n2601 VSS.n2321 0.00134872
R39392 VSS.n2602 VSS.n2601 0.00134872
R39393 VSS.n2604 VSS.n2320 0.00134872
R39394 VSS.n2605 VSS.n2604 0.00134872
R39395 VSS.n2609 VSS.n2319 0.00134872
R39396 VSS.n2610 VSS.n2609 0.00134872
R39397 VSS.n2612 VSS.n2318 0.00134872
R39398 VSS.n2613 VSS.n2612 0.00134872
R39399 VSS.n2617 VSS.n2317 0.00134872
R39400 VSS.n2618 VSS.n2617 0.00134872
R39401 VSS.n2620 VSS.n2316 0.00134872
R39402 VSS.n2621 VSS.n2620 0.00134872
R39403 VSS.n2625 VSS.n2315 0.00134872
R39404 VSS.n2626 VSS.n2625 0.00134872
R39405 VSS.n2628 VSS.n2314 0.00134872
R39406 VSS.n2629 VSS.n2628 0.00134872
R39407 VSS.n2633 VSS.n2313 0.00134872
R39408 VSS.n2634 VSS.n2633 0.00134872
R39409 VSS.n2636 VSS.n2312 0.00134872
R39410 VSS.n2637 VSS.n2636 0.00134872
R39411 VSS.n2640 VSS.n2311 0.00134872
R39412 VSS.n2641 VSS.n2640 0.00134872
R39413 VSS.n2643 VSS.n2310 0.00134872
R39414 VSS.n2644 VSS.n2643 0.00134872
R39415 VSS.n2648 VSS.n2309 0.00134872
R39416 VSS.n2649 VSS.n2648 0.00134872
R39417 VSS.n2651 VSS.n2308 0.00134872
R39418 VSS.n2652 VSS.n2651 0.00134872
R39419 VSS.n2656 VSS.n2307 0.00134872
R39420 VSS.n2657 VSS.n2656 0.00134872
R39421 VSS.n2659 VSS.n2306 0.00134872
R39422 VSS.n2660 VSS.n2659 0.00134872
R39423 VSS.n2664 VSS.n2305 0.00134872
R39424 VSS.n2665 VSS.n2664 0.00134872
R39425 VSS.n2667 VSS.n2304 0.00134872
R39426 VSS.n2668 VSS.n2667 0.00134872
R39427 VSS.n2672 VSS.n2303 0.00134872
R39428 VSS.n2673 VSS.n2672 0.00134872
R39429 VSS.n2675 VSS.n2302 0.00134872
R39430 VSS.n2676 VSS.n2675 0.00134872
R39431 VSS.n2680 VSS.n2301 0.00134872
R39432 VSS.n2681 VSS.n2680 0.00134872
R39433 VSS.n2683 VSS.n2300 0.00134872
R39434 VSS.n2684 VSS.n2683 0.00134872
R39435 VSS.n2688 VSS.n2299 0.00134872
R39436 VSS.n2689 VSS.n2688 0.00134872
R39437 VSS.n2691 VSS.n2298 0.00134872
R39438 VSS.n2692 VSS.n2691 0.00134872
R39439 VSS.n2696 VSS.n2297 0.00134872
R39440 VSS.n2697 VSS.n2696 0.00134872
R39441 VSS.n2699 VSS.n2296 0.00134872
R39442 VSS.n2700 VSS.n2699 0.00134872
R39443 VSS.n2704 VSS.n2295 0.00134872
R39444 VSS.n2705 VSS.n2704 0.00134872
R39445 VSS.n2707 VSS.n2294 0.00134872
R39446 VSS.n2708 VSS.n2707 0.00134872
R39447 VSS.n2712 VSS.n2293 0.00134872
R39448 VSS.n2713 VSS.n2712 0.00134872
R39449 VSS.n2715 VSS.n2292 0.00134872
R39450 VSS.n2716 VSS.n2715 0.00134872
R39451 VSS.n2720 VSS.n2291 0.00134872
R39452 VSS.n2721 VSS.n2720 0.00134872
R39453 VSS.n2723 VSS.n2290 0.00134872
R39454 VSS.n2724 VSS.n2723 0.00134872
R39455 VSS.n2791 VSS.n2289 0.00134872
R39456 VSS.n2792 VSS.n2791 0.00134872
R39457 VSS.n2858 VSS.n2288 0.00134872
R39458 VSS.n3052 VSS.n3051 0.00134872
R39459 VSS.n2483 VSS.n2350 0.00134872
R39460 VSS.n2486 VSS.n2349 0.00134872
R39461 VSS.n2491 VSS.n2348 0.00134872
R39462 VSS.n2494 VSS.n2347 0.00134872
R39463 VSS.n2499 VSS.n2346 0.00134872
R39464 VSS.n2502 VSS.n2345 0.00134872
R39465 VSS.n2507 VSS.n2344 0.00134872
R39466 VSS.n2510 VSS.n2343 0.00134872
R39467 VSS.n2515 VSS.n2342 0.00134872
R39468 VSS.n2518 VSS.n2341 0.00134872
R39469 VSS.n2523 VSS.n2340 0.00134872
R39470 VSS.n2526 VSS.n2339 0.00134872
R39471 VSS.n2531 VSS.n2338 0.00134872
R39472 VSS.n2534 VSS.n2337 0.00134872
R39473 VSS.n2539 VSS.n2336 0.00134872
R39474 VSS.n2542 VSS.n2335 0.00134872
R39475 VSS.n2547 VSS.n2334 0.00134872
R39476 VSS.n2550 VSS.n2333 0.00134872
R39477 VSS.n2555 VSS.n2332 0.00134872
R39478 VSS.n2558 VSS.n2331 0.00134872
R39479 VSS.n2563 VSS.n2330 0.00134872
R39480 VSS.n2566 VSS.n2329 0.00134872
R39481 VSS.n2571 VSS.n2328 0.00134872
R39482 VSS.n2574 VSS.n2327 0.00134872
R39483 VSS.n2579 VSS.n2326 0.00134872
R39484 VSS.n2582 VSS.n2325 0.00134872
R39485 VSS.n2587 VSS.n2324 0.00134872
R39486 VSS.n2590 VSS.n2323 0.00134872
R39487 VSS.n2595 VSS.n2322 0.00134872
R39488 VSS.n2598 VSS.n2321 0.00134872
R39489 VSS.n2603 VSS.n2320 0.00134872
R39490 VSS.n2606 VSS.n2319 0.00134872
R39491 VSS.n2611 VSS.n2318 0.00134872
R39492 VSS.n2614 VSS.n2317 0.00134872
R39493 VSS.n2619 VSS.n2316 0.00134872
R39494 VSS.n2622 VSS.n2315 0.00134872
R39495 VSS.n2627 VSS.n2314 0.00134872
R39496 VSS.n2630 VSS.n2313 0.00134872
R39497 VSS.n2635 VSS.n2312 0.00134872
R39498 VSS.n2638 VSS.n2311 0.00134872
R39499 VSS.n2642 VSS.n2310 0.00134872
R39500 VSS.n2645 VSS.n2309 0.00134872
R39501 VSS.n2650 VSS.n2308 0.00134872
R39502 VSS.n2653 VSS.n2307 0.00134872
R39503 VSS.n2658 VSS.n2306 0.00134872
R39504 VSS.n2661 VSS.n2305 0.00134872
R39505 VSS.n2666 VSS.n2304 0.00134872
R39506 VSS.n2669 VSS.n2303 0.00134872
R39507 VSS.n2674 VSS.n2302 0.00134872
R39508 VSS.n2677 VSS.n2301 0.00134872
R39509 VSS.n2682 VSS.n2300 0.00134872
R39510 VSS.n2685 VSS.n2299 0.00134872
R39511 VSS.n2690 VSS.n2298 0.00134872
R39512 VSS.n2693 VSS.n2297 0.00134872
R39513 VSS.n2698 VSS.n2296 0.00134872
R39514 VSS.n2701 VSS.n2295 0.00134872
R39515 VSS.n2706 VSS.n2294 0.00134872
R39516 VSS.n2709 VSS.n2293 0.00134872
R39517 VSS.n2714 VSS.n2292 0.00134872
R39518 VSS.n2717 VSS.n2291 0.00134872
R39519 VSS.n2722 VSS.n2290 0.00134872
R39520 VSS.n2725 VSS.n2289 0.00134872
R39521 VSS.n2793 VSS.n2288 0.00134872
R39522 VSS.n2483 VSS.n2482 0.00134872
R39523 VSS.n2486 VSS.n2485 0.00134872
R39524 VSS.n2491 VSS.n2490 0.00134872
R39525 VSS.n2494 VSS.n2493 0.00134872
R39526 VSS.n2499 VSS.n2498 0.00134872
R39527 VSS.n2502 VSS.n2501 0.00134872
R39528 VSS.n2507 VSS.n2506 0.00134872
R39529 VSS.n2510 VSS.n2509 0.00134872
R39530 VSS.n2515 VSS.n2514 0.00134872
R39531 VSS.n2518 VSS.n2517 0.00134872
R39532 VSS.n2523 VSS.n2522 0.00134872
R39533 VSS.n2526 VSS.n2525 0.00134872
R39534 VSS.n2531 VSS.n2530 0.00134872
R39535 VSS.n2534 VSS.n2533 0.00134872
R39536 VSS.n2539 VSS.n2538 0.00134872
R39537 VSS.n2542 VSS.n2541 0.00134872
R39538 VSS.n2547 VSS.n2546 0.00134872
R39539 VSS.n2550 VSS.n2549 0.00134872
R39540 VSS.n2555 VSS.n2554 0.00134872
R39541 VSS.n2558 VSS.n2557 0.00134872
R39542 VSS.n2563 VSS.n2562 0.00134872
R39543 VSS.n2566 VSS.n2565 0.00134872
R39544 VSS.n2571 VSS.n2570 0.00134872
R39545 VSS.n2574 VSS.n2573 0.00134872
R39546 VSS.n2579 VSS.n2578 0.00134872
R39547 VSS.n2582 VSS.n2581 0.00134872
R39548 VSS.n2587 VSS.n2586 0.00134872
R39549 VSS.n2590 VSS.n2589 0.00134872
R39550 VSS.n2595 VSS.n2594 0.00134872
R39551 VSS.n2598 VSS.n2597 0.00134872
R39552 VSS.n2603 VSS.n2602 0.00134872
R39553 VSS.n2606 VSS.n2605 0.00134872
R39554 VSS.n2611 VSS.n2610 0.00134872
R39555 VSS.n2614 VSS.n2613 0.00134872
R39556 VSS.n2619 VSS.n2618 0.00134872
R39557 VSS.n2622 VSS.n2621 0.00134872
R39558 VSS.n2627 VSS.n2626 0.00134872
R39559 VSS.n2630 VSS.n2629 0.00134872
R39560 VSS.n2635 VSS.n2634 0.00134872
R39561 VSS.n2638 VSS.n2637 0.00134872
R39562 VSS.n2642 VSS.n2641 0.00134872
R39563 VSS.n2645 VSS.n2644 0.00134872
R39564 VSS.n2650 VSS.n2649 0.00134872
R39565 VSS.n2653 VSS.n2652 0.00134872
R39566 VSS.n2658 VSS.n2657 0.00134872
R39567 VSS.n2661 VSS.n2660 0.00134872
R39568 VSS.n2666 VSS.n2665 0.00134872
R39569 VSS.n2669 VSS.n2668 0.00134872
R39570 VSS.n2674 VSS.n2673 0.00134872
R39571 VSS.n2677 VSS.n2676 0.00134872
R39572 VSS.n2682 VSS.n2681 0.00134872
R39573 VSS.n2685 VSS.n2684 0.00134872
R39574 VSS.n2690 VSS.n2689 0.00134872
R39575 VSS.n2693 VSS.n2692 0.00134872
R39576 VSS.n2698 VSS.n2697 0.00134872
R39577 VSS.n2701 VSS.n2700 0.00134872
R39578 VSS.n2706 VSS.n2705 0.00134872
R39579 VSS.n2709 VSS.n2708 0.00134872
R39580 VSS.n2714 VSS.n2713 0.00134872
R39581 VSS.n2717 VSS.n2716 0.00134872
R39582 VSS.n2722 VSS.n2721 0.00134872
R39583 VSS.n2725 VSS.n2724 0.00134872
R39584 VSS.n2793 VSS.n2792 0.00134872
R39585 VSS.n2416 VSS.n2287 0.00134872
R39586 VSS.n2794 VSS.n2415 0.00134872
R39587 VSS.n2790 VSS.n2417 0.00134872
R39588 VSS.n2795 VSS.n2414 0.00134872
R39589 VSS.n2789 VSS.n2418 0.00134872
R39590 VSS.n2796 VSS.n2413 0.00134872
R39591 VSS.n2788 VSS.n2419 0.00134872
R39592 VSS.n2797 VSS.n2412 0.00134872
R39593 VSS.n2787 VSS.n2420 0.00134872
R39594 VSS.n2798 VSS.n2411 0.00134872
R39595 VSS.n2786 VSS.n2421 0.00134872
R39596 VSS.n2799 VSS.n2410 0.00134872
R39597 VSS.n2785 VSS.n2422 0.00134872
R39598 VSS.n2800 VSS.n2409 0.00134872
R39599 VSS.n2784 VSS.n2423 0.00134872
R39600 VSS.n2801 VSS.n2408 0.00134872
R39601 VSS.n2783 VSS.n2424 0.00134872
R39602 VSS.n2802 VSS.n2407 0.00134872
R39603 VSS.n2782 VSS.n2425 0.00134872
R39604 VSS.n2803 VSS.n2406 0.00134872
R39605 VSS.n2781 VSS.n2426 0.00134872
R39606 VSS.n2804 VSS.n2405 0.00134872
R39607 VSS.n2780 VSS.n2427 0.00134872
R39608 VSS.n2805 VSS.n2404 0.00134872
R39609 VSS.n2779 VSS.n2428 0.00134872
R39610 VSS.n2806 VSS.n2403 0.00134872
R39611 VSS.n2778 VSS.n2429 0.00134872
R39612 VSS.n2807 VSS.n2402 0.00134872
R39613 VSS.n2777 VSS.n2430 0.00134872
R39614 VSS.n2808 VSS.n2401 0.00134872
R39615 VSS.n2776 VSS.n2431 0.00134872
R39616 VSS.n2809 VSS.n2400 0.00134872
R39617 VSS.n2775 VSS.n2432 0.00134872
R39618 VSS.n2810 VSS.n2399 0.00134872
R39619 VSS.n2774 VSS.n2433 0.00134872
R39620 VSS.n2811 VSS.n2398 0.00134872
R39621 VSS.n2773 VSS.n2434 0.00134872
R39622 VSS.n2812 VSS.n2397 0.00134872
R39623 VSS.n2772 VSS.n2435 0.00134872
R39624 VSS.n2813 VSS.n2396 0.00134872
R39625 VSS.n2771 VSS.n2436 0.00134872
R39626 VSS.n2814 VSS.n2395 0.00134872
R39627 VSS.n2770 VSS.n2437 0.00134872
R39628 VSS.n2815 VSS.n2394 0.00134872
R39629 VSS.n2769 VSS.n2438 0.00134872
R39630 VSS.n2816 VSS.n2393 0.00134872
R39631 VSS.n2768 VSS.n2439 0.00134872
R39632 VSS.n2817 VSS.n2392 0.00134872
R39633 VSS.n2767 VSS.n2440 0.00134872
R39634 VSS.n2818 VSS.n2391 0.00134872
R39635 VSS.n2766 VSS.n2441 0.00134872
R39636 VSS.n2819 VSS.n2390 0.00134872
R39637 VSS.n2765 VSS.n2442 0.00134872
R39638 VSS.n2820 VSS.n2389 0.00134872
R39639 VSS.n2764 VSS.n2443 0.00134872
R39640 VSS.n2821 VSS.n2388 0.00134872
R39641 VSS.n2763 VSS.n2444 0.00134872
R39642 VSS.n2822 VSS.n2387 0.00134872
R39643 VSS.n2762 VSS.n2445 0.00134872
R39644 VSS.n2823 VSS.n2386 0.00134872
R39645 VSS.n2761 VSS.n2446 0.00134872
R39646 VSS.n2824 VSS.n2385 0.00134872
R39647 VSS.n2760 VSS.n2447 0.00134872
R39648 VSS.n2825 VSS.n2384 0.00134872
R39649 VSS.n2759 VSS.n2448 0.00134872
R39650 VSS.n2826 VSS.n2383 0.00134872
R39651 VSS.n2758 VSS.n2449 0.00134872
R39652 VSS.n2827 VSS.n2382 0.00134872
R39653 VSS.n2757 VSS.n2450 0.00134872
R39654 VSS.n2828 VSS.n2381 0.00134872
R39655 VSS.n2756 VSS.n2451 0.00134872
R39656 VSS.n2829 VSS.n2380 0.00134872
R39657 VSS.n2755 VSS.n2452 0.00134872
R39658 VSS.n2830 VSS.n2379 0.00134872
R39659 VSS.n2754 VSS.n2453 0.00134872
R39660 VSS.n2831 VSS.n2378 0.00134872
R39661 VSS.n2753 VSS.n2454 0.00134872
R39662 VSS.n2832 VSS.n2377 0.00134872
R39663 VSS.n2752 VSS.n2455 0.00134872
R39664 VSS.n2833 VSS.n2376 0.00134872
R39665 VSS.n2751 VSS.n2456 0.00134872
R39666 VSS.n2834 VSS.n2375 0.00134872
R39667 VSS.n2750 VSS.n2457 0.00134872
R39668 VSS.n2835 VSS.n2374 0.00134872
R39669 VSS.n2749 VSS.n2458 0.00134872
R39670 VSS.n2836 VSS.n2373 0.00134872
R39671 VSS.n2748 VSS.n2459 0.00134872
R39672 VSS.n2837 VSS.n2372 0.00134872
R39673 VSS.n2747 VSS.n2460 0.00134872
R39674 VSS.n2838 VSS.n2371 0.00134872
R39675 VSS.n2746 VSS.n2461 0.00134872
R39676 VSS.n2839 VSS.n2370 0.00134872
R39677 VSS.n2745 VSS.n2462 0.00134872
R39678 VSS.n2840 VSS.n2369 0.00134872
R39679 VSS.n2744 VSS.n2463 0.00134872
R39680 VSS.n2841 VSS.n2368 0.00134872
R39681 VSS.n2743 VSS.n2464 0.00134872
R39682 VSS.n2842 VSS.n2367 0.00134872
R39683 VSS.n2742 VSS.n2465 0.00134872
R39684 VSS.n2843 VSS.n2366 0.00134872
R39685 VSS.n2741 VSS.n2466 0.00134872
R39686 VSS.n2844 VSS.n2365 0.00134872
R39687 VSS.n2740 VSS.n2467 0.00134872
R39688 VSS.n2845 VSS.n2364 0.00134872
R39689 VSS.n2739 VSS.n2468 0.00134872
R39690 VSS.n2846 VSS.n2363 0.00134872
R39691 VSS.n2738 VSS.n2469 0.00134872
R39692 VSS.n2847 VSS.n2362 0.00134872
R39693 VSS.n2737 VSS.n2470 0.00134872
R39694 VSS.n2848 VSS.n2361 0.00134872
R39695 VSS.n2736 VSS.n2471 0.00134872
R39696 VSS.n2849 VSS.n2360 0.00134872
R39697 VSS.n2735 VSS.n2472 0.00134872
R39698 VSS.n2850 VSS.n2359 0.00134872
R39699 VSS.n2734 VSS.n2473 0.00134872
R39700 VSS.n2851 VSS.n2358 0.00134872
R39701 VSS.n2733 VSS.n2474 0.00134872
R39702 VSS.n2852 VSS.n2357 0.00134872
R39703 VSS.n2732 VSS.n2475 0.00134872
R39704 VSS.n2853 VSS.n2356 0.00134872
R39705 VSS.n2731 VSS.n2476 0.00134872
R39706 VSS.n2854 VSS.n2355 0.00134872
R39707 VSS.n2730 VSS.n2477 0.00134872
R39708 VSS.n2855 VSS.n2354 0.00134872
R39709 VSS.n2729 VSS.n2478 0.00134872
R39710 VSS.n2856 VSS.n2353 0.00134872
R39711 VSS.n2728 VSS.n2479 0.00134872
R39712 VSS.n2857 VSS.n2352 0.00134872
R39713 VSS.n4413 VSS.n4252 0.00134303
R39714 VSS.n4500 VSS.n384 0.00134303
R39715 VSS.n2861 VSS.n2860 0.00134303
R39716 VSS.n4411 VSS.n4252 0.0011975
R39717 VSS.n4411 VSS.n4410 0.0011975
R39718 VSS.n4410 VSS.n4409 0.0011975
R39719 VSS.n4409 VSS.n4408 0.0011975
R39720 VSS.n4408 VSS.n4407 0.0011975
R39721 VSS.n4407 VSS.n4406 0.0011975
R39722 VSS.n4406 VSS.n4405 0.0011975
R39723 VSS.n4405 VSS.n4404 0.0011975
R39724 VSS.n4404 VSS.n4403 0.0011975
R39725 VSS.n4403 VSS.n4402 0.0011975
R39726 VSS.n4402 VSS.n4401 0.0011975
R39727 VSS.n4401 VSS.n4400 0.0011975
R39728 VSS.n4400 VSS.n4399 0.0011975
R39729 VSS.n4399 VSS.n4398 0.0011975
R39730 VSS.n4398 VSS.n4397 0.0011975
R39731 VSS.n4397 VSS.n4396 0.0011975
R39732 VSS.n4396 VSS.n4395 0.0011975
R39733 VSS.n4395 VSS.n4394 0.0011975
R39734 VSS.n4394 VSS.n4393 0.0011975
R39735 VSS.n4393 VSS.n4392 0.0011975
R39736 VSS.n4392 VSS.n4391 0.0011975
R39737 VSS.n4391 VSS.n4390 0.0011975
R39738 VSS.n4390 VSS.n4389 0.0011975
R39739 VSS.n4389 VSS.n4388 0.0011975
R39740 VSS.n4388 VSS.n4387 0.0011975
R39741 VSS.n4387 VSS.n4386 0.0011975
R39742 VSS.n4386 VSS.n4385 0.0011975
R39743 VSS.n4385 VSS.n4384 0.0011975
R39744 VSS.n4384 VSS.n4383 0.0011975
R39745 VSS.n4383 VSS.n4382 0.0011975
R39746 VSS.n4382 VSS.n4381 0.0011975
R39747 VSS.n4381 VSS.n4380 0.0011975
R39748 VSS.n4380 VSS.n4379 0.0011975
R39749 VSS.n4379 VSS.n4378 0.0011975
R39750 VSS.n4378 VSS.n4377 0.0011975
R39751 VSS.n4377 VSS.n4376 0.0011975
R39752 VSS.n4376 VSS.n4375 0.0011975
R39753 VSS.n4375 VSS.n4374 0.0011975
R39754 VSS.n4374 VSS.n4373 0.0011975
R39755 VSS.n4373 VSS.n4372 0.0011975
R39756 VSS.n4372 VSS.n4371 0.0011975
R39757 VSS.n4371 VSS.n4370 0.0011975
R39758 VSS.n4370 VSS.n4369 0.0011975
R39759 VSS.n4369 VSS.n4368 0.0011975
R39760 VSS.n4368 VSS.n4367 0.0011975
R39761 VSS.n4367 VSS.n4366 0.0011975
R39762 VSS.n4366 VSS.n4365 0.0011975
R39763 VSS.n4365 VSS.n4364 0.0011975
R39764 VSS.n4364 VSS.n4363 0.0011975
R39765 VSS.n4363 VSS.n4362 0.0011975
R39766 VSS.n4362 VSS.n4361 0.0011975
R39767 VSS.n4361 VSS.n4360 0.0011975
R39768 VSS.n4360 VSS.n4359 0.0011975
R39769 VSS.n4359 VSS.n4358 0.0011975
R39770 VSS.n4358 VSS.n4357 0.0011975
R39771 VSS.n4357 VSS.n4356 0.0011975
R39772 VSS.n4356 VSS.n4355 0.0011975
R39773 VSS.n4355 VSS.n4354 0.0011975
R39774 VSS.n4354 VSS.n4353 0.0011975
R39775 VSS.n4353 VSS.n4352 0.0011975
R39776 VSS.n4352 VSS.n4351 0.0011975
R39777 VSS.n4351 VSS.n4350 0.0011975
R39778 VSS.n4350 VSS.n4349 0.0011975
R39779 VSS.n4349 VSS.n4348 0.0011975
R39780 VSS.n4348 VSS.n4347 0.0011975
R39781 VSS.n4347 VSS.n4346 0.0011975
R39782 VSS.n4346 VSS.n4345 0.0011975
R39783 VSS.n4345 VSS.n4344 0.0011975
R39784 VSS.n4344 VSS.n4343 0.0011975
R39785 VSS.n4343 VSS.n4342 0.0011975
R39786 VSS.n4342 VSS.n4341 0.0011975
R39787 VSS.n4341 VSS.n4340 0.0011975
R39788 VSS.n4340 VSS.n4339 0.0011975
R39789 VSS.n4339 VSS.n4338 0.0011975
R39790 VSS.n4338 VSS.n4337 0.0011975
R39791 VSS.n4337 VSS.n4336 0.0011975
R39792 VSS.n4336 VSS.n4335 0.0011975
R39793 VSS.n4335 VSS.n4334 0.0011975
R39794 VSS.n4334 VSS.n4333 0.0011975
R39795 VSS.n4333 VSS.n4332 0.0011975
R39796 VSS.n4332 VSS.n2 0.0011975
R39797 VSS.n4507 VSS.n2 0.0011975
R39798 VSS.n4507 VSS.n3 0.0011975
R39799 VSS.n4437 VSS.n3 0.0011975
R39800 VSS.n4440 VSS.n4437 0.0011975
R39801 VSS.n4441 VSS.n4440 0.0011975
R39802 VSS.n4442 VSS.n4441 0.0011975
R39803 VSS.n4442 VSS.n4435 0.0011975
R39804 VSS.n4446 VSS.n4435 0.0011975
R39805 VSS.n4447 VSS.n4446 0.0011975
R39806 VSS.n4448 VSS.n4447 0.0011975
R39807 VSS.n4448 VSS.n4433 0.0011975
R39808 VSS.n4452 VSS.n4433 0.0011975
R39809 VSS.n4453 VSS.n4452 0.0011975
R39810 VSS.n4454 VSS.n4453 0.0011975
R39811 VSS.n4454 VSS.n4431 0.0011975
R39812 VSS.n4458 VSS.n4431 0.0011975
R39813 VSS.n4459 VSS.n4458 0.0011975
R39814 VSS.n4460 VSS.n4459 0.0011975
R39815 VSS.n4460 VSS.n4429 0.0011975
R39816 VSS.n4464 VSS.n4429 0.0011975
R39817 VSS.n4465 VSS.n4464 0.0011975
R39818 VSS.n4466 VSS.n4465 0.0011975
R39819 VSS.n4466 VSS.n4427 0.0011975
R39820 VSS.n4470 VSS.n4427 0.0011975
R39821 VSS.n4471 VSS.n4470 0.0011975
R39822 VSS.n4472 VSS.n4471 0.0011975
R39823 VSS.n4472 VSS.n4425 0.0011975
R39824 VSS.n4476 VSS.n4425 0.0011975
R39825 VSS.n4477 VSS.n4476 0.0011975
R39826 VSS.n4478 VSS.n4477 0.0011975
R39827 VSS.n4478 VSS.n4423 0.0011975
R39828 VSS.n4482 VSS.n4423 0.0011975
R39829 VSS.n4483 VSS.n4482 0.0011975
R39830 VSS.n4484 VSS.n4483 0.0011975
R39831 VSS.n4484 VSS.n4421 0.0011975
R39832 VSS.n4488 VSS.n4421 0.0011975
R39833 VSS.n4489 VSS.n4488 0.0011975
R39834 VSS.n4490 VSS.n4489 0.0011975
R39835 VSS.n4490 VSS.n4419 0.0011975
R39836 VSS.n4494 VSS.n4419 0.0011975
R39837 VSS.n4495 VSS.n4494 0.0011975
R39838 VSS.n4496 VSS.n4495 0.0011975
R39839 VSS.n4496 VSS.n4417 0.0011975
R39840 VSS.n4501 VSS.n4417 0.0011975
R39841 VSS.n4501 VSS.n4500 0.0011975
R39842 VSS.n4504 VSS.n321 0.0011975
R39843 VSS.n2859 VSS.n2858 0.0011975
R39844 VSS.n3048 VSS.n2480 0.0011975
R39845 VSS.n3048 VSS.n3047 0.0011975
R39846 VSS.n3047 VSS.n3046 0.0011975
R39847 VSS.n3046 VSS.n2487 0.0011975
R39848 VSS.n3042 VSS.n2487 0.0011975
R39849 VSS.n3042 VSS.n3041 0.0011975
R39850 VSS.n3041 VSS.n3040 0.0011975
R39851 VSS.n3040 VSS.n2495 0.0011975
R39852 VSS.n3036 VSS.n2495 0.0011975
R39853 VSS.n3036 VSS.n3035 0.0011975
R39854 VSS.n3035 VSS.n3034 0.0011975
R39855 VSS.n3034 VSS.n2503 0.0011975
R39856 VSS.n3030 VSS.n2503 0.0011975
R39857 VSS.n3030 VSS.n3029 0.0011975
R39858 VSS.n3029 VSS.n3028 0.0011975
R39859 VSS.n3028 VSS.n2511 0.0011975
R39860 VSS.n3024 VSS.n2511 0.0011975
R39861 VSS.n3024 VSS.n3023 0.0011975
R39862 VSS.n3023 VSS.n3022 0.0011975
R39863 VSS.n3022 VSS.n2519 0.0011975
R39864 VSS.n3018 VSS.n2519 0.0011975
R39865 VSS.n3018 VSS.n3017 0.0011975
R39866 VSS.n3017 VSS.n3016 0.0011975
R39867 VSS.n3016 VSS.n2527 0.0011975
R39868 VSS.n3012 VSS.n2527 0.0011975
R39869 VSS.n3012 VSS.n3011 0.0011975
R39870 VSS.n3011 VSS.n3010 0.0011975
R39871 VSS.n3010 VSS.n2535 0.0011975
R39872 VSS.n3006 VSS.n2535 0.0011975
R39873 VSS.n3006 VSS.n3005 0.0011975
R39874 VSS.n3005 VSS.n3004 0.0011975
R39875 VSS.n3004 VSS.n2543 0.0011975
R39876 VSS.n3000 VSS.n2543 0.0011975
R39877 VSS.n3000 VSS.n2999 0.0011975
R39878 VSS.n2999 VSS.n2998 0.0011975
R39879 VSS.n2998 VSS.n2551 0.0011975
R39880 VSS.n2994 VSS.n2551 0.0011975
R39881 VSS.n2994 VSS.n2993 0.0011975
R39882 VSS.n2993 VSS.n2992 0.0011975
R39883 VSS.n2992 VSS.n2559 0.0011975
R39884 VSS.n2988 VSS.n2559 0.0011975
R39885 VSS.n2988 VSS.n2987 0.0011975
R39886 VSS.n2987 VSS.n2986 0.0011975
R39887 VSS.n2986 VSS.n2567 0.0011975
R39888 VSS.n2982 VSS.n2567 0.0011975
R39889 VSS.n2982 VSS.n2981 0.0011975
R39890 VSS.n2981 VSS.n2980 0.0011975
R39891 VSS.n2980 VSS.n2575 0.0011975
R39892 VSS.n2976 VSS.n2575 0.0011975
R39893 VSS.n2976 VSS.n2975 0.0011975
R39894 VSS.n2975 VSS.n2974 0.0011975
R39895 VSS.n2974 VSS.n2583 0.0011975
R39896 VSS.n2970 VSS.n2583 0.0011975
R39897 VSS.n2970 VSS.n2969 0.0011975
R39898 VSS.n2969 VSS.n2968 0.0011975
R39899 VSS.n2968 VSS.n2591 0.0011975
R39900 VSS.n2964 VSS.n2591 0.0011975
R39901 VSS.n2964 VSS.n2963 0.0011975
R39902 VSS.n2963 VSS.n2962 0.0011975
R39903 VSS.n2962 VSS.n2599 0.0011975
R39904 VSS.n2958 VSS.n2599 0.0011975
R39905 VSS.n2958 VSS.n2957 0.0011975
R39906 VSS.n2957 VSS.n2956 0.0011975
R39907 VSS.n2956 VSS.n2607 0.0011975
R39908 VSS.n2952 VSS.n2607 0.0011975
R39909 VSS.n2952 VSS.n2951 0.0011975
R39910 VSS.n2951 VSS.n2950 0.0011975
R39911 VSS.n2950 VSS.n2615 0.0011975
R39912 VSS.n2946 VSS.n2615 0.0011975
R39913 VSS.n2946 VSS.n2945 0.0011975
R39914 VSS.n2945 VSS.n2944 0.0011975
R39915 VSS.n2944 VSS.n2623 0.0011975
R39916 VSS.n2940 VSS.n2623 0.0011975
R39917 VSS.n2940 VSS.n2939 0.0011975
R39918 VSS.n2939 VSS.n2938 0.0011975
R39919 VSS.n2938 VSS.n2631 0.0011975
R39920 VSS.n2934 VSS.n2631 0.0011975
R39921 VSS.n2934 VSS.n2933 0.0011975
R39922 VSS.n2933 VSS.n2932 0.0011975
R39923 VSS.n2932 VSS.n2639 0.0011975
R39924 VSS.n2928 VSS.n2639 0.0011975
R39925 VSS.n2928 VSS.n2927 0.0011975
R39926 VSS.n2927 VSS.n2646 0.0011975
R39927 VSS.n2923 VSS.n2646 0.0011975
R39928 VSS.n2923 VSS.n2922 0.0011975
R39929 VSS.n2922 VSS.n2921 0.0011975
R39930 VSS.n2921 VSS.n2654 0.0011975
R39931 VSS.n2917 VSS.n2654 0.0011975
R39932 VSS.n2917 VSS.n2916 0.0011975
R39933 VSS.n2916 VSS.n2915 0.0011975
R39934 VSS.n2915 VSS.n2662 0.0011975
R39935 VSS.n2911 VSS.n2662 0.0011975
R39936 VSS.n2911 VSS.n2910 0.0011975
R39937 VSS.n2910 VSS.n2909 0.0011975
R39938 VSS.n2909 VSS.n2670 0.0011975
R39939 VSS.n2905 VSS.n2670 0.0011975
R39940 VSS.n2905 VSS.n2904 0.0011975
R39941 VSS.n2904 VSS.n2903 0.0011975
R39942 VSS.n2903 VSS.n2678 0.0011975
R39943 VSS.n2899 VSS.n2678 0.0011975
R39944 VSS.n2899 VSS.n2898 0.0011975
R39945 VSS.n2898 VSS.n2897 0.0011975
R39946 VSS.n2897 VSS.n2686 0.0011975
R39947 VSS.n2893 VSS.n2686 0.0011975
R39948 VSS.n2893 VSS.n2892 0.0011975
R39949 VSS.n2892 VSS.n2891 0.0011975
R39950 VSS.n2891 VSS.n2694 0.0011975
R39951 VSS.n2887 VSS.n2694 0.0011975
R39952 VSS.n2887 VSS.n2886 0.0011975
R39953 VSS.n2886 VSS.n2885 0.0011975
R39954 VSS.n2885 VSS.n2702 0.0011975
R39955 VSS.n2881 VSS.n2702 0.0011975
R39956 VSS.n2881 VSS.n2880 0.0011975
R39957 VSS.n2880 VSS.n2879 0.0011975
R39958 VSS.n2879 VSS.n2710 0.0011975
R39959 VSS.n2875 VSS.n2710 0.0011975
R39960 VSS.n2875 VSS.n2874 0.0011975
R39961 VSS.n2874 VSS.n2873 0.0011975
R39962 VSS.n2873 VSS.n2718 0.0011975
R39963 VSS.n2869 VSS.n2718 0.0011975
R39964 VSS.n2869 VSS.n2868 0.0011975
R39965 VSS.n2868 VSS.n2867 0.0011975
R39966 VSS.n2867 VSS.n2726 0.0011975
R39967 VSS.n2863 VSS.n2726 0.0011975
R39968 VSS.n2863 VSS.n2862 0.0011975
R39969 VSS.n2862 VSS.n2861 0.0011975
R39970 VSS.n4412 VSS.n4253 0.000965
R39971 VSS.n4254 VSS.n4253 0.000965
R39972 VSS.n4255 VSS.n4254 0.000965
R39973 VSS.n4256 VSS.n4255 0.000965
R39974 VSS.n4257 VSS.n4256 0.000965
R39975 VSS.n4258 VSS.n4257 0.000965
R39976 VSS.n4259 VSS.n4258 0.000965
R39977 VSS.n4260 VSS.n4259 0.000965
R39978 VSS.n4261 VSS.n4260 0.000965
R39979 VSS.n4262 VSS.n4261 0.000965
R39980 VSS.n4263 VSS.n4262 0.000965
R39981 VSS.n4264 VSS.n4263 0.000965
R39982 VSS.n4265 VSS.n4264 0.000965
R39983 VSS.n4266 VSS.n4265 0.000965
R39984 VSS.n4267 VSS.n4266 0.000965
R39985 VSS.n4268 VSS.n4267 0.000965
R39986 VSS.n4269 VSS.n4268 0.000965
R39987 VSS.n4270 VSS.n4269 0.000965
R39988 VSS.n4271 VSS.n4270 0.000965
R39989 VSS.n4272 VSS.n4271 0.000965
R39990 VSS.n4273 VSS.n4272 0.000965
R39991 VSS.n4274 VSS.n4273 0.000965
R39992 VSS.n4275 VSS.n4274 0.000965
R39993 VSS.n4276 VSS.n4275 0.000965
R39994 VSS.n4277 VSS.n4276 0.000965
R39995 VSS.n4278 VSS.n4277 0.000965
R39996 VSS.n4279 VSS.n4278 0.000965
R39997 VSS.n4280 VSS.n4279 0.000965
R39998 VSS.n4281 VSS.n4280 0.000965
R39999 VSS.n4282 VSS.n4281 0.000965
R40000 VSS.n4283 VSS.n4282 0.000965
R40001 VSS.n4284 VSS.n4283 0.000965
R40002 VSS.n4285 VSS.n4284 0.000965
R40003 VSS.n4286 VSS.n4285 0.000965
R40004 VSS.n4287 VSS.n4286 0.000965
R40005 VSS.n4288 VSS.n4287 0.000965
R40006 VSS.n4289 VSS.n4288 0.000965
R40007 VSS.n4290 VSS.n4289 0.000965
R40008 VSS.n4291 VSS.n4290 0.000965
R40009 VSS.n4292 VSS.n4291 0.000965
R40010 VSS.n4293 VSS.n4292 0.000965
R40011 VSS.n4294 VSS.n4293 0.000965
R40012 VSS.n4295 VSS.n4294 0.000965
R40013 VSS.n4296 VSS.n4295 0.000965
R40014 VSS.n4297 VSS.n4296 0.000965
R40015 VSS.n4298 VSS.n4297 0.000965
R40016 VSS.n4299 VSS.n4298 0.000965
R40017 VSS.n4300 VSS.n4299 0.000965
R40018 VSS.n4301 VSS.n4300 0.000965
R40019 VSS.n4302 VSS.n4301 0.000965
R40020 VSS.n4303 VSS.n4302 0.000965
R40021 VSS.n4304 VSS.n4303 0.000965
R40022 VSS.n4305 VSS.n4304 0.000965
R40023 VSS.n4306 VSS.n4305 0.000965
R40024 VSS.n4307 VSS.n4306 0.000965
R40025 VSS.n4308 VSS.n4307 0.000965
R40026 VSS.n4309 VSS.n4308 0.000965
R40027 VSS.n4310 VSS.n4309 0.000965
R40028 VSS.n4311 VSS.n4310 0.000965
R40029 VSS.n4312 VSS.n4311 0.000965
R40030 VSS.n4313 VSS.n4312 0.000965
R40031 VSS.n4314 VSS.n4313 0.000965
R40032 VSS.n4315 VSS.n4314 0.000965
R40033 VSS.n4316 VSS.n4315 0.000965
R40034 VSS.n4317 VSS.n4316 0.000965
R40035 VSS.n4318 VSS.n4317 0.000965
R40036 VSS.n4319 VSS.n4318 0.000965
R40037 VSS.n4320 VSS.n4319 0.000965
R40038 VSS.n4321 VSS.n4320 0.000965
R40039 VSS.n4322 VSS.n4321 0.000965
R40040 VSS.n4323 VSS.n4322 0.000965
R40041 VSS.n4324 VSS.n4323 0.000965
R40042 VSS.n4325 VSS.n4324 0.000965
R40043 VSS.n4326 VSS.n4325 0.000965
R40044 VSS.n4327 VSS.n4326 0.000965
R40045 VSS.n4328 VSS.n4327 0.000965
R40046 VSS.n4329 VSS.n4328 0.000965
R40047 VSS.n4330 VSS.n4329 0.000965
R40048 VSS.n4331 VSS.n4330 0.000965
R40049 VSS.n4331 VSS.n0 0.000965
R40050 VSS.n4508 VSS.n1 0.000965
R40051 VSS.n4438 VSS.n1 0.000965
R40052 VSS.n4439 VSS.n4438 0.000965
R40053 VSS.n4439 VSS.n4436 0.000965
R40054 VSS.n4443 VSS.n4436 0.000965
R40055 VSS.n4444 VSS.n4443 0.000965
R40056 VSS.n4445 VSS.n4444 0.000965
R40057 VSS.n4445 VSS.n4434 0.000965
R40058 VSS.n4449 VSS.n4434 0.000965
R40059 VSS.n4450 VSS.n4449 0.000965
R40060 VSS.n4451 VSS.n4450 0.000965
R40061 VSS.n4451 VSS.n4432 0.000965
R40062 VSS.n4455 VSS.n4432 0.000965
R40063 VSS.n4456 VSS.n4455 0.000965
R40064 VSS.n4457 VSS.n4456 0.000965
R40065 VSS.n4457 VSS.n4430 0.000965
R40066 VSS.n4461 VSS.n4430 0.000965
R40067 VSS.n4462 VSS.n4461 0.000965
R40068 VSS.n4463 VSS.n4462 0.000965
R40069 VSS.n4463 VSS.n4428 0.000965
R40070 VSS.n4467 VSS.n4428 0.000965
R40071 VSS.n4468 VSS.n4467 0.000965
R40072 VSS.n4469 VSS.n4468 0.000965
R40073 VSS.n4469 VSS.n4426 0.000965
R40074 VSS.n4473 VSS.n4426 0.000965
R40075 VSS.n4474 VSS.n4473 0.000965
R40076 VSS.n4475 VSS.n4474 0.000965
R40077 VSS.n4475 VSS.n4424 0.000965
R40078 VSS.n4479 VSS.n4424 0.000965
R40079 VSS.n4480 VSS.n4479 0.000965
R40080 VSS.n4481 VSS.n4480 0.000965
R40081 VSS.n4481 VSS.n4422 0.000965
R40082 VSS.n4485 VSS.n4422 0.000965
R40083 VSS.n4486 VSS.n4485 0.000965
R40084 VSS.n4487 VSS.n4486 0.000965
R40085 VSS.n4487 VSS.n4420 0.000965
R40086 VSS.n4491 VSS.n4420 0.000965
R40087 VSS.n4492 VSS.n4491 0.000965
R40088 VSS.n4493 VSS.n4492 0.000965
R40089 VSS.n4493 VSS.n4418 0.000965
R40090 VSS.n4497 VSS.n4418 0.000965
R40091 VSS.n4498 VSS.n4497 0.000965
R40092 VSS.n4499 VSS.n4498 0.000965
R40093 VSS.n3049 VSS.n2481 0.000965
R40094 VSS.n3045 VSS.n2481 0.000965
R40095 VSS.n3045 VSS.n3044 0.000965
R40096 VSS.n3044 VSS.n3043 0.000965
R40097 VSS.n3043 VSS.n2488 0.000965
R40098 VSS.n3039 VSS.n2488 0.000965
R40099 VSS.n3039 VSS.n3038 0.000965
R40100 VSS.n3038 VSS.n3037 0.000965
R40101 VSS.n3037 VSS.n2496 0.000965
R40102 VSS.n3033 VSS.n2496 0.000965
R40103 VSS.n3033 VSS.n3032 0.000965
R40104 VSS.n3032 VSS.n3031 0.000965
R40105 VSS.n3031 VSS.n2504 0.000965
R40106 VSS.n3027 VSS.n2504 0.000965
R40107 VSS.n3027 VSS.n3026 0.000965
R40108 VSS.n3026 VSS.n3025 0.000965
R40109 VSS.n3025 VSS.n2512 0.000965
R40110 VSS.n3021 VSS.n2512 0.000965
R40111 VSS.n3021 VSS.n3020 0.000965
R40112 VSS.n3020 VSS.n3019 0.000965
R40113 VSS.n3019 VSS.n2520 0.000965
R40114 VSS.n3015 VSS.n2520 0.000965
R40115 VSS.n3015 VSS.n3014 0.000965
R40116 VSS.n3014 VSS.n3013 0.000965
R40117 VSS.n3013 VSS.n2528 0.000965
R40118 VSS.n3009 VSS.n2528 0.000965
R40119 VSS.n3009 VSS.n3008 0.000965
R40120 VSS.n3008 VSS.n3007 0.000965
R40121 VSS.n3007 VSS.n2536 0.000965
R40122 VSS.n3003 VSS.n2536 0.000965
R40123 VSS.n3003 VSS.n3002 0.000965
R40124 VSS.n3002 VSS.n3001 0.000965
R40125 VSS.n3001 VSS.n2544 0.000965
R40126 VSS.n2997 VSS.n2544 0.000965
R40127 VSS.n2997 VSS.n2996 0.000965
R40128 VSS.n2996 VSS.n2995 0.000965
R40129 VSS.n2995 VSS.n2552 0.000965
R40130 VSS.n2991 VSS.n2552 0.000965
R40131 VSS.n2991 VSS.n2990 0.000965
R40132 VSS.n2990 VSS.n2989 0.000965
R40133 VSS.n2989 VSS.n2560 0.000965
R40134 VSS.n2985 VSS.n2560 0.000965
R40135 VSS.n2985 VSS.n2984 0.000965
R40136 VSS.n2984 VSS.n2983 0.000965
R40137 VSS.n2983 VSS.n2568 0.000965
R40138 VSS.n2979 VSS.n2568 0.000965
R40139 VSS.n2979 VSS.n2978 0.000965
R40140 VSS.n2978 VSS.n2977 0.000965
R40141 VSS.n2977 VSS.n2576 0.000965
R40142 VSS.n2973 VSS.n2576 0.000965
R40143 VSS.n2973 VSS.n2972 0.000965
R40144 VSS.n2972 VSS.n2971 0.000965
R40145 VSS.n2971 VSS.n2584 0.000965
R40146 VSS.n2967 VSS.n2584 0.000965
R40147 VSS.n2967 VSS.n2966 0.000965
R40148 VSS.n2966 VSS.n2965 0.000965
R40149 VSS.n2965 VSS.n2592 0.000965
R40150 VSS.n2961 VSS.n2592 0.000965
R40151 VSS.n2961 VSS.n2960 0.000965
R40152 VSS.n2960 VSS.n2959 0.000965
R40153 VSS.n2959 VSS.n2600 0.000965
R40154 VSS.n2955 VSS.n2600 0.000965
R40155 VSS.n2955 VSS.n2954 0.000965
R40156 VSS.n2954 VSS.n2953 0.000965
R40157 VSS.n2953 VSS.n2608 0.000965
R40158 VSS.n2949 VSS.n2608 0.000965
R40159 VSS.n2949 VSS.n2948 0.000965
R40160 VSS.n2948 VSS.n2947 0.000965
R40161 VSS.n2947 VSS.n2616 0.000965
R40162 VSS.n2943 VSS.n2616 0.000965
R40163 VSS.n2943 VSS.n2942 0.000965
R40164 VSS.n2942 VSS.n2941 0.000965
R40165 VSS.n2941 VSS.n2624 0.000965
R40166 VSS.n2937 VSS.n2624 0.000965
R40167 VSS.n2937 VSS.n2936 0.000965
R40168 VSS.n2936 VSS.n2935 0.000965
R40169 VSS.n2935 VSS.n2632 0.000965
R40170 VSS.n2931 VSS.n2632 0.000965
R40171 VSS.n2931 VSS.n2930 0.000965
R40172 VSS.n2930 VSS.n2929 0.000965
R40173 VSS.n2926 VSS.n2925 0.000965
R40174 VSS.n2925 VSS.n2924 0.000965
R40175 VSS.n2924 VSS.n2647 0.000965
R40176 VSS.n2920 VSS.n2647 0.000965
R40177 VSS.n2920 VSS.n2919 0.000965
R40178 VSS.n2919 VSS.n2918 0.000965
R40179 VSS.n2918 VSS.n2655 0.000965
R40180 VSS.n2914 VSS.n2655 0.000965
R40181 VSS.n2914 VSS.n2913 0.000965
R40182 VSS.n2913 VSS.n2912 0.000965
R40183 VSS.n2912 VSS.n2663 0.000965
R40184 VSS.n2908 VSS.n2663 0.000965
R40185 VSS.n2908 VSS.n2907 0.000965
R40186 VSS.n2907 VSS.n2906 0.000965
R40187 VSS.n2906 VSS.n2671 0.000965
R40188 VSS.n2902 VSS.n2671 0.000965
R40189 VSS.n2902 VSS.n2901 0.000965
R40190 VSS.n2901 VSS.n2900 0.000965
R40191 VSS.n2900 VSS.n2679 0.000965
R40192 VSS.n2896 VSS.n2679 0.000965
R40193 VSS.n2896 VSS.n2895 0.000965
R40194 VSS.n2895 VSS.n2894 0.000965
R40195 VSS.n2894 VSS.n2687 0.000965
R40196 VSS.n2890 VSS.n2687 0.000965
R40197 VSS.n2890 VSS.n2889 0.000965
R40198 VSS.n2889 VSS.n2888 0.000965
R40199 VSS.n2888 VSS.n2695 0.000965
R40200 VSS.n2884 VSS.n2695 0.000965
R40201 VSS.n2884 VSS.n2883 0.000965
R40202 VSS.n2883 VSS.n2882 0.000965
R40203 VSS.n2882 VSS.n2703 0.000965
R40204 VSS.n2878 VSS.n2703 0.000965
R40205 VSS.n2878 VSS.n2877 0.000965
R40206 VSS.n2877 VSS.n2876 0.000965
R40207 VSS.n2876 VSS.n2711 0.000965
R40208 VSS.n2872 VSS.n2711 0.000965
R40209 VSS.n2872 VSS.n2871 0.000965
R40210 VSS.n2871 VSS.n2870 0.000965
R40211 VSS.n2870 VSS.n2719 0.000965
R40212 VSS.n2866 VSS.n2719 0.000965
R40213 VSS.n2866 VSS.n2865 0.000965
R40214 VSS.n2865 VSS.n2864 0.000965
R40215 VSS.n2864 VSS.n2727 0.000965
R40216 VSS VSS.n0 0.00089
R40217 VSS.n2929 VSS 0.00089
R40218 VSS VSS.n4508 0.000575
R40219 VSS.n2926 VSS 0.000575
R40220 a_n1924_n43526.n1 a_n1924_n43526.t5 45.8581
R40221 a_n1924_n43526.n1 a_n1924_n43526.t4 45.8463
R40222 a_n1924_n43526.n1 a_n1924_n43526.t7 45.5929
R40223 a_n1924_n43526.n2 a_n1924_n43526.t2 45.5905
R40224 a_n1924_n43526.n1 a_n1924_n43526.t6 45.5905
R40225 a_n1924_n43526.n0 a_n1924_n43526.t1 9.52626
R40226 a_n1924_n43526.n2 a_n1924_n43526.t3 9.36673
R40227 a_n1924_n43526.n0 a_n1924_n43526.n1 9.34387
R40228 a_n1924_n43526.t0 a_n1924_n43526.n0 9.32226
R40229 a_n1924_n43526.n0 a_n1924_n43526.n2 4.41355
R40230 a_16582_n43566.t1 a_16582_n43566.n0 8.35926
R40231 a_16582_n43566.n0 a_16582_n43566.t0 8.19126
R40232 a_16582_n43566.n0 a_16582_n43566.t2 0.891842
R40233 VINP.n67 VINP.t14 41.7352
R40234 VINP.n67 VINP.t9 41.638
R40235 VINP.n68 VINP.t17 41.638
R40236 VINP.n69 VINP.t1 41.638
R40237 VINP.n70 VINP.t8 41.638
R40238 VINP.n71 VINP.t3 41.638
R40239 VINP.n72 VINP.t16 41.638
R40240 VINP.n73 VINP.t11 41.638
R40241 VINP.n74 VINP.t4 41.638
R40242 VINP.n75 VINP.t13 41.638
R40243 VINP.n76 VINP.t7 41.638
R40244 VINP.n77 VINP.t2 41.638
R40245 VINP.n78 VINP.t18 41.638
R40246 VINP.n79 VINP.t12 41.638
R40247 VINP.n80 VINP.t0 41.638
R40248 VINP.n81 VINP.t15 41.638
R40249 VINP.n82 VINP.t10 41.638
R40250 VINP.n83 VINP.t5 41.638
R40251 VINP.n84 VINP.t19 41.638
R40252 VINP.n85 VINP.t6 41.638
R40253 VINP.n86 VINP.n85 10.0188
R40254 VINP.n276 VINP.n151 4.5005
R40255 VINP.n656 VINP.n151 4.5005
R40256 VINP.n151 VINP.n0 4.5005
R40257 VINP.n280 VINP.n149 4.5005
R40258 VINP.n275 VINP.n149 4.5005
R40259 VINP.n282 VINP.n149 4.5005
R40260 VINP.n274 VINP.n149 4.5005
R40261 VINP.n284 VINP.n149 4.5005
R40262 VINP.n273 VINP.n149 4.5005
R40263 VINP.n286 VINP.n149 4.5005
R40264 VINP.n272 VINP.n149 4.5005
R40265 VINP.n288 VINP.n149 4.5005
R40266 VINP.n271 VINP.n149 4.5005
R40267 VINP.n290 VINP.n149 4.5005
R40268 VINP.n270 VINP.n149 4.5005
R40269 VINP.n292 VINP.n149 4.5005
R40270 VINP.n269 VINP.n149 4.5005
R40271 VINP.n294 VINP.n149 4.5005
R40272 VINP.n268 VINP.n149 4.5005
R40273 VINP.n296 VINP.n149 4.5005
R40274 VINP.n267 VINP.n149 4.5005
R40275 VINP.n298 VINP.n149 4.5005
R40276 VINP.n266 VINP.n149 4.5005
R40277 VINP.n300 VINP.n149 4.5005
R40278 VINP.n265 VINP.n149 4.5005
R40279 VINP.n302 VINP.n149 4.5005
R40280 VINP.n264 VINP.n149 4.5005
R40281 VINP.n304 VINP.n149 4.5005
R40282 VINP.n263 VINP.n149 4.5005
R40283 VINP.n306 VINP.n149 4.5005
R40284 VINP.n262 VINP.n149 4.5005
R40285 VINP.n308 VINP.n149 4.5005
R40286 VINP.n261 VINP.n149 4.5005
R40287 VINP.n310 VINP.n149 4.5005
R40288 VINP.n260 VINP.n149 4.5005
R40289 VINP.n312 VINP.n149 4.5005
R40290 VINP.n259 VINP.n149 4.5005
R40291 VINP.n314 VINP.n149 4.5005
R40292 VINP.n258 VINP.n149 4.5005
R40293 VINP.n316 VINP.n149 4.5005
R40294 VINP.n257 VINP.n149 4.5005
R40295 VINP.n318 VINP.n149 4.5005
R40296 VINP.n256 VINP.n149 4.5005
R40297 VINP.n320 VINP.n149 4.5005
R40298 VINP.n255 VINP.n149 4.5005
R40299 VINP.n322 VINP.n149 4.5005
R40300 VINP.n254 VINP.n149 4.5005
R40301 VINP.n324 VINP.n149 4.5005
R40302 VINP.n253 VINP.n149 4.5005
R40303 VINP.n326 VINP.n149 4.5005
R40304 VINP.n252 VINP.n149 4.5005
R40305 VINP.n328 VINP.n149 4.5005
R40306 VINP.n251 VINP.n149 4.5005
R40307 VINP.n330 VINP.n149 4.5005
R40308 VINP.n250 VINP.n149 4.5005
R40309 VINP.n332 VINP.n149 4.5005
R40310 VINP.n249 VINP.n149 4.5005
R40311 VINP.n334 VINP.n149 4.5005
R40312 VINP.n248 VINP.n149 4.5005
R40313 VINP.n336 VINP.n149 4.5005
R40314 VINP.n247 VINP.n149 4.5005
R40315 VINP.n338 VINP.n149 4.5005
R40316 VINP.n246 VINP.n149 4.5005
R40317 VINP.n340 VINP.n149 4.5005
R40318 VINP.n245 VINP.n149 4.5005
R40319 VINP.n342 VINP.n149 4.5005
R40320 VINP.n244 VINP.n149 4.5005
R40321 VINP.n344 VINP.n149 4.5005
R40322 VINP.n243 VINP.n149 4.5005
R40323 VINP.n346 VINP.n149 4.5005
R40324 VINP.n242 VINP.n149 4.5005
R40325 VINP.n348 VINP.n149 4.5005
R40326 VINP.n241 VINP.n149 4.5005
R40327 VINP.n350 VINP.n149 4.5005
R40328 VINP.n240 VINP.n149 4.5005
R40329 VINP.n352 VINP.n149 4.5005
R40330 VINP.n239 VINP.n149 4.5005
R40331 VINP.n354 VINP.n149 4.5005
R40332 VINP.n238 VINP.n149 4.5005
R40333 VINP.n356 VINP.n149 4.5005
R40334 VINP.n237 VINP.n149 4.5005
R40335 VINP.n358 VINP.n149 4.5005
R40336 VINP.n236 VINP.n149 4.5005
R40337 VINP.n360 VINP.n149 4.5005
R40338 VINP.n235 VINP.n149 4.5005
R40339 VINP.n362 VINP.n149 4.5005
R40340 VINP.n234 VINP.n149 4.5005
R40341 VINP.n364 VINP.n149 4.5005
R40342 VINP.n233 VINP.n149 4.5005
R40343 VINP.n366 VINP.n149 4.5005
R40344 VINP.n232 VINP.n149 4.5005
R40345 VINP.n368 VINP.n149 4.5005
R40346 VINP.n231 VINP.n149 4.5005
R40347 VINP.n370 VINP.n149 4.5005
R40348 VINP.n230 VINP.n149 4.5005
R40349 VINP.n372 VINP.n149 4.5005
R40350 VINP.n229 VINP.n149 4.5005
R40351 VINP.n374 VINP.n149 4.5005
R40352 VINP.n228 VINP.n149 4.5005
R40353 VINP.n376 VINP.n149 4.5005
R40354 VINP.n227 VINP.n149 4.5005
R40355 VINP.n378 VINP.n149 4.5005
R40356 VINP.n226 VINP.n149 4.5005
R40357 VINP.n380 VINP.n149 4.5005
R40358 VINP.n225 VINP.n149 4.5005
R40359 VINP.n382 VINP.n149 4.5005
R40360 VINP.n224 VINP.n149 4.5005
R40361 VINP.n384 VINP.n149 4.5005
R40362 VINP.n223 VINP.n149 4.5005
R40363 VINP.n386 VINP.n149 4.5005
R40364 VINP.n222 VINP.n149 4.5005
R40365 VINP.n388 VINP.n149 4.5005
R40366 VINP.n221 VINP.n149 4.5005
R40367 VINP.n390 VINP.n149 4.5005
R40368 VINP.n220 VINP.n149 4.5005
R40369 VINP.n392 VINP.n149 4.5005
R40370 VINP.n219 VINP.n149 4.5005
R40371 VINP.n394 VINP.n149 4.5005
R40372 VINP.n218 VINP.n149 4.5005
R40373 VINP.n396 VINP.n149 4.5005
R40374 VINP.n217 VINP.n149 4.5005
R40375 VINP.n398 VINP.n149 4.5005
R40376 VINP.n216 VINP.n149 4.5005
R40377 VINP.n400 VINP.n149 4.5005
R40378 VINP.n215 VINP.n149 4.5005
R40379 VINP.n654 VINP.n149 4.5005
R40380 VINP.n656 VINP.n149 4.5005
R40381 VINP.n149 VINP.n0 4.5005
R40382 VINP.n278 VINP.n152 4.5005
R40383 VINP.n276 VINP.n152 4.5005
R40384 VINP.n280 VINP.n152 4.5005
R40385 VINP.n275 VINP.n152 4.5005
R40386 VINP.n282 VINP.n152 4.5005
R40387 VINP.n274 VINP.n152 4.5005
R40388 VINP.n284 VINP.n152 4.5005
R40389 VINP.n273 VINP.n152 4.5005
R40390 VINP.n286 VINP.n152 4.5005
R40391 VINP.n272 VINP.n152 4.5005
R40392 VINP.n288 VINP.n152 4.5005
R40393 VINP.n271 VINP.n152 4.5005
R40394 VINP.n290 VINP.n152 4.5005
R40395 VINP.n270 VINP.n152 4.5005
R40396 VINP.n292 VINP.n152 4.5005
R40397 VINP.n269 VINP.n152 4.5005
R40398 VINP.n294 VINP.n152 4.5005
R40399 VINP.n268 VINP.n152 4.5005
R40400 VINP.n296 VINP.n152 4.5005
R40401 VINP.n267 VINP.n152 4.5005
R40402 VINP.n298 VINP.n152 4.5005
R40403 VINP.n266 VINP.n152 4.5005
R40404 VINP.n300 VINP.n152 4.5005
R40405 VINP.n265 VINP.n152 4.5005
R40406 VINP.n302 VINP.n152 4.5005
R40407 VINP.n264 VINP.n152 4.5005
R40408 VINP.n304 VINP.n152 4.5005
R40409 VINP.n263 VINP.n152 4.5005
R40410 VINP.n306 VINP.n152 4.5005
R40411 VINP.n262 VINP.n152 4.5005
R40412 VINP.n308 VINP.n152 4.5005
R40413 VINP.n261 VINP.n152 4.5005
R40414 VINP.n310 VINP.n152 4.5005
R40415 VINP.n260 VINP.n152 4.5005
R40416 VINP.n312 VINP.n152 4.5005
R40417 VINP.n259 VINP.n152 4.5005
R40418 VINP.n314 VINP.n152 4.5005
R40419 VINP.n258 VINP.n152 4.5005
R40420 VINP.n316 VINP.n152 4.5005
R40421 VINP.n257 VINP.n152 4.5005
R40422 VINP.n318 VINP.n152 4.5005
R40423 VINP.n256 VINP.n152 4.5005
R40424 VINP.n320 VINP.n152 4.5005
R40425 VINP.n255 VINP.n152 4.5005
R40426 VINP.n322 VINP.n152 4.5005
R40427 VINP.n254 VINP.n152 4.5005
R40428 VINP.n324 VINP.n152 4.5005
R40429 VINP.n253 VINP.n152 4.5005
R40430 VINP.n326 VINP.n152 4.5005
R40431 VINP.n252 VINP.n152 4.5005
R40432 VINP.n328 VINP.n152 4.5005
R40433 VINP.n251 VINP.n152 4.5005
R40434 VINP.n330 VINP.n152 4.5005
R40435 VINP.n250 VINP.n152 4.5005
R40436 VINP.n332 VINP.n152 4.5005
R40437 VINP.n249 VINP.n152 4.5005
R40438 VINP.n334 VINP.n152 4.5005
R40439 VINP.n248 VINP.n152 4.5005
R40440 VINP.n336 VINP.n152 4.5005
R40441 VINP.n247 VINP.n152 4.5005
R40442 VINP.n338 VINP.n152 4.5005
R40443 VINP.n246 VINP.n152 4.5005
R40444 VINP.n340 VINP.n152 4.5005
R40445 VINP.n245 VINP.n152 4.5005
R40446 VINP.n342 VINP.n152 4.5005
R40447 VINP.n244 VINP.n152 4.5005
R40448 VINP.n344 VINP.n152 4.5005
R40449 VINP.n243 VINP.n152 4.5005
R40450 VINP.n346 VINP.n152 4.5005
R40451 VINP.n242 VINP.n152 4.5005
R40452 VINP.n348 VINP.n152 4.5005
R40453 VINP.n241 VINP.n152 4.5005
R40454 VINP.n350 VINP.n152 4.5005
R40455 VINP.n240 VINP.n152 4.5005
R40456 VINP.n352 VINP.n152 4.5005
R40457 VINP.n239 VINP.n152 4.5005
R40458 VINP.n354 VINP.n152 4.5005
R40459 VINP.n238 VINP.n152 4.5005
R40460 VINP.n356 VINP.n152 4.5005
R40461 VINP.n237 VINP.n152 4.5005
R40462 VINP.n358 VINP.n152 4.5005
R40463 VINP.n236 VINP.n152 4.5005
R40464 VINP.n360 VINP.n152 4.5005
R40465 VINP.n235 VINP.n152 4.5005
R40466 VINP.n362 VINP.n152 4.5005
R40467 VINP.n234 VINP.n152 4.5005
R40468 VINP.n364 VINP.n152 4.5005
R40469 VINP.n233 VINP.n152 4.5005
R40470 VINP.n366 VINP.n152 4.5005
R40471 VINP.n232 VINP.n152 4.5005
R40472 VINP.n368 VINP.n152 4.5005
R40473 VINP.n231 VINP.n152 4.5005
R40474 VINP.n370 VINP.n152 4.5005
R40475 VINP.n230 VINP.n152 4.5005
R40476 VINP.n372 VINP.n152 4.5005
R40477 VINP.n229 VINP.n152 4.5005
R40478 VINP.n374 VINP.n152 4.5005
R40479 VINP.n228 VINP.n152 4.5005
R40480 VINP.n376 VINP.n152 4.5005
R40481 VINP.n227 VINP.n152 4.5005
R40482 VINP.n378 VINP.n152 4.5005
R40483 VINP.n226 VINP.n152 4.5005
R40484 VINP.n380 VINP.n152 4.5005
R40485 VINP.n225 VINP.n152 4.5005
R40486 VINP.n382 VINP.n152 4.5005
R40487 VINP.n224 VINP.n152 4.5005
R40488 VINP.n384 VINP.n152 4.5005
R40489 VINP.n223 VINP.n152 4.5005
R40490 VINP.n386 VINP.n152 4.5005
R40491 VINP.n222 VINP.n152 4.5005
R40492 VINP.n388 VINP.n152 4.5005
R40493 VINP.n221 VINP.n152 4.5005
R40494 VINP.n390 VINP.n152 4.5005
R40495 VINP.n220 VINP.n152 4.5005
R40496 VINP.n392 VINP.n152 4.5005
R40497 VINP.n219 VINP.n152 4.5005
R40498 VINP.n394 VINP.n152 4.5005
R40499 VINP.n218 VINP.n152 4.5005
R40500 VINP.n396 VINP.n152 4.5005
R40501 VINP.n217 VINP.n152 4.5005
R40502 VINP.n398 VINP.n152 4.5005
R40503 VINP.n216 VINP.n152 4.5005
R40504 VINP.n400 VINP.n152 4.5005
R40505 VINP.n215 VINP.n152 4.5005
R40506 VINP.n654 VINP.n152 4.5005
R40507 VINP.n656 VINP.n152 4.5005
R40508 VINP.n152 VINP.n0 4.5005
R40509 VINP.n278 VINP.n148 4.5005
R40510 VINP.n276 VINP.n148 4.5005
R40511 VINP.n280 VINP.n148 4.5005
R40512 VINP.n275 VINP.n148 4.5005
R40513 VINP.n282 VINP.n148 4.5005
R40514 VINP.n274 VINP.n148 4.5005
R40515 VINP.n284 VINP.n148 4.5005
R40516 VINP.n273 VINP.n148 4.5005
R40517 VINP.n286 VINP.n148 4.5005
R40518 VINP.n272 VINP.n148 4.5005
R40519 VINP.n288 VINP.n148 4.5005
R40520 VINP.n271 VINP.n148 4.5005
R40521 VINP.n290 VINP.n148 4.5005
R40522 VINP.n270 VINP.n148 4.5005
R40523 VINP.n292 VINP.n148 4.5005
R40524 VINP.n269 VINP.n148 4.5005
R40525 VINP.n294 VINP.n148 4.5005
R40526 VINP.n268 VINP.n148 4.5005
R40527 VINP.n296 VINP.n148 4.5005
R40528 VINP.n267 VINP.n148 4.5005
R40529 VINP.n298 VINP.n148 4.5005
R40530 VINP.n266 VINP.n148 4.5005
R40531 VINP.n300 VINP.n148 4.5005
R40532 VINP.n265 VINP.n148 4.5005
R40533 VINP.n302 VINP.n148 4.5005
R40534 VINP.n264 VINP.n148 4.5005
R40535 VINP.n304 VINP.n148 4.5005
R40536 VINP.n263 VINP.n148 4.5005
R40537 VINP.n306 VINP.n148 4.5005
R40538 VINP.n262 VINP.n148 4.5005
R40539 VINP.n308 VINP.n148 4.5005
R40540 VINP.n261 VINP.n148 4.5005
R40541 VINP.n310 VINP.n148 4.5005
R40542 VINP.n260 VINP.n148 4.5005
R40543 VINP.n312 VINP.n148 4.5005
R40544 VINP.n259 VINP.n148 4.5005
R40545 VINP.n314 VINP.n148 4.5005
R40546 VINP.n258 VINP.n148 4.5005
R40547 VINP.n316 VINP.n148 4.5005
R40548 VINP.n257 VINP.n148 4.5005
R40549 VINP.n318 VINP.n148 4.5005
R40550 VINP.n256 VINP.n148 4.5005
R40551 VINP.n320 VINP.n148 4.5005
R40552 VINP.n255 VINP.n148 4.5005
R40553 VINP.n322 VINP.n148 4.5005
R40554 VINP.n254 VINP.n148 4.5005
R40555 VINP.n324 VINP.n148 4.5005
R40556 VINP.n253 VINP.n148 4.5005
R40557 VINP.n326 VINP.n148 4.5005
R40558 VINP.n252 VINP.n148 4.5005
R40559 VINP.n328 VINP.n148 4.5005
R40560 VINP.n251 VINP.n148 4.5005
R40561 VINP.n330 VINP.n148 4.5005
R40562 VINP.n250 VINP.n148 4.5005
R40563 VINP.n332 VINP.n148 4.5005
R40564 VINP.n249 VINP.n148 4.5005
R40565 VINP.n334 VINP.n148 4.5005
R40566 VINP.n248 VINP.n148 4.5005
R40567 VINP.n336 VINP.n148 4.5005
R40568 VINP.n247 VINP.n148 4.5005
R40569 VINP.n338 VINP.n148 4.5005
R40570 VINP.n246 VINP.n148 4.5005
R40571 VINP.n340 VINP.n148 4.5005
R40572 VINP.n245 VINP.n148 4.5005
R40573 VINP.n342 VINP.n148 4.5005
R40574 VINP.n244 VINP.n148 4.5005
R40575 VINP.n344 VINP.n148 4.5005
R40576 VINP.n243 VINP.n148 4.5005
R40577 VINP.n346 VINP.n148 4.5005
R40578 VINP.n242 VINP.n148 4.5005
R40579 VINP.n348 VINP.n148 4.5005
R40580 VINP.n241 VINP.n148 4.5005
R40581 VINP.n350 VINP.n148 4.5005
R40582 VINP.n240 VINP.n148 4.5005
R40583 VINP.n352 VINP.n148 4.5005
R40584 VINP.n239 VINP.n148 4.5005
R40585 VINP.n354 VINP.n148 4.5005
R40586 VINP.n238 VINP.n148 4.5005
R40587 VINP.n356 VINP.n148 4.5005
R40588 VINP.n237 VINP.n148 4.5005
R40589 VINP.n358 VINP.n148 4.5005
R40590 VINP.n236 VINP.n148 4.5005
R40591 VINP.n360 VINP.n148 4.5005
R40592 VINP.n235 VINP.n148 4.5005
R40593 VINP.n362 VINP.n148 4.5005
R40594 VINP.n234 VINP.n148 4.5005
R40595 VINP.n364 VINP.n148 4.5005
R40596 VINP.n233 VINP.n148 4.5005
R40597 VINP.n366 VINP.n148 4.5005
R40598 VINP.n232 VINP.n148 4.5005
R40599 VINP.n368 VINP.n148 4.5005
R40600 VINP.n231 VINP.n148 4.5005
R40601 VINP.n370 VINP.n148 4.5005
R40602 VINP.n230 VINP.n148 4.5005
R40603 VINP.n372 VINP.n148 4.5005
R40604 VINP.n229 VINP.n148 4.5005
R40605 VINP.n374 VINP.n148 4.5005
R40606 VINP.n228 VINP.n148 4.5005
R40607 VINP.n376 VINP.n148 4.5005
R40608 VINP.n227 VINP.n148 4.5005
R40609 VINP.n378 VINP.n148 4.5005
R40610 VINP.n226 VINP.n148 4.5005
R40611 VINP.n380 VINP.n148 4.5005
R40612 VINP.n225 VINP.n148 4.5005
R40613 VINP.n382 VINP.n148 4.5005
R40614 VINP.n224 VINP.n148 4.5005
R40615 VINP.n384 VINP.n148 4.5005
R40616 VINP.n223 VINP.n148 4.5005
R40617 VINP.n386 VINP.n148 4.5005
R40618 VINP.n222 VINP.n148 4.5005
R40619 VINP.n388 VINP.n148 4.5005
R40620 VINP.n221 VINP.n148 4.5005
R40621 VINP.n390 VINP.n148 4.5005
R40622 VINP.n220 VINP.n148 4.5005
R40623 VINP.n392 VINP.n148 4.5005
R40624 VINP.n219 VINP.n148 4.5005
R40625 VINP.n394 VINP.n148 4.5005
R40626 VINP.n218 VINP.n148 4.5005
R40627 VINP.n396 VINP.n148 4.5005
R40628 VINP.n217 VINP.n148 4.5005
R40629 VINP.n398 VINP.n148 4.5005
R40630 VINP.n216 VINP.n148 4.5005
R40631 VINP.n400 VINP.n148 4.5005
R40632 VINP.n215 VINP.n148 4.5005
R40633 VINP.n654 VINP.n148 4.5005
R40634 VINP.n656 VINP.n148 4.5005
R40635 VINP.n148 VINP.n0 4.5005
R40636 VINP.n278 VINP.n153 4.5005
R40637 VINP.n276 VINP.n153 4.5005
R40638 VINP.n280 VINP.n153 4.5005
R40639 VINP.n275 VINP.n153 4.5005
R40640 VINP.n282 VINP.n153 4.5005
R40641 VINP.n274 VINP.n153 4.5005
R40642 VINP.n284 VINP.n153 4.5005
R40643 VINP.n273 VINP.n153 4.5005
R40644 VINP.n286 VINP.n153 4.5005
R40645 VINP.n272 VINP.n153 4.5005
R40646 VINP.n288 VINP.n153 4.5005
R40647 VINP.n271 VINP.n153 4.5005
R40648 VINP.n290 VINP.n153 4.5005
R40649 VINP.n270 VINP.n153 4.5005
R40650 VINP.n292 VINP.n153 4.5005
R40651 VINP.n269 VINP.n153 4.5005
R40652 VINP.n294 VINP.n153 4.5005
R40653 VINP.n268 VINP.n153 4.5005
R40654 VINP.n296 VINP.n153 4.5005
R40655 VINP.n267 VINP.n153 4.5005
R40656 VINP.n298 VINP.n153 4.5005
R40657 VINP.n266 VINP.n153 4.5005
R40658 VINP.n300 VINP.n153 4.5005
R40659 VINP.n265 VINP.n153 4.5005
R40660 VINP.n302 VINP.n153 4.5005
R40661 VINP.n264 VINP.n153 4.5005
R40662 VINP.n304 VINP.n153 4.5005
R40663 VINP.n263 VINP.n153 4.5005
R40664 VINP.n306 VINP.n153 4.5005
R40665 VINP.n262 VINP.n153 4.5005
R40666 VINP.n308 VINP.n153 4.5005
R40667 VINP.n261 VINP.n153 4.5005
R40668 VINP.n310 VINP.n153 4.5005
R40669 VINP.n260 VINP.n153 4.5005
R40670 VINP.n312 VINP.n153 4.5005
R40671 VINP.n259 VINP.n153 4.5005
R40672 VINP.n314 VINP.n153 4.5005
R40673 VINP.n258 VINP.n153 4.5005
R40674 VINP.n316 VINP.n153 4.5005
R40675 VINP.n257 VINP.n153 4.5005
R40676 VINP.n318 VINP.n153 4.5005
R40677 VINP.n256 VINP.n153 4.5005
R40678 VINP.n320 VINP.n153 4.5005
R40679 VINP.n255 VINP.n153 4.5005
R40680 VINP.n322 VINP.n153 4.5005
R40681 VINP.n254 VINP.n153 4.5005
R40682 VINP.n324 VINP.n153 4.5005
R40683 VINP.n253 VINP.n153 4.5005
R40684 VINP.n326 VINP.n153 4.5005
R40685 VINP.n252 VINP.n153 4.5005
R40686 VINP.n328 VINP.n153 4.5005
R40687 VINP.n251 VINP.n153 4.5005
R40688 VINP.n330 VINP.n153 4.5005
R40689 VINP.n250 VINP.n153 4.5005
R40690 VINP.n332 VINP.n153 4.5005
R40691 VINP.n249 VINP.n153 4.5005
R40692 VINP.n334 VINP.n153 4.5005
R40693 VINP.n248 VINP.n153 4.5005
R40694 VINP.n336 VINP.n153 4.5005
R40695 VINP.n247 VINP.n153 4.5005
R40696 VINP.n338 VINP.n153 4.5005
R40697 VINP.n246 VINP.n153 4.5005
R40698 VINP.n340 VINP.n153 4.5005
R40699 VINP.n245 VINP.n153 4.5005
R40700 VINP.n342 VINP.n153 4.5005
R40701 VINP.n244 VINP.n153 4.5005
R40702 VINP.n344 VINP.n153 4.5005
R40703 VINP.n243 VINP.n153 4.5005
R40704 VINP.n346 VINP.n153 4.5005
R40705 VINP.n242 VINP.n153 4.5005
R40706 VINP.n348 VINP.n153 4.5005
R40707 VINP.n241 VINP.n153 4.5005
R40708 VINP.n350 VINP.n153 4.5005
R40709 VINP.n240 VINP.n153 4.5005
R40710 VINP.n352 VINP.n153 4.5005
R40711 VINP.n239 VINP.n153 4.5005
R40712 VINP.n354 VINP.n153 4.5005
R40713 VINP.n238 VINP.n153 4.5005
R40714 VINP.n356 VINP.n153 4.5005
R40715 VINP.n237 VINP.n153 4.5005
R40716 VINP.n358 VINP.n153 4.5005
R40717 VINP.n236 VINP.n153 4.5005
R40718 VINP.n360 VINP.n153 4.5005
R40719 VINP.n235 VINP.n153 4.5005
R40720 VINP.n362 VINP.n153 4.5005
R40721 VINP.n234 VINP.n153 4.5005
R40722 VINP.n364 VINP.n153 4.5005
R40723 VINP.n233 VINP.n153 4.5005
R40724 VINP.n366 VINP.n153 4.5005
R40725 VINP.n232 VINP.n153 4.5005
R40726 VINP.n368 VINP.n153 4.5005
R40727 VINP.n231 VINP.n153 4.5005
R40728 VINP.n370 VINP.n153 4.5005
R40729 VINP.n230 VINP.n153 4.5005
R40730 VINP.n372 VINP.n153 4.5005
R40731 VINP.n229 VINP.n153 4.5005
R40732 VINP.n374 VINP.n153 4.5005
R40733 VINP.n228 VINP.n153 4.5005
R40734 VINP.n376 VINP.n153 4.5005
R40735 VINP.n227 VINP.n153 4.5005
R40736 VINP.n378 VINP.n153 4.5005
R40737 VINP.n226 VINP.n153 4.5005
R40738 VINP.n380 VINP.n153 4.5005
R40739 VINP.n225 VINP.n153 4.5005
R40740 VINP.n382 VINP.n153 4.5005
R40741 VINP.n224 VINP.n153 4.5005
R40742 VINP.n384 VINP.n153 4.5005
R40743 VINP.n223 VINP.n153 4.5005
R40744 VINP.n386 VINP.n153 4.5005
R40745 VINP.n222 VINP.n153 4.5005
R40746 VINP.n388 VINP.n153 4.5005
R40747 VINP.n221 VINP.n153 4.5005
R40748 VINP.n390 VINP.n153 4.5005
R40749 VINP.n220 VINP.n153 4.5005
R40750 VINP.n392 VINP.n153 4.5005
R40751 VINP.n219 VINP.n153 4.5005
R40752 VINP.n394 VINP.n153 4.5005
R40753 VINP.n218 VINP.n153 4.5005
R40754 VINP.n396 VINP.n153 4.5005
R40755 VINP.n217 VINP.n153 4.5005
R40756 VINP.n398 VINP.n153 4.5005
R40757 VINP.n216 VINP.n153 4.5005
R40758 VINP.n400 VINP.n153 4.5005
R40759 VINP.n215 VINP.n153 4.5005
R40760 VINP.n654 VINP.n153 4.5005
R40761 VINP.n656 VINP.n153 4.5005
R40762 VINP.n153 VINP.n0 4.5005
R40763 VINP.n278 VINP.n147 4.5005
R40764 VINP.n276 VINP.n147 4.5005
R40765 VINP.n280 VINP.n147 4.5005
R40766 VINP.n275 VINP.n147 4.5005
R40767 VINP.n282 VINP.n147 4.5005
R40768 VINP.n274 VINP.n147 4.5005
R40769 VINP.n284 VINP.n147 4.5005
R40770 VINP.n273 VINP.n147 4.5005
R40771 VINP.n286 VINP.n147 4.5005
R40772 VINP.n272 VINP.n147 4.5005
R40773 VINP.n288 VINP.n147 4.5005
R40774 VINP.n271 VINP.n147 4.5005
R40775 VINP.n290 VINP.n147 4.5005
R40776 VINP.n270 VINP.n147 4.5005
R40777 VINP.n292 VINP.n147 4.5005
R40778 VINP.n269 VINP.n147 4.5005
R40779 VINP.n294 VINP.n147 4.5005
R40780 VINP.n268 VINP.n147 4.5005
R40781 VINP.n296 VINP.n147 4.5005
R40782 VINP.n267 VINP.n147 4.5005
R40783 VINP.n298 VINP.n147 4.5005
R40784 VINP.n266 VINP.n147 4.5005
R40785 VINP.n300 VINP.n147 4.5005
R40786 VINP.n265 VINP.n147 4.5005
R40787 VINP.n302 VINP.n147 4.5005
R40788 VINP.n264 VINP.n147 4.5005
R40789 VINP.n304 VINP.n147 4.5005
R40790 VINP.n263 VINP.n147 4.5005
R40791 VINP.n306 VINP.n147 4.5005
R40792 VINP.n262 VINP.n147 4.5005
R40793 VINP.n308 VINP.n147 4.5005
R40794 VINP.n261 VINP.n147 4.5005
R40795 VINP.n310 VINP.n147 4.5005
R40796 VINP.n260 VINP.n147 4.5005
R40797 VINP.n312 VINP.n147 4.5005
R40798 VINP.n259 VINP.n147 4.5005
R40799 VINP.n314 VINP.n147 4.5005
R40800 VINP.n258 VINP.n147 4.5005
R40801 VINP.n316 VINP.n147 4.5005
R40802 VINP.n257 VINP.n147 4.5005
R40803 VINP.n318 VINP.n147 4.5005
R40804 VINP.n256 VINP.n147 4.5005
R40805 VINP.n320 VINP.n147 4.5005
R40806 VINP.n255 VINP.n147 4.5005
R40807 VINP.n322 VINP.n147 4.5005
R40808 VINP.n254 VINP.n147 4.5005
R40809 VINP.n324 VINP.n147 4.5005
R40810 VINP.n253 VINP.n147 4.5005
R40811 VINP.n326 VINP.n147 4.5005
R40812 VINP.n252 VINP.n147 4.5005
R40813 VINP.n328 VINP.n147 4.5005
R40814 VINP.n251 VINP.n147 4.5005
R40815 VINP.n330 VINP.n147 4.5005
R40816 VINP.n250 VINP.n147 4.5005
R40817 VINP.n332 VINP.n147 4.5005
R40818 VINP.n249 VINP.n147 4.5005
R40819 VINP.n334 VINP.n147 4.5005
R40820 VINP.n248 VINP.n147 4.5005
R40821 VINP.n336 VINP.n147 4.5005
R40822 VINP.n247 VINP.n147 4.5005
R40823 VINP.n338 VINP.n147 4.5005
R40824 VINP.n246 VINP.n147 4.5005
R40825 VINP.n340 VINP.n147 4.5005
R40826 VINP.n245 VINP.n147 4.5005
R40827 VINP.n342 VINP.n147 4.5005
R40828 VINP.n244 VINP.n147 4.5005
R40829 VINP.n344 VINP.n147 4.5005
R40830 VINP.n243 VINP.n147 4.5005
R40831 VINP.n346 VINP.n147 4.5005
R40832 VINP.n242 VINP.n147 4.5005
R40833 VINP.n348 VINP.n147 4.5005
R40834 VINP.n241 VINP.n147 4.5005
R40835 VINP.n350 VINP.n147 4.5005
R40836 VINP.n240 VINP.n147 4.5005
R40837 VINP.n352 VINP.n147 4.5005
R40838 VINP.n239 VINP.n147 4.5005
R40839 VINP.n354 VINP.n147 4.5005
R40840 VINP.n238 VINP.n147 4.5005
R40841 VINP.n356 VINP.n147 4.5005
R40842 VINP.n237 VINP.n147 4.5005
R40843 VINP.n358 VINP.n147 4.5005
R40844 VINP.n236 VINP.n147 4.5005
R40845 VINP.n360 VINP.n147 4.5005
R40846 VINP.n235 VINP.n147 4.5005
R40847 VINP.n362 VINP.n147 4.5005
R40848 VINP.n234 VINP.n147 4.5005
R40849 VINP.n364 VINP.n147 4.5005
R40850 VINP.n233 VINP.n147 4.5005
R40851 VINP.n366 VINP.n147 4.5005
R40852 VINP.n232 VINP.n147 4.5005
R40853 VINP.n368 VINP.n147 4.5005
R40854 VINP.n231 VINP.n147 4.5005
R40855 VINP.n370 VINP.n147 4.5005
R40856 VINP.n230 VINP.n147 4.5005
R40857 VINP.n372 VINP.n147 4.5005
R40858 VINP.n229 VINP.n147 4.5005
R40859 VINP.n374 VINP.n147 4.5005
R40860 VINP.n228 VINP.n147 4.5005
R40861 VINP.n376 VINP.n147 4.5005
R40862 VINP.n227 VINP.n147 4.5005
R40863 VINP.n378 VINP.n147 4.5005
R40864 VINP.n226 VINP.n147 4.5005
R40865 VINP.n380 VINP.n147 4.5005
R40866 VINP.n225 VINP.n147 4.5005
R40867 VINP.n382 VINP.n147 4.5005
R40868 VINP.n224 VINP.n147 4.5005
R40869 VINP.n384 VINP.n147 4.5005
R40870 VINP.n223 VINP.n147 4.5005
R40871 VINP.n386 VINP.n147 4.5005
R40872 VINP.n222 VINP.n147 4.5005
R40873 VINP.n388 VINP.n147 4.5005
R40874 VINP.n221 VINP.n147 4.5005
R40875 VINP.n390 VINP.n147 4.5005
R40876 VINP.n220 VINP.n147 4.5005
R40877 VINP.n392 VINP.n147 4.5005
R40878 VINP.n219 VINP.n147 4.5005
R40879 VINP.n394 VINP.n147 4.5005
R40880 VINP.n218 VINP.n147 4.5005
R40881 VINP.n396 VINP.n147 4.5005
R40882 VINP.n217 VINP.n147 4.5005
R40883 VINP.n398 VINP.n147 4.5005
R40884 VINP.n216 VINP.n147 4.5005
R40885 VINP.n400 VINP.n147 4.5005
R40886 VINP.n215 VINP.n147 4.5005
R40887 VINP.n654 VINP.n147 4.5005
R40888 VINP.n656 VINP.n147 4.5005
R40889 VINP.n147 VINP.n0 4.5005
R40890 VINP.n278 VINP.n154 4.5005
R40891 VINP.n276 VINP.n154 4.5005
R40892 VINP.n280 VINP.n154 4.5005
R40893 VINP.n275 VINP.n154 4.5005
R40894 VINP.n282 VINP.n154 4.5005
R40895 VINP.n274 VINP.n154 4.5005
R40896 VINP.n284 VINP.n154 4.5005
R40897 VINP.n273 VINP.n154 4.5005
R40898 VINP.n286 VINP.n154 4.5005
R40899 VINP.n272 VINP.n154 4.5005
R40900 VINP.n288 VINP.n154 4.5005
R40901 VINP.n271 VINP.n154 4.5005
R40902 VINP.n290 VINP.n154 4.5005
R40903 VINP.n270 VINP.n154 4.5005
R40904 VINP.n292 VINP.n154 4.5005
R40905 VINP.n269 VINP.n154 4.5005
R40906 VINP.n294 VINP.n154 4.5005
R40907 VINP.n268 VINP.n154 4.5005
R40908 VINP.n296 VINP.n154 4.5005
R40909 VINP.n267 VINP.n154 4.5005
R40910 VINP.n298 VINP.n154 4.5005
R40911 VINP.n266 VINP.n154 4.5005
R40912 VINP.n300 VINP.n154 4.5005
R40913 VINP.n265 VINP.n154 4.5005
R40914 VINP.n302 VINP.n154 4.5005
R40915 VINP.n264 VINP.n154 4.5005
R40916 VINP.n304 VINP.n154 4.5005
R40917 VINP.n263 VINP.n154 4.5005
R40918 VINP.n306 VINP.n154 4.5005
R40919 VINP.n262 VINP.n154 4.5005
R40920 VINP.n308 VINP.n154 4.5005
R40921 VINP.n261 VINP.n154 4.5005
R40922 VINP.n310 VINP.n154 4.5005
R40923 VINP.n260 VINP.n154 4.5005
R40924 VINP.n312 VINP.n154 4.5005
R40925 VINP.n259 VINP.n154 4.5005
R40926 VINP.n314 VINP.n154 4.5005
R40927 VINP.n258 VINP.n154 4.5005
R40928 VINP.n316 VINP.n154 4.5005
R40929 VINP.n257 VINP.n154 4.5005
R40930 VINP.n318 VINP.n154 4.5005
R40931 VINP.n256 VINP.n154 4.5005
R40932 VINP.n320 VINP.n154 4.5005
R40933 VINP.n255 VINP.n154 4.5005
R40934 VINP.n322 VINP.n154 4.5005
R40935 VINP.n254 VINP.n154 4.5005
R40936 VINP.n324 VINP.n154 4.5005
R40937 VINP.n253 VINP.n154 4.5005
R40938 VINP.n326 VINP.n154 4.5005
R40939 VINP.n252 VINP.n154 4.5005
R40940 VINP.n328 VINP.n154 4.5005
R40941 VINP.n251 VINP.n154 4.5005
R40942 VINP.n330 VINP.n154 4.5005
R40943 VINP.n250 VINP.n154 4.5005
R40944 VINP.n332 VINP.n154 4.5005
R40945 VINP.n249 VINP.n154 4.5005
R40946 VINP.n334 VINP.n154 4.5005
R40947 VINP.n248 VINP.n154 4.5005
R40948 VINP.n336 VINP.n154 4.5005
R40949 VINP.n247 VINP.n154 4.5005
R40950 VINP.n338 VINP.n154 4.5005
R40951 VINP.n246 VINP.n154 4.5005
R40952 VINP.n340 VINP.n154 4.5005
R40953 VINP.n245 VINP.n154 4.5005
R40954 VINP.n342 VINP.n154 4.5005
R40955 VINP.n244 VINP.n154 4.5005
R40956 VINP.n344 VINP.n154 4.5005
R40957 VINP.n243 VINP.n154 4.5005
R40958 VINP.n346 VINP.n154 4.5005
R40959 VINP.n242 VINP.n154 4.5005
R40960 VINP.n348 VINP.n154 4.5005
R40961 VINP.n241 VINP.n154 4.5005
R40962 VINP.n350 VINP.n154 4.5005
R40963 VINP.n240 VINP.n154 4.5005
R40964 VINP.n352 VINP.n154 4.5005
R40965 VINP.n239 VINP.n154 4.5005
R40966 VINP.n354 VINP.n154 4.5005
R40967 VINP.n238 VINP.n154 4.5005
R40968 VINP.n356 VINP.n154 4.5005
R40969 VINP.n237 VINP.n154 4.5005
R40970 VINP.n358 VINP.n154 4.5005
R40971 VINP.n236 VINP.n154 4.5005
R40972 VINP.n360 VINP.n154 4.5005
R40973 VINP.n235 VINP.n154 4.5005
R40974 VINP.n362 VINP.n154 4.5005
R40975 VINP.n234 VINP.n154 4.5005
R40976 VINP.n364 VINP.n154 4.5005
R40977 VINP.n233 VINP.n154 4.5005
R40978 VINP.n366 VINP.n154 4.5005
R40979 VINP.n232 VINP.n154 4.5005
R40980 VINP.n368 VINP.n154 4.5005
R40981 VINP.n231 VINP.n154 4.5005
R40982 VINP.n370 VINP.n154 4.5005
R40983 VINP.n230 VINP.n154 4.5005
R40984 VINP.n372 VINP.n154 4.5005
R40985 VINP.n229 VINP.n154 4.5005
R40986 VINP.n374 VINP.n154 4.5005
R40987 VINP.n228 VINP.n154 4.5005
R40988 VINP.n376 VINP.n154 4.5005
R40989 VINP.n227 VINP.n154 4.5005
R40990 VINP.n378 VINP.n154 4.5005
R40991 VINP.n226 VINP.n154 4.5005
R40992 VINP.n380 VINP.n154 4.5005
R40993 VINP.n225 VINP.n154 4.5005
R40994 VINP.n382 VINP.n154 4.5005
R40995 VINP.n224 VINP.n154 4.5005
R40996 VINP.n384 VINP.n154 4.5005
R40997 VINP.n223 VINP.n154 4.5005
R40998 VINP.n386 VINP.n154 4.5005
R40999 VINP.n222 VINP.n154 4.5005
R41000 VINP.n388 VINP.n154 4.5005
R41001 VINP.n221 VINP.n154 4.5005
R41002 VINP.n390 VINP.n154 4.5005
R41003 VINP.n220 VINP.n154 4.5005
R41004 VINP.n392 VINP.n154 4.5005
R41005 VINP.n219 VINP.n154 4.5005
R41006 VINP.n394 VINP.n154 4.5005
R41007 VINP.n218 VINP.n154 4.5005
R41008 VINP.n396 VINP.n154 4.5005
R41009 VINP.n217 VINP.n154 4.5005
R41010 VINP.n398 VINP.n154 4.5005
R41011 VINP.n216 VINP.n154 4.5005
R41012 VINP.n400 VINP.n154 4.5005
R41013 VINP.n215 VINP.n154 4.5005
R41014 VINP.n654 VINP.n154 4.5005
R41015 VINP.n656 VINP.n154 4.5005
R41016 VINP.n154 VINP.n0 4.5005
R41017 VINP.n278 VINP.n146 4.5005
R41018 VINP.n276 VINP.n146 4.5005
R41019 VINP.n280 VINP.n146 4.5005
R41020 VINP.n275 VINP.n146 4.5005
R41021 VINP.n282 VINP.n146 4.5005
R41022 VINP.n274 VINP.n146 4.5005
R41023 VINP.n284 VINP.n146 4.5005
R41024 VINP.n273 VINP.n146 4.5005
R41025 VINP.n286 VINP.n146 4.5005
R41026 VINP.n272 VINP.n146 4.5005
R41027 VINP.n288 VINP.n146 4.5005
R41028 VINP.n271 VINP.n146 4.5005
R41029 VINP.n290 VINP.n146 4.5005
R41030 VINP.n270 VINP.n146 4.5005
R41031 VINP.n292 VINP.n146 4.5005
R41032 VINP.n269 VINP.n146 4.5005
R41033 VINP.n294 VINP.n146 4.5005
R41034 VINP.n268 VINP.n146 4.5005
R41035 VINP.n296 VINP.n146 4.5005
R41036 VINP.n267 VINP.n146 4.5005
R41037 VINP.n298 VINP.n146 4.5005
R41038 VINP.n266 VINP.n146 4.5005
R41039 VINP.n300 VINP.n146 4.5005
R41040 VINP.n265 VINP.n146 4.5005
R41041 VINP.n302 VINP.n146 4.5005
R41042 VINP.n264 VINP.n146 4.5005
R41043 VINP.n304 VINP.n146 4.5005
R41044 VINP.n263 VINP.n146 4.5005
R41045 VINP.n306 VINP.n146 4.5005
R41046 VINP.n262 VINP.n146 4.5005
R41047 VINP.n308 VINP.n146 4.5005
R41048 VINP.n261 VINP.n146 4.5005
R41049 VINP.n310 VINP.n146 4.5005
R41050 VINP.n260 VINP.n146 4.5005
R41051 VINP.n312 VINP.n146 4.5005
R41052 VINP.n259 VINP.n146 4.5005
R41053 VINP.n314 VINP.n146 4.5005
R41054 VINP.n258 VINP.n146 4.5005
R41055 VINP.n316 VINP.n146 4.5005
R41056 VINP.n257 VINP.n146 4.5005
R41057 VINP.n318 VINP.n146 4.5005
R41058 VINP.n256 VINP.n146 4.5005
R41059 VINP.n320 VINP.n146 4.5005
R41060 VINP.n255 VINP.n146 4.5005
R41061 VINP.n322 VINP.n146 4.5005
R41062 VINP.n254 VINP.n146 4.5005
R41063 VINP.n324 VINP.n146 4.5005
R41064 VINP.n253 VINP.n146 4.5005
R41065 VINP.n326 VINP.n146 4.5005
R41066 VINP.n252 VINP.n146 4.5005
R41067 VINP.n328 VINP.n146 4.5005
R41068 VINP.n251 VINP.n146 4.5005
R41069 VINP.n330 VINP.n146 4.5005
R41070 VINP.n250 VINP.n146 4.5005
R41071 VINP.n332 VINP.n146 4.5005
R41072 VINP.n249 VINP.n146 4.5005
R41073 VINP.n334 VINP.n146 4.5005
R41074 VINP.n248 VINP.n146 4.5005
R41075 VINP.n336 VINP.n146 4.5005
R41076 VINP.n247 VINP.n146 4.5005
R41077 VINP.n338 VINP.n146 4.5005
R41078 VINP.n246 VINP.n146 4.5005
R41079 VINP.n340 VINP.n146 4.5005
R41080 VINP.n245 VINP.n146 4.5005
R41081 VINP.n342 VINP.n146 4.5005
R41082 VINP.n244 VINP.n146 4.5005
R41083 VINP.n344 VINP.n146 4.5005
R41084 VINP.n243 VINP.n146 4.5005
R41085 VINP.n346 VINP.n146 4.5005
R41086 VINP.n242 VINP.n146 4.5005
R41087 VINP.n348 VINP.n146 4.5005
R41088 VINP.n241 VINP.n146 4.5005
R41089 VINP.n350 VINP.n146 4.5005
R41090 VINP.n240 VINP.n146 4.5005
R41091 VINP.n352 VINP.n146 4.5005
R41092 VINP.n239 VINP.n146 4.5005
R41093 VINP.n354 VINP.n146 4.5005
R41094 VINP.n238 VINP.n146 4.5005
R41095 VINP.n356 VINP.n146 4.5005
R41096 VINP.n237 VINP.n146 4.5005
R41097 VINP.n358 VINP.n146 4.5005
R41098 VINP.n236 VINP.n146 4.5005
R41099 VINP.n360 VINP.n146 4.5005
R41100 VINP.n235 VINP.n146 4.5005
R41101 VINP.n362 VINP.n146 4.5005
R41102 VINP.n234 VINP.n146 4.5005
R41103 VINP.n364 VINP.n146 4.5005
R41104 VINP.n233 VINP.n146 4.5005
R41105 VINP.n366 VINP.n146 4.5005
R41106 VINP.n232 VINP.n146 4.5005
R41107 VINP.n368 VINP.n146 4.5005
R41108 VINP.n231 VINP.n146 4.5005
R41109 VINP.n370 VINP.n146 4.5005
R41110 VINP.n230 VINP.n146 4.5005
R41111 VINP.n372 VINP.n146 4.5005
R41112 VINP.n229 VINP.n146 4.5005
R41113 VINP.n374 VINP.n146 4.5005
R41114 VINP.n228 VINP.n146 4.5005
R41115 VINP.n376 VINP.n146 4.5005
R41116 VINP.n227 VINP.n146 4.5005
R41117 VINP.n378 VINP.n146 4.5005
R41118 VINP.n226 VINP.n146 4.5005
R41119 VINP.n380 VINP.n146 4.5005
R41120 VINP.n225 VINP.n146 4.5005
R41121 VINP.n382 VINP.n146 4.5005
R41122 VINP.n224 VINP.n146 4.5005
R41123 VINP.n384 VINP.n146 4.5005
R41124 VINP.n223 VINP.n146 4.5005
R41125 VINP.n386 VINP.n146 4.5005
R41126 VINP.n222 VINP.n146 4.5005
R41127 VINP.n388 VINP.n146 4.5005
R41128 VINP.n221 VINP.n146 4.5005
R41129 VINP.n390 VINP.n146 4.5005
R41130 VINP.n220 VINP.n146 4.5005
R41131 VINP.n392 VINP.n146 4.5005
R41132 VINP.n219 VINP.n146 4.5005
R41133 VINP.n394 VINP.n146 4.5005
R41134 VINP.n218 VINP.n146 4.5005
R41135 VINP.n396 VINP.n146 4.5005
R41136 VINP.n217 VINP.n146 4.5005
R41137 VINP.n398 VINP.n146 4.5005
R41138 VINP.n216 VINP.n146 4.5005
R41139 VINP.n400 VINP.n146 4.5005
R41140 VINP.n215 VINP.n146 4.5005
R41141 VINP.n654 VINP.n146 4.5005
R41142 VINP.n656 VINP.n146 4.5005
R41143 VINP.n146 VINP.n0 4.5005
R41144 VINP.n278 VINP.n155 4.5005
R41145 VINP.n276 VINP.n155 4.5005
R41146 VINP.n280 VINP.n155 4.5005
R41147 VINP.n275 VINP.n155 4.5005
R41148 VINP.n282 VINP.n155 4.5005
R41149 VINP.n274 VINP.n155 4.5005
R41150 VINP.n284 VINP.n155 4.5005
R41151 VINP.n273 VINP.n155 4.5005
R41152 VINP.n286 VINP.n155 4.5005
R41153 VINP.n272 VINP.n155 4.5005
R41154 VINP.n288 VINP.n155 4.5005
R41155 VINP.n271 VINP.n155 4.5005
R41156 VINP.n290 VINP.n155 4.5005
R41157 VINP.n270 VINP.n155 4.5005
R41158 VINP.n292 VINP.n155 4.5005
R41159 VINP.n269 VINP.n155 4.5005
R41160 VINP.n294 VINP.n155 4.5005
R41161 VINP.n268 VINP.n155 4.5005
R41162 VINP.n296 VINP.n155 4.5005
R41163 VINP.n267 VINP.n155 4.5005
R41164 VINP.n298 VINP.n155 4.5005
R41165 VINP.n266 VINP.n155 4.5005
R41166 VINP.n300 VINP.n155 4.5005
R41167 VINP.n265 VINP.n155 4.5005
R41168 VINP.n302 VINP.n155 4.5005
R41169 VINP.n264 VINP.n155 4.5005
R41170 VINP.n304 VINP.n155 4.5005
R41171 VINP.n263 VINP.n155 4.5005
R41172 VINP.n306 VINP.n155 4.5005
R41173 VINP.n262 VINP.n155 4.5005
R41174 VINP.n308 VINP.n155 4.5005
R41175 VINP.n261 VINP.n155 4.5005
R41176 VINP.n310 VINP.n155 4.5005
R41177 VINP.n260 VINP.n155 4.5005
R41178 VINP.n312 VINP.n155 4.5005
R41179 VINP.n259 VINP.n155 4.5005
R41180 VINP.n314 VINP.n155 4.5005
R41181 VINP.n258 VINP.n155 4.5005
R41182 VINP.n316 VINP.n155 4.5005
R41183 VINP.n257 VINP.n155 4.5005
R41184 VINP.n318 VINP.n155 4.5005
R41185 VINP.n256 VINP.n155 4.5005
R41186 VINP.n320 VINP.n155 4.5005
R41187 VINP.n255 VINP.n155 4.5005
R41188 VINP.n322 VINP.n155 4.5005
R41189 VINP.n254 VINP.n155 4.5005
R41190 VINP.n324 VINP.n155 4.5005
R41191 VINP.n253 VINP.n155 4.5005
R41192 VINP.n326 VINP.n155 4.5005
R41193 VINP.n252 VINP.n155 4.5005
R41194 VINP.n328 VINP.n155 4.5005
R41195 VINP.n251 VINP.n155 4.5005
R41196 VINP.n330 VINP.n155 4.5005
R41197 VINP.n250 VINP.n155 4.5005
R41198 VINP.n332 VINP.n155 4.5005
R41199 VINP.n249 VINP.n155 4.5005
R41200 VINP.n334 VINP.n155 4.5005
R41201 VINP.n248 VINP.n155 4.5005
R41202 VINP.n336 VINP.n155 4.5005
R41203 VINP.n247 VINP.n155 4.5005
R41204 VINP.n338 VINP.n155 4.5005
R41205 VINP.n246 VINP.n155 4.5005
R41206 VINP.n340 VINP.n155 4.5005
R41207 VINP.n245 VINP.n155 4.5005
R41208 VINP.n342 VINP.n155 4.5005
R41209 VINP.n244 VINP.n155 4.5005
R41210 VINP.n344 VINP.n155 4.5005
R41211 VINP.n243 VINP.n155 4.5005
R41212 VINP.n346 VINP.n155 4.5005
R41213 VINP.n242 VINP.n155 4.5005
R41214 VINP.n348 VINP.n155 4.5005
R41215 VINP.n241 VINP.n155 4.5005
R41216 VINP.n350 VINP.n155 4.5005
R41217 VINP.n240 VINP.n155 4.5005
R41218 VINP.n352 VINP.n155 4.5005
R41219 VINP.n239 VINP.n155 4.5005
R41220 VINP.n354 VINP.n155 4.5005
R41221 VINP.n238 VINP.n155 4.5005
R41222 VINP.n356 VINP.n155 4.5005
R41223 VINP.n237 VINP.n155 4.5005
R41224 VINP.n358 VINP.n155 4.5005
R41225 VINP.n236 VINP.n155 4.5005
R41226 VINP.n360 VINP.n155 4.5005
R41227 VINP.n235 VINP.n155 4.5005
R41228 VINP.n362 VINP.n155 4.5005
R41229 VINP.n234 VINP.n155 4.5005
R41230 VINP.n364 VINP.n155 4.5005
R41231 VINP.n233 VINP.n155 4.5005
R41232 VINP.n366 VINP.n155 4.5005
R41233 VINP.n232 VINP.n155 4.5005
R41234 VINP.n368 VINP.n155 4.5005
R41235 VINP.n231 VINP.n155 4.5005
R41236 VINP.n370 VINP.n155 4.5005
R41237 VINP.n230 VINP.n155 4.5005
R41238 VINP.n372 VINP.n155 4.5005
R41239 VINP.n229 VINP.n155 4.5005
R41240 VINP.n374 VINP.n155 4.5005
R41241 VINP.n228 VINP.n155 4.5005
R41242 VINP.n376 VINP.n155 4.5005
R41243 VINP.n227 VINP.n155 4.5005
R41244 VINP.n378 VINP.n155 4.5005
R41245 VINP.n226 VINP.n155 4.5005
R41246 VINP.n380 VINP.n155 4.5005
R41247 VINP.n225 VINP.n155 4.5005
R41248 VINP.n382 VINP.n155 4.5005
R41249 VINP.n224 VINP.n155 4.5005
R41250 VINP.n384 VINP.n155 4.5005
R41251 VINP.n223 VINP.n155 4.5005
R41252 VINP.n386 VINP.n155 4.5005
R41253 VINP.n222 VINP.n155 4.5005
R41254 VINP.n388 VINP.n155 4.5005
R41255 VINP.n221 VINP.n155 4.5005
R41256 VINP.n390 VINP.n155 4.5005
R41257 VINP.n220 VINP.n155 4.5005
R41258 VINP.n392 VINP.n155 4.5005
R41259 VINP.n219 VINP.n155 4.5005
R41260 VINP.n394 VINP.n155 4.5005
R41261 VINP.n218 VINP.n155 4.5005
R41262 VINP.n396 VINP.n155 4.5005
R41263 VINP.n217 VINP.n155 4.5005
R41264 VINP.n398 VINP.n155 4.5005
R41265 VINP.n216 VINP.n155 4.5005
R41266 VINP.n400 VINP.n155 4.5005
R41267 VINP.n215 VINP.n155 4.5005
R41268 VINP.n654 VINP.n155 4.5005
R41269 VINP.n656 VINP.n155 4.5005
R41270 VINP.n155 VINP.n0 4.5005
R41271 VINP.n278 VINP.n145 4.5005
R41272 VINP.n276 VINP.n145 4.5005
R41273 VINP.n280 VINP.n145 4.5005
R41274 VINP.n275 VINP.n145 4.5005
R41275 VINP.n282 VINP.n145 4.5005
R41276 VINP.n274 VINP.n145 4.5005
R41277 VINP.n284 VINP.n145 4.5005
R41278 VINP.n273 VINP.n145 4.5005
R41279 VINP.n286 VINP.n145 4.5005
R41280 VINP.n272 VINP.n145 4.5005
R41281 VINP.n288 VINP.n145 4.5005
R41282 VINP.n271 VINP.n145 4.5005
R41283 VINP.n290 VINP.n145 4.5005
R41284 VINP.n270 VINP.n145 4.5005
R41285 VINP.n292 VINP.n145 4.5005
R41286 VINP.n269 VINP.n145 4.5005
R41287 VINP.n294 VINP.n145 4.5005
R41288 VINP.n268 VINP.n145 4.5005
R41289 VINP.n296 VINP.n145 4.5005
R41290 VINP.n267 VINP.n145 4.5005
R41291 VINP.n298 VINP.n145 4.5005
R41292 VINP.n266 VINP.n145 4.5005
R41293 VINP.n300 VINP.n145 4.5005
R41294 VINP.n265 VINP.n145 4.5005
R41295 VINP.n302 VINP.n145 4.5005
R41296 VINP.n264 VINP.n145 4.5005
R41297 VINP.n304 VINP.n145 4.5005
R41298 VINP.n263 VINP.n145 4.5005
R41299 VINP.n306 VINP.n145 4.5005
R41300 VINP.n262 VINP.n145 4.5005
R41301 VINP.n308 VINP.n145 4.5005
R41302 VINP.n261 VINP.n145 4.5005
R41303 VINP.n310 VINP.n145 4.5005
R41304 VINP.n260 VINP.n145 4.5005
R41305 VINP.n312 VINP.n145 4.5005
R41306 VINP.n259 VINP.n145 4.5005
R41307 VINP.n314 VINP.n145 4.5005
R41308 VINP.n258 VINP.n145 4.5005
R41309 VINP.n316 VINP.n145 4.5005
R41310 VINP.n257 VINP.n145 4.5005
R41311 VINP.n318 VINP.n145 4.5005
R41312 VINP.n256 VINP.n145 4.5005
R41313 VINP.n320 VINP.n145 4.5005
R41314 VINP.n255 VINP.n145 4.5005
R41315 VINP.n322 VINP.n145 4.5005
R41316 VINP.n254 VINP.n145 4.5005
R41317 VINP.n324 VINP.n145 4.5005
R41318 VINP.n253 VINP.n145 4.5005
R41319 VINP.n326 VINP.n145 4.5005
R41320 VINP.n252 VINP.n145 4.5005
R41321 VINP.n328 VINP.n145 4.5005
R41322 VINP.n251 VINP.n145 4.5005
R41323 VINP.n330 VINP.n145 4.5005
R41324 VINP.n250 VINP.n145 4.5005
R41325 VINP.n332 VINP.n145 4.5005
R41326 VINP.n249 VINP.n145 4.5005
R41327 VINP.n334 VINP.n145 4.5005
R41328 VINP.n248 VINP.n145 4.5005
R41329 VINP.n336 VINP.n145 4.5005
R41330 VINP.n247 VINP.n145 4.5005
R41331 VINP.n338 VINP.n145 4.5005
R41332 VINP.n246 VINP.n145 4.5005
R41333 VINP.n340 VINP.n145 4.5005
R41334 VINP.n245 VINP.n145 4.5005
R41335 VINP.n342 VINP.n145 4.5005
R41336 VINP.n244 VINP.n145 4.5005
R41337 VINP.n344 VINP.n145 4.5005
R41338 VINP.n243 VINP.n145 4.5005
R41339 VINP.n346 VINP.n145 4.5005
R41340 VINP.n242 VINP.n145 4.5005
R41341 VINP.n348 VINP.n145 4.5005
R41342 VINP.n241 VINP.n145 4.5005
R41343 VINP.n350 VINP.n145 4.5005
R41344 VINP.n240 VINP.n145 4.5005
R41345 VINP.n352 VINP.n145 4.5005
R41346 VINP.n239 VINP.n145 4.5005
R41347 VINP.n354 VINP.n145 4.5005
R41348 VINP.n238 VINP.n145 4.5005
R41349 VINP.n356 VINP.n145 4.5005
R41350 VINP.n237 VINP.n145 4.5005
R41351 VINP.n358 VINP.n145 4.5005
R41352 VINP.n236 VINP.n145 4.5005
R41353 VINP.n360 VINP.n145 4.5005
R41354 VINP.n235 VINP.n145 4.5005
R41355 VINP.n362 VINP.n145 4.5005
R41356 VINP.n234 VINP.n145 4.5005
R41357 VINP.n364 VINP.n145 4.5005
R41358 VINP.n233 VINP.n145 4.5005
R41359 VINP.n366 VINP.n145 4.5005
R41360 VINP.n232 VINP.n145 4.5005
R41361 VINP.n368 VINP.n145 4.5005
R41362 VINP.n231 VINP.n145 4.5005
R41363 VINP.n370 VINP.n145 4.5005
R41364 VINP.n230 VINP.n145 4.5005
R41365 VINP.n372 VINP.n145 4.5005
R41366 VINP.n229 VINP.n145 4.5005
R41367 VINP.n374 VINP.n145 4.5005
R41368 VINP.n228 VINP.n145 4.5005
R41369 VINP.n376 VINP.n145 4.5005
R41370 VINP.n227 VINP.n145 4.5005
R41371 VINP.n378 VINP.n145 4.5005
R41372 VINP.n226 VINP.n145 4.5005
R41373 VINP.n380 VINP.n145 4.5005
R41374 VINP.n225 VINP.n145 4.5005
R41375 VINP.n382 VINP.n145 4.5005
R41376 VINP.n224 VINP.n145 4.5005
R41377 VINP.n384 VINP.n145 4.5005
R41378 VINP.n223 VINP.n145 4.5005
R41379 VINP.n386 VINP.n145 4.5005
R41380 VINP.n222 VINP.n145 4.5005
R41381 VINP.n388 VINP.n145 4.5005
R41382 VINP.n221 VINP.n145 4.5005
R41383 VINP.n390 VINP.n145 4.5005
R41384 VINP.n220 VINP.n145 4.5005
R41385 VINP.n392 VINP.n145 4.5005
R41386 VINP.n219 VINP.n145 4.5005
R41387 VINP.n394 VINP.n145 4.5005
R41388 VINP.n218 VINP.n145 4.5005
R41389 VINP.n396 VINP.n145 4.5005
R41390 VINP.n217 VINP.n145 4.5005
R41391 VINP.n398 VINP.n145 4.5005
R41392 VINP.n216 VINP.n145 4.5005
R41393 VINP.n400 VINP.n145 4.5005
R41394 VINP.n215 VINP.n145 4.5005
R41395 VINP.n654 VINP.n145 4.5005
R41396 VINP.n656 VINP.n145 4.5005
R41397 VINP.n145 VINP.n0 4.5005
R41398 VINP.n278 VINP.n156 4.5005
R41399 VINP.n276 VINP.n156 4.5005
R41400 VINP.n280 VINP.n156 4.5005
R41401 VINP.n275 VINP.n156 4.5005
R41402 VINP.n282 VINP.n156 4.5005
R41403 VINP.n274 VINP.n156 4.5005
R41404 VINP.n284 VINP.n156 4.5005
R41405 VINP.n273 VINP.n156 4.5005
R41406 VINP.n286 VINP.n156 4.5005
R41407 VINP.n272 VINP.n156 4.5005
R41408 VINP.n288 VINP.n156 4.5005
R41409 VINP.n271 VINP.n156 4.5005
R41410 VINP.n290 VINP.n156 4.5005
R41411 VINP.n270 VINP.n156 4.5005
R41412 VINP.n292 VINP.n156 4.5005
R41413 VINP.n269 VINP.n156 4.5005
R41414 VINP.n294 VINP.n156 4.5005
R41415 VINP.n268 VINP.n156 4.5005
R41416 VINP.n296 VINP.n156 4.5005
R41417 VINP.n267 VINP.n156 4.5005
R41418 VINP.n298 VINP.n156 4.5005
R41419 VINP.n266 VINP.n156 4.5005
R41420 VINP.n300 VINP.n156 4.5005
R41421 VINP.n265 VINP.n156 4.5005
R41422 VINP.n302 VINP.n156 4.5005
R41423 VINP.n264 VINP.n156 4.5005
R41424 VINP.n304 VINP.n156 4.5005
R41425 VINP.n263 VINP.n156 4.5005
R41426 VINP.n306 VINP.n156 4.5005
R41427 VINP.n262 VINP.n156 4.5005
R41428 VINP.n308 VINP.n156 4.5005
R41429 VINP.n261 VINP.n156 4.5005
R41430 VINP.n310 VINP.n156 4.5005
R41431 VINP.n260 VINP.n156 4.5005
R41432 VINP.n312 VINP.n156 4.5005
R41433 VINP.n259 VINP.n156 4.5005
R41434 VINP.n314 VINP.n156 4.5005
R41435 VINP.n258 VINP.n156 4.5005
R41436 VINP.n316 VINP.n156 4.5005
R41437 VINP.n257 VINP.n156 4.5005
R41438 VINP.n318 VINP.n156 4.5005
R41439 VINP.n256 VINP.n156 4.5005
R41440 VINP.n320 VINP.n156 4.5005
R41441 VINP.n255 VINP.n156 4.5005
R41442 VINP.n322 VINP.n156 4.5005
R41443 VINP.n254 VINP.n156 4.5005
R41444 VINP.n324 VINP.n156 4.5005
R41445 VINP.n253 VINP.n156 4.5005
R41446 VINP.n326 VINP.n156 4.5005
R41447 VINP.n252 VINP.n156 4.5005
R41448 VINP.n328 VINP.n156 4.5005
R41449 VINP.n251 VINP.n156 4.5005
R41450 VINP.n330 VINP.n156 4.5005
R41451 VINP.n250 VINP.n156 4.5005
R41452 VINP.n332 VINP.n156 4.5005
R41453 VINP.n249 VINP.n156 4.5005
R41454 VINP.n334 VINP.n156 4.5005
R41455 VINP.n248 VINP.n156 4.5005
R41456 VINP.n336 VINP.n156 4.5005
R41457 VINP.n247 VINP.n156 4.5005
R41458 VINP.n338 VINP.n156 4.5005
R41459 VINP.n246 VINP.n156 4.5005
R41460 VINP.n340 VINP.n156 4.5005
R41461 VINP.n245 VINP.n156 4.5005
R41462 VINP.n342 VINP.n156 4.5005
R41463 VINP.n244 VINP.n156 4.5005
R41464 VINP.n344 VINP.n156 4.5005
R41465 VINP.n243 VINP.n156 4.5005
R41466 VINP.n346 VINP.n156 4.5005
R41467 VINP.n242 VINP.n156 4.5005
R41468 VINP.n348 VINP.n156 4.5005
R41469 VINP.n241 VINP.n156 4.5005
R41470 VINP.n350 VINP.n156 4.5005
R41471 VINP.n240 VINP.n156 4.5005
R41472 VINP.n352 VINP.n156 4.5005
R41473 VINP.n239 VINP.n156 4.5005
R41474 VINP.n354 VINP.n156 4.5005
R41475 VINP.n238 VINP.n156 4.5005
R41476 VINP.n356 VINP.n156 4.5005
R41477 VINP.n237 VINP.n156 4.5005
R41478 VINP.n358 VINP.n156 4.5005
R41479 VINP.n236 VINP.n156 4.5005
R41480 VINP.n360 VINP.n156 4.5005
R41481 VINP.n235 VINP.n156 4.5005
R41482 VINP.n362 VINP.n156 4.5005
R41483 VINP.n234 VINP.n156 4.5005
R41484 VINP.n364 VINP.n156 4.5005
R41485 VINP.n233 VINP.n156 4.5005
R41486 VINP.n366 VINP.n156 4.5005
R41487 VINP.n232 VINP.n156 4.5005
R41488 VINP.n368 VINP.n156 4.5005
R41489 VINP.n231 VINP.n156 4.5005
R41490 VINP.n370 VINP.n156 4.5005
R41491 VINP.n230 VINP.n156 4.5005
R41492 VINP.n372 VINP.n156 4.5005
R41493 VINP.n229 VINP.n156 4.5005
R41494 VINP.n374 VINP.n156 4.5005
R41495 VINP.n228 VINP.n156 4.5005
R41496 VINP.n376 VINP.n156 4.5005
R41497 VINP.n227 VINP.n156 4.5005
R41498 VINP.n378 VINP.n156 4.5005
R41499 VINP.n226 VINP.n156 4.5005
R41500 VINP.n380 VINP.n156 4.5005
R41501 VINP.n225 VINP.n156 4.5005
R41502 VINP.n382 VINP.n156 4.5005
R41503 VINP.n224 VINP.n156 4.5005
R41504 VINP.n384 VINP.n156 4.5005
R41505 VINP.n223 VINP.n156 4.5005
R41506 VINP.n386 VINP.n156 4.5005
R41507 VINP.n222 VINP.n156 4.5005
R41508 VINP.n388 VINP.n156 4.5005
R41509 VINP.n221 VINP.n156 4.5005
R41510 VINP.n390 VINP.n156 4.5005
R41511 VINP.n220 VINP.n156 4.5005
R41512 VINP.n392 VINP.n156 4.5005
R41513 VINP.n219 VINP.n156 4.5005
R41514 VINP.n394 VINP.n156 4.5005
R41515 VINP.n218 VINP.n156 4.5005
R41516 VINP.n396 VINP.n156 4.5005
R41517 VINP.n217 VINP.n156 4.5005
R41518 VINP.n398 VINP.n156 4.5005
R41519 VINP.n216 VINP.n156 4.5005
R41520 VINP.n400 VINP.n156 4.5005
R41521 VINP.n215 VINP.n156 4.5005
R41522 VINP.n654 VINP.n156 4.5005
R41523 VINP.n656 VINP.n156 4.5005
R41524 VINP.n156 VINP.n0 4.5005
R41525 VINP.n278 VINP.n144 4.5005
R41526 VINP.n276 VINP.n144 4.5005
R41527 VINP.n280 VINP.n144 4.5005
R41528 VINP.n275 VINP.n144 4.5005
R41529 VINP.n282 VINP.n144 4.5005
R41530 VINP.n274 VINP.n144 4.5005
R41531 VINP.n284 VINP.n144 4.5005
R41532 VINP.n273 VINP.n144 4.5005
R41533 VINP.n286 VINP.n144 4.5005
R41534 VINP.n272 VINP.n144 4.5005
R41535 VINP.n288 VINP.n144 4.5005
R41536 VINP.n271 VINP.n144 4.5005
R41537 VINP.n290 VINP.n144 4.5005
R41538 VINP.n270 VINP.n144 4.5005
R41539 VINP.n292 VINP.n144 4.5005
R41540 VINP.n269 VINP.n144 4.5005
R41541 VINP.n294 VINP.n144 4.5005
R41542 VINP.n268 VINP.n144 4.5005
R41543 VINP.n296 VINP.n144 4.5005
R41544 VINP.n267 VINP.n144 4.5005
R41545 VINP.n298 VINP.n144 4.5005
R41546 VINP.n266 VINP.n144 4.5005
R41547 VINP.n300 VINP.n144 4.5005
R41548 VINP.n265 VINP.n144 4.5005
R41549 VINP.n302 VINP.n144 4.5005
R41550 VINP.n264 VINP.n144 4.5005
R41551 VINP.n304 VINP.n144 4.5005
R41552 VINP.n263 VINP.n144 4.5005
R41553 VINP.n306 VINP.n144 4.5005
R41554 VINP.n262 VINP.n144 4.5005
R41555 VINP.n308 VINP.n144 4.5005
R41556 VINP.n261 VINP.n144 4.5005
R41557 VINP.n310 VINP.n144 4.5005
R41558 VINP.n260 VINP.n144 4.5005
R41559 VINP.n312 VINP.n144 4.5005
R41560 VINP.n259 VINP.n144 4.5005
R41561 VINP.n314 VINP.n144 4.5005
R41562 VINP.n258 VINP.n144 4.5005
R41563 VINP.n316 VINP.n144 4.5005
R41564 VINP.n257 VINP.n144 4.5005
R41565 VINP.n318 VINP.n144 4.5005
R41566 VINP.n256 VINP.n144 4.5005
R41567 VINP.n320 VINP.n144 4.5005
R41568 VINP.n255 VINP.n144 4.5005
R41569 VINP.n322 VINP.n144 4.5005
R41570 VINP.n254 VINP.n144 4.5005
R41571 VINP.n324 VINP.n144 4.5005
R41572 VINP.n253 VINP.n144 4.5005
R41573 VINP.n326 VINP.n144 4.5005
R41574 VINP.n252 VINP.n144 4.5005
R41575 VINP.n328 VINP.n144 4.5005
R41576 VINP.n251 VINP.n144 4.5005
R41577 VINP.n330 VINP.n144 4.5005
R41578 VINP.n250 VINP.n144 4.5005
R41579 VINP.n332 VINP.n144 4.5005
R41580 VINP.n249 VINP.n144 4.5005
R41581 VINP.n334 VINP.n144 4.5005
R41582 VINP.n248 VINP.n144 4.5005
R41583 VINP.n336 VINP.n144 4.5005
R41584 VINP.n247 VINP.n144 4.5005
R41585 VINP.n338 VINP.n144 4.5005
R41586 VINP.n246 VINP.n144 4.5005
R41587 VINP.n340 VINP.n144 4.5005
R41588 VINP.n245 VINP.n144 4.5005
R41589 VINP.n342 VINP.n144 4.5005
R41590 VINP.n244 VINP.n144 4.5005
R41591 VINP.n344 VINP.n144 4.5005
R41592 VINP.n243 VINP.n144 4.5005
R41593 VINP.n346 VINP.n144 4.5005
R41594 VINP.n242 VINP.n144 4.5005
R41595 VINP.n348 VINP.n144 4.5005
R41596 VINP.n241 VINP.n144 4.5005
R41597 VINP.n350 VINP.n144 4.5005
R41598 VINP.n240 VINP.n144 4.5005
R41599 VINP.n352 VINP.n144 4.5005
R41600 VINP.n239 VINP.n144 4.5005
R41601 VINP.n354 VINP.n144 4.5005
R41602 VINP.n238 VINP.n144 4.5005
R41603 VINP.n356 VINP.n144 4.5005
R41604 VINP.n237 VINP.n144 4.5005
R41605 VINP.n358 VINP.n144 4.5005
R41606 VINP.n236 VINP.n144 4.5005
R41607 VINP.n360 VINP.n144 4.5005
R41608 VINP.n235 VINP.n144 4.5005
R41609 VINP.n362 VINP.n144 4.5005
R41610 VINP.n234 VINP.n144 4.5005
R41611 VINP.n364 VINP.n144 4.5005
R41612 VINP.n233 VINP.n144 4.5005
R41613 VINP.n366 VINP.n144 4.5005
R41614 VINP.n232 VINP.n144 4.5005
R41615 VINP.n368 VINP.n144 4.5005
R41616 VINP.n231 VINP.n144 4.5005
R41617 VINP.n370 VINP.n144 4.5005
R41618 VINP.n230 VINP.n144 4.5005
R41619 VINP.n372 VINP.n144 4.5005
R41620 VINP.n229 VINP.n144 4.5005
R41621 VINP.n374 VINP.n144 4.5005
R41622 VINP.n228 VINP.n144 4.5005
R41623 VINP.n376 VINP.n144 4.5005
R41624 VINP.n227 VINP.n144 4.5005
R41625 VINP.n378 VINP.n144 4.5005
R41626 VINP.n226 VINP.n144 4.5005
R41627 VINP.n380 VINP.n144 4.5005
R41628 VINP.n225 VINP.n144 4.5005
R41629 VINP.n382 VINP.n144 4.5005
R41630 VINP.n224 VINP.n144 4.5005
R41631 VINP.n384 VINP.n144 4.5005
R41632 VINP.n223 VINP.n144 4.5005
R41633 VINP.n386 VINP.n144 4.5005
R41634 VINP.n222 VINP.n144 4.5005
R41635 VINP.n388 VINP.n144 4.5005
R41636 VINP.n221 VINP.n144 4.5005
R41637 VINP.n390 VINP.n144 4.5005
R41638 VINP.n220 VINP.n144 4.5005
R41639 VINP.n392 VINP.n144 4.5005
R41640 VINP.n219 VINP.n144 4.5005
R41641 VINP.n394 VINP.n144 4.5005
R41642 VINP.n218 VINP.n144 4.5005
R41643 VINP.n396 VINP.n144 4.5005
R41644 VINP.n217 VINP.n144 4.5005
R41645 VINP.n398 VINP.n144 4.5005
R41646 VINP.n216 VINP.n144 4.5005
R41647 VINP.n400 VINP.n144 4.5005
R41648 VINP.n215 VINP.n144 4.5005
R41649 VINP.n654 VINP.n144 4.5005
R41650 VINP.n656 VINP.n144 4.5005
R41651 VINP.n144 VINP.n0 4.5005
R41652 VINP.n278 VINP.n157 4.5005
R41653 VINP.n276 VINP.n157 4.5005
R41654 VINP.n280 VINP.n157 4.5005
R41655 VINP.n275 VINP.n157 4.5005
R41656 VINP.n282 VINP.n157 4.5005
R41657 VINP.n274 VINP.n157 4.5005
R41658 VINP.n284 VINP.n157 4.5005
R41659 VINP.n273 VINP.n157 4.5005
R41660 VINP.n286 VINP.n157 4.5005
R41661 VINP.n272 VINP.n157 4.5005
R41662 VINP.n288 VINP.n157 4.5005
R41663 VINP.n271 VINP.n157 4.5005
R41664 VINP.n290 VINP.n157 4.5005
R41665 VINP.n270 VINP.n157 4.5005
R41666 VINP.n292 VINP.n157 4.5005
R41667 VINP.n269 VINP.n157 4.5005
R41668 VINP.n294 VINP.n157 4.5005
R41669 VINP.n268 VINP.n157 4.5005
R41670 VINP.n296 VINP.n157 4.5005
R41671 VINP.n267 VINP.n157 4.5005
R41672 VINP.n298 VINP.n157 4.5005
R41673 VINP.n266 VINP.n157 4.5005
R41674 VINP.n300 VINP.n157 4.5005
R41675 VINP.n265 VINP.n157 4.5005
R41676 VINP.n302 VINP.n157 4.5005
R41677 VINP.n264 VINP.n157 4.5005
R41678 VINP.n304 VINP.n157 4.5005
R41679 VINP.n263 VINP.n157 4.5005
R41680 VINP.n306 VINP.n157 4.5005
R41681 VINP.n262 VINP.n157 4.5005
R41682 VINP.n308 VINP.n157 4.5005
R41683 VINP.n261 VINP.n157 4.5005
R41684 VINP.n310 VINP.n157 4.5005
R41685 VINP.n260 VINP.n157 4.5005
R41686 VINP.n312 VINP.n157 4.5005
R41687 VINP.n259 VINP.n157 4.5005
R41688 VINP.n314 VINP.n157 4.5005
R41689 VINP.n258 VINP.n157 4.5005
R41690 VINP.n316 VINP.n157 4.5005
R41691 VINP.n257 VINP.n157 4.5005
R41692 VINP.n318 VINP.n157 4.5005
R41693 VINP.n256 VINP.n157 4.5005
R41694 VINP.n320 VINP.n157 4.5005
R41695 VINP.n255 VINP.n157 4.5005
R41696 VINP.n322 VINP.n157 4.5005
R41697 VINP.n254 VINP.n157 4.5005
R41698 VINP.n324 VINP.n157 4.5005
R41699 VINP.n253 VINP.n157 4.5005
R41700 VINP.n326 VINP.n157 4.5005
R41701 VINP.n252 VINP.n157 4.5005
R41702 VINP.n328 VINP.n157 4.5005
R41703 VINP.n251 VINP.n157 4.5005
R41704 VINP.n330 VINP.n157 4.5005
R41705 VINP.n250 VINP.n157 4.5005
R41706 VINP.n332 VINP.n157 4.5005
R41707 VINP.n249 VINP.n157 4.5005
R41708 VINP.n334 VINP.n157 4.5005
R41709 VINP.n248 VINP.n157 4.5005
R41710 VINP.n336 VINP.n157 4.5005
R41711 VINP.n247 VINP.n157 4.5005
R41712 VINP.n338 VINP.n157 4.5005
R41713 VINP.n246 VINP.n157 4.5005
R41714 VINP.n340 VINP.n157 4.5005
R41715 VINP.n245 VINP.n157 4.5005
R41716 VINP.n342 VINP.n157 4.5005
R41717 VINP.n244 VINP.n157 4.5005
R41718 VINP.n344 VINP.n157 4.5005
R41719 VINP.n243 VINP.n157 4.5005
R41720 VINP.n346 VINP.n157 4.5005
R41721 VINP.n242 VINP.n157 4.5005
R41722 VINP.n348 VINP.n157 4.5005
R41723 VINP.n241 VINP.n157 4.5005
R41724 VINP.n350 VINP.n157 4.5005
R41725 VINP.n240 VINP.n157 4.5005
R41726 VINP.n352 VINP.n157 4.5005
R41727 VINP.n239 VINP.n157 4.5005
R41728 VINP.n354 VINP.n157 4.5005
R41729 VINP.n238 VINP.n157 4.5005
R41730 VINP.n356 VINP.n157 4.5005
R41731 VINP.n237 VINP.n157 4.5005
R41732 VINP.n358 VINP.n157 4.5005
R41733 VINP.n236 VINP.n157 4.5005
R41734 VINP.n360 VINP.n157 4.5005
R41735 VINP.n235 VINP.n157 4.5005
R41736 VINP.n362 VINP.n157 4.5005
R41737 VINP.n234 VINP.n157 4.5005
R41738 VINP.n364 VINP.n157 4.5005
R41739 VINP.n233 VINP.n157 4.5005
R41740 VINP.n366 VINP.n157 4.5005
R41741 VINP.n232 VINP.n157 4.5005
R41742 VINP.n368 VINP.n157 4.5005
R41743 VINP.n231 VINP.n157 4.5005
R41744 VINP.n370 VINP.n157 4.5005
R41745 VINP.n230 VINP.n157 4.5005
R41746 VINP.n372 VINP.n157 4.5005
R41747 VINP.n229 VINP.n157 4.5005
R41748 VINP.n374 VINP.n157 4.5005
R41749 VINP.n228 VINP.n157 4.5005
R41750 VINP.n376 VINP.n157 4.5005
R41751 VINP.n227 VINP.n157 4.5005
R41752 VINP.n378 VINP.n157 4.5005
R41753 VINP.n226 VINP.n157 4.5005
R41754 VINP.n380 VINP.n157 4.5005
R41755 VINP.n225 VINP.n157 4.5005
R41756 VINP.n382 VINP.n157 4.5005
R41757 VINP.n224 VINP.n157 4.5005
R41758 VINP.n384 VINP.n157 4.5005
R41759 VINP.n223 VINP.n157 4.5005
R41760 VINP.n386 VINP.n157 4.5005
R41761 VINP.n222 VINP.n157 4.5005
R41762 VINP.n388 VINP.n157 4.5005
R41763 VINP.n221 VINP.n157 4.5005
R41764 VINP.n390 VINP.n157 4.5005
R41765 VINP.n220 VINP.n157 4.5005
R41766 VINP.n392 VINP.n157 4.5005
R41767 VINP.n219 VINP.n157 4.5005
R41768 VINP.n394 VINP.n157 4.5005
R41769 VINP.n218 VINP.n157 4.5005
R41770 VINP.n396 VINP.n157 4.5005
R41771 VINP.n217 VINP.n157 4.5005
R41772 VINP.n398 VINP.n157 4.5005
R41773 VINP.n216 VINP.n157 4.5005
R41774 VINP.n400 VINP.n157 4.5005
R41775 VINP.n215 VINP.n157 4.5005
R41776 VINP.n654 VINP.n157 4.5005
R41777 VINP.n656 VINP.n157 4.5005
R41778 VINP.n157 VINP.n0 4.5005
R41779 VINP.n278 VINP.n143 4.5005
R41780 VINP.n276 VINP.n143 4.5005
R41781 VINP.n280 VINP.n143 4.5005
R41782 VINP.n275 VINP.n143 4.5005
R41783 VINP.n282 VINP.n143 4.5005
R41784 VINP.n274 VINP.n143 4.5005
R41785 VINP.n284 VINP.n143 4.5005
R41786 VINP.n273 VINP.n143 4.5005
R41787 VINP.n286 VINP.n143 4.5005
R41788 VINP.n272 VINP.n143 4.5005
R41789 VINP.n288 VINP.n143 4.5005
R41790 VINP.n271 VINP.n143 4.5005
R41791 VINP.n290 VINP.n143 4.5005
R41792 VINP.n270 VINP.n143 4.5005
R41793 VINP.n292 VINP.n143 4.5005
R41794 VINP.n269 VINP.n143 4.5005
R41795 VINP.n294 VINP.n143 4.5005
R41796 VINP.n268 VINP.n143 4.5005
R41797 VINP.n296 VINP.n143 4.5005
R41798 VINP.n267 VINP.n143 4.5005
R41799 VINP.n298 VINP.n143 4.5005
R41800 VINP.n266 VINP.n143 4.5005
R41801 VINP.n300 VINP.n143 4.5005
R41802 VINP.n265 VINP.n143 4.5005
R41803 VINP.n302 VINP.n143 4.5005
R41804 VINP.n264 VINP.n143 4.5005
R41805 VINP.n304 VINP.n143 4.5005
R41806 VINP.n263 VINP.n143 4.5005
R41807 VINP.n306 VINP.n143 4.5005
R41808 VINP.n262 VINP.n143 4.5005
R41809 VINP.n308 VINP.n143 4.5005
R41810 VINP.n261 VINP.n143 4.5005
R41811 VINP.n310 VINP.n143 4.5005
R41812 VINP.n260 VINP.n143 4.5005
R41813 VINP.n312 VINP.n143 4.5005
R41814 VINP.n259 VINP.n143 4.5005
R41815 VINP.n314 VINP.n143 4.5005
R41816 VINP.n258 VINP.n143 4.5005
R41817 VINP.n316 VINP.n143 4.5005
R41818 VINP.n257 VINP.n143 4.5005
R41819 VINP.n318 VINP.n143 4.5005
R41820 VINP.n256 VINP.n143 4.5005
R41821 VINP.n320 VINP.n143 4.5005
R41822 VINP.n255 VINP.n143 4.5005
R41823 VINP.n322 VINP.n143 4.5005
R41824 VINP.n254 VINP.n143 4.5005
R41825 VINP.n324 VINP.n143 4.5005
R41826 VINP.n253 VINP.n143 4.5005
R41827 VINP.n326 VINP.n143 4.5005
R41828 VINP.n252 VINP.n143 4.5005
R41829 VINP.n328 VINP.n143 4.5005
R41830 VINP.n251 VINP.n143 4.5005
R41831 VINP.n330 VINP.n143 4.5005
R41832 VINP.n250 VINP.n143 4.5005
R41833 VINP.n332 VINP.n143 4.5005
R41834 VINP.n249 VINP.n143 4.5005
R41835 VINP.n334 VINP.n143 4.5005
R41836 VINP.n248 VINP.n143 4.5005
R41837 VINP.n336 VINP.n143 4.5005
R41838 VINP.n247 VINP.n143 4.5005
R41839 VINP.n338 VINP.n143 4.5005
R41840 VINP.n246 VINP.n143 4.5005
R41841 VINP.n340 VINP.n143 4.5005
R41842 VINP.n245 VINP.n143 4.5005
R41843 VINP.n342 VINP.n143 4.5005
R41844 VINP.n244 VINP.n143 4.5005
R41845 VINP.n344 VINP.n143 4.5005
R41846 VINP.n243 VINP.n143 4.5005
R41847 VINP.n346 VINP.n143 4.5005
R41848 VINP.n242 VINP.n143 4.5005
R41849 VINP.n348 VINP.n143 4.5005
R41850 VINP.n241 VINP.n143 4.5005
R41851 VINP.n350 VINP.n143 4.5005
R41852 VINP.n240 VINP.n143 4.5005
R41853 VINP.n352 VINP.n143 4.5005
R41854 VINP.n239 VINP.n143 4.5005
R41855 VINP.n354 VINP.n143 4.5005
R41856 VINP.n238 VINP.n143 4.5005
R41857 VINP.n356 VINP.n143 4.5005
R41858 VINP.n237 VINP.n143 4.5005
R41859 VINP.n358 VINP.n143 4.5005
R41860 VINP.n236 VINP.n143 4.5005
R41861 VINP.n360 VINP.n143 4.5005
R41862 VINP.n235 VINP.n143 4.5005
R41863 VINP.n362 VINP.n143 4.5005
R41864 VINP.n234 VINP.n143 4.5005
R41865 VINP.n364 VINP.n143 4.5005
R41866 VINP.n233 VINP.n143 4.5005
R41867 VINP.n366 VINP.n143 4.5005
R41868 VINP.n232 VINP.n143 4.5005
R41869 VINP.n368 VINP.n143 4.5005
R41870 VINP.n231 VINP.n143 4.5005
R41871 VINP.n370 VINP.n143 4.5005
R41872 VINP.n230 VINP.n143 4.5005
R41873 VINP.n372 VINP.n143 4.5005
R41874 VINP.n229 VINP.n143 4.5005
R41875 VINP.n374 VINP.n143 4.5005
R41876 VINP.n228 VINP.n143 4.5005
R41877 VINP.n376 VINP.n143 4.5005
R41878 VINP.n227 VINP.n143 4.5005
R41879 VINP.n378 VINP.n143 4.5005
R41880 VINP.n226 VINP.n143 4.5005
R41881 VINP.n380 VINP.n143 4.5005
R41882 VINP.n225 VINP.n143 4.5005
R41883 VINP.n382 VINP.n143 4.5005
R41884 VINP.n224 VINP.n143 4.5005
R41885 VINP.n384 VINP.n143 4.5005
R41886 VINP.n223 VINP.n143 4.5005
R41887 VINP.n386 VINP.n143 4.5005
R41888 VINP.n222 VINP.n143 4.5005
R41889 VINP.n388 VINP.n143 4.5005
R41890 VINP.n221 VINP.n143 4.5005
R41891 VINP.n390 VINP.n143 4.5005
R41892 VINP.n220 VINP.n143 4.5005
R41893 VINP.n392 VINP.n143 4.5005
R41894 VINP.n219 VINP.n143 4.5005
R41895 VINP.n394 VINP.n143 4.5005
R41896 VINP.n218 VINP.n143 4.5005
R41897 VINP.n396 VINP.n143 4.5005
R41898 VINP.n217 VINP.n143 4.5005
R41899 VINP.n398 VINP.n143 4.5005
R41900 VINP.n216 VINP.n143 4.5005
R41901 VINP.n400 VINP.n143 4.5005
R41902 VINP.n215 VINP.n143 4.5005
R41903 VINP.n654 VINP.n143 4.5005
R41904 VINP.n656 VINP.n143 4.5005
R41905 VINP.n143 VINP.n0 4.5005
R41906 VINP.n278 VINP.n158 4.5005
R41907 VINP.n276 VINP.n158 4.5005
R41908 VINP.n280 VINP.n158 4.5005
R41909 VINP.n275 VINP.n158 4.5005
R41910 VINP.n282 VINP.n158 4.5005
R41911 VINP.n274 VINP.n158 4.5005
R41912 VINP.n284 VINP.n158 4.5005
R41913 VINP.n273 VINP.n158 4.5005
R41914 VINP.n286 VINP.n158 4.5005
R41915 VINP.n272 VINP.n158 4.5005
R41916 VINP.n288 VINP.n158 4.5005
R41917 VINP.n271 VINP.n158 4.5005
R41918 VINP.n290 VINP.n158 4.5005
R41919 VINP.n270 VINP.n158 4.5005
R41920 VINP.n292 VINP.n158 4.5005
R41921 VINP.n269 VINP.n158 4.5005
R41922 VINP.n294 VINP.n158 4.5005
R41923 VINP.n268 VINP.n158 4.5005
R41924 VINP.n296 VINP.n158 4.5005
R41925 VINP.n267 VINP.n158 4.5005
R41926 VINP.n298 VINP.n158 4.5005
R41927 VINP.n266 VINP.n158 4.5005
R41928 VINP.n300 VINP.n158 4.5005
R41929 VINP.n265 VINP.n158 4.5005
R41930 VINP.n302 VINP.n158 4.5005
R41931 VINP.n264 VINP.n158 4.5005
R41932 VINP.n304 VINP.n158 4.5005
R41933 VINP.n263 VINP.n158 4.5005
R41934 VINP.n306 VINP.n158 4.5005
R41935 VINP.n262 VINP.n158 4.5005
R41936 VINP.n308 VINP.n158 4.5005
R41937 VINP.n261 VINP.n158 4.5005
R41938 VINP.n310 VINP.n158 4.5005
R41939 VINP.n260 VINP.n158 4.5005
R41940 VINP.n312 VINP.n158 4.5005
R41941 VINP.n259 VINP.n158 4.5005
R41942 VINP.n314 VINP.n158 4.5005
R41943 VINP.n258 VINP.n158 4.5005
R41944 VINP.n316 VINP.n158 4.5005
R41945 VINP.n257 VINP.n158 4.5005
R41946 VINP.n318 VINP.n158 4.5005
R41947 VINP.n256 VINP.n158 4.5005
R41948 VINP.n320 VINP.n158 4.5005
R41949 VINP.n255 VINP.n158 4.5005
R41950 VINP.n322 VINP.n158 4.5005
R41951 VINP.n254 VINP.n158 4.5005
R41952 VINP.n324 VINP.n158 4.5005
R41953 VINP.n253 VINP.n158 4.5005
R41954 VINP.n326 VINP.n158 4.5005
R41955 VINP.n252 VINP.n158 4.5005
R41956 VINP.n328 VINP.n158 4.5005
R41957 VINP.n251 VINP.n158 4.5005
R41958 VINP.n330 VINP.n158 4.5005
R41959 VINP.n250 VINP.n158 4.5005
R41960 VINP.n332 VINP.n158 4.5005
R41961 VINP.n249 VINP.n158 4.5005
R41962 VINP.n334 VINP.n158 4.5005
R41963 VINP.n248 VINP.n158 4.5005
R41964 VINP.n336 VINP.n158 4.5005
R41965 VINP.n247 VINP.n158 4.5005
R41966 VINP.n338 VINP.n158 4.5005
R41967 VINP.n246 VINP.n158 4.5005
R41968 VINP.n340 VINP.n158 4.5005
R41969 VINP.n245 VINP.n158 4.5005
R41970 VINP.n342 VINP.n158 4.5005
R41971 VINP.n244 VINP.n158 4.5005
R41972 VINP.n344 VINP.n158 4.5005
R41973 VINP.n243 VINP.n158 4.5005
R41974 VINP.n346 VINP.n158 4.5005
R41975 VINP.n242 VINP.n158 4.5005
R41976 VINP.n348 VINP.n158 4.5005
R41977 VINP.n241 VINP.n158 4.5005
R41978 VINP.n350 VINP.n158 4.5005
R41979 VINP.n240 VINP.n158 4.5005
R41980 VINP.n352 VINP.n158 4.5005
R41981 VINP.n239 VINP.n158 4.5005
R41982 VINP.n354 VINP.n158 4.5005
R41983 VINP.n238 VINP.n158 4.5005
R41984 VINP.n356 VINP.n158 4.5005
R41985 VINP.n237 VINP.n158 4.5005
R41986 VINP.n358 VINP.n158 4.5005
R41987 VINP.n236 VINP.n158 4.5005
R41988 VINP.n360 VINP.n158 4.5005
R41989 VINP.n235 VINP.n158 4.5005
R41990 VINP.n362 VINP.n158 4.5005
R41991 VINP.n234 VINP.n158 4.5005
R41992 VINP.n364 VINP.n158 4.5005
R41993 VINP.n233 VINP.n158 4.5005
R41994 VINP.n366 VINP.n158 4.5005
R41995 VINP.n232 VINP.n158 4.5005
R41996 VINP.n368 VINP.n158 4.5005
R41997 VINP.n231 VINP.n158 4.5005
R41998 VINP.n370 VINP.n158 4.5005
R41999 VINP.n230 VINP.n158 4.5005
R42000 VINP.n372 VINP.n158 4.5005
R42001 VINP.n229 VINP.n158 4.5005
R42002 VINP.n374 VINP.n158 4.5005
R42003 VINP.n228 VINP.n158 4.5005
R42004 VINP.n376 VINP.n158 4.5005
R42005 VINP.n227 VINP.n158 4.5005
R42006 VINP.n378 VINP.n158 4.5005
R42007 VINP.n226 VINP.n158 4.5005
R42008 VINP.n380 VINP.n158 4.5005
R42009 VINP.n225 VINP.n158 4.5005
R42010 VINP.n382 VINP.n158 4.5005
R42011 VINP.n224 VINP.n158 4.5005
R42012 VINP.n384 VINP.n158 4.5005
R42013 VINP.n223 VINP.n158 4.5005
R42014 VINP.n386 VINP.n158 4.5005
R42015 VINP.n222 VINP.n158 4.5005
R42016 VINP.n388 VINP.n158 4.5005
R42017 VINP.n221 VINP.n158 4.5005
R42018 VINP.n390 VINP.n158 4.5005
R42019 VINP.n220 VINP.n158 4.5005
R42020 VINP.n392 VINP.n158 4.5005
R42021 VINP.n219 VINP.n158 4.5005
R42022 VINP.n394 VINP.n158 4.5005
R42023 VINP.n218 VINP.n158 4.5005
R42024 VINP.n396 VINP.n158 4.5005
R42025 VINP.n217 VINP.n158 4.5005
R42026 VINP.n398 VINP.n158 4.5005
R42027 VINP.n216 VINP.n158 4.5005
R42028 VINP.n400 VINP.n158 4.5005
R42029 VINP.n215 VINP.n158 4.5005
R42030 VINP.n654 VINP.n158 4.5005
R42031 VINP.n656 VINP.n158 4.5005
R42032 VINP.n158 VINP.n0 4.5005
R42033 VINP.n278 VINP.n142 4.5005
R42034 VINP.n276 VINP.n142 4.5005
R42035 VINP.n280 VINP.n142 4.5005
R42036 VINP.n275 VINP.n142 4.5005
R42037 VINP.n282 VINP.n142 4.5005
R42038 VINP.n274 VINP.n142 4.5005
R42039 VINP.n284 VINP.n142 4.5005
R42040 VINP.n273 VINP.n142 4.5005
R42041 VINP.n286 VINP.n142 4.5005
R42042 VINP.n272 VINP.n142 4.5005
R42043 VINP.n288 VINP.n142 4.5005
R42044 VINP.n271 VINP.n142 4.5005
R42045 VINP.n290 VINP.n142 4.5005
R42046 VINP.n270 VINP.n142 4.5005
R42047 VINP.n292 VINP.n142 4.5005
R42048 VINP.n269 VINP.n142 4.5005
R42049 VINP.n294 VINP.n142 4.5005
R42050 VINP.n268 VINP.n142 4.5005
R42051 VINP.n296 VINP.n142 4.5005
R42052 VINP.n267 VINP.n142 4.5005
R42053 VINP.n298 VINP.n142 4.5005
R42054 VINP.n266 VINP.n142 4.5005
R42055 VINP.n300 VINP.n142 4.5005
R42056 VINP.n265 VINP.n142 4.5005
R42057 VINP.n302 VINP.n142 4.5005
R42058 VINP.n264 VINP.n142 4.5005
R42059 VINP.n304 VINP.n142 4.5005
R42060 VINP.n263 VINP.n142 4.5005
R42061 VINP.n306 VINP.n142 4.5005
R42062 VINP.n262 VINP.n142 4.5005
R42063 VINP.n308 VINP.n142 4.5005
R42064 VINP.n261 VINP.n142 4.5005
R42065 VINP.n310 VINP.n142 4.5005
R42066 VINP.n260 VINP.n142 4.5005
R42067 VINP.n312 VINP.n142 4.5005
R42068 VINP.n259 VINP.n142 4.5005
R42069 VINP.n314 VINP.n142 4.5005
R42070 VINP.n258 VINP.n142 4.5005
R42071 VINP.n316 VINP.n142 4.5005
R42072 VINP.n257 VINP.n142 4.5005
R42073 VINP.n318 VINP.n142 4.5005
R42074 VINP.n256 VINP.n142 4.5005
R42075 VINP.n320 VINP.n142 4.5005
R42076 VINP.n255 VINP.n142 4.5005
R42077 VINP.n322 VINP.n142 4.5005
R42078 VINP.n254 VINP.n142 4.5005
R42079 VINP.n324 VINP.n142 4.5005
R42080 VINP.n253 VINP.n142 4.5005
R42081 VINP.n326 VINP.n142 4.5005
R42082 VINP.n252 VINP.n142 4.5005
R42083 VINP.n328 VINP.n142 4.5005
R42084 VINP.n251 VINP.n142 4.5005
R42085 VINP.n330 VINP.n142 4.5005
R42086 VINP.n250 VINP.n142 4.5005
R42087 VINP.n332 VINP.n142 4.5005
R42088 VINP.n249 VINP.n142 4.5005
R42089 VINP.n334 VINP.n142 4.5005
R42090 VINP.n248 VINP.n142 4.5005
R42091 VINP.n336 VINP.n142 4.5005
R42092 VINP.n247 VINP.n142 4.5005
R42093 VINP.n338 VINP.n142 4.5005
R42094 VINP.n246 VINP.n142 4.5005
R42095 VINP.n340 VINP.n142 4.5005
R42096 VINP.n245 VINP.n142 4.5005
R42097 VINP.n342 VINP.n142 4.5005
R42098 VINP.n244 VINP.n142 4.5005
R42099 VINP.n344 VINP.n142 4.5005
R42100 VINP.n243 VINP.n142 4.5005
R42101 VINP.n346 VINP.n142 4.5005
R42102 VINP.n242 VINP.n142 4.5005
R42103 VINP.n348 VINP.n142 4.5005
R42104 VINP.n241 VINP.n142 4.5005
R42105 VINP.n350 VINP.n142 4.5005
R42106 VINP.n240 VINP.n142 4.5005
R42107 VINP.n352 VINP.n142 4.5005
R42108 VINP.n239 VINP.n142 4.5005
R42109 VINP.n354 VINP.n142 4.5005
R42110 VINP.n238 VINP.n142 4.5005
R42111 VINP.n356 VINP.n142 4.5005
R42112 VINP.n237 VINP.n142 4.5005
R42113 VINP.n358 VINP.n142 4.5005
R42114 VINP.n236 VINP.n142 4.5005
R42115 VINP.n360 VINP.n142 4.5005
R42116 VINP.n235 VINP.n142 4.5005
R42117 VINP.n362 VINP.n142 4.5005
R42118 VINP.n234 VINP.n142 4.5005
R42119 VINP.n364 VINP.n142 4.5005
R42120 VINP.n233 VINP.n142 4.5005
R42121 VINP.n366 VINP.n142 4.5005
R42122 VINP.n232 VINP.n142 4.5005
R42123 VINP.n368 VINP.n142 4.5005
R42124 VINP.n231 VINP.n142 4.5005
R42125 VINP.n370 VINP.n142 4.5005
R42126 VINP.n230 VINP.n142 4.5005
R42127 VINP.n372 VINP.n142 4.5005
R42128 VINP.n229 VINP.n142 4.5005
R42129 VINP.n374 VINP.n142 4.5005
R42130 VINP.n228 VINP.n142 4.5005
R42131 VINP.n376 VINP.n142 4.5005
R42132 VINP.n227 VINP.n142 4.5005
R42133 VINP.n378 VINP.n142 4.5005
R42134 VINP.n226 VINP.n142 4.5005
R42135 VINP.n380 VINP.n142 4.5005
R42136 VINP.n225 VINP.n142 4.5005
R42137 VINP.n382 VINP.n142 4.5005
R42138 VINP.n224 VINP.n142 4.5005
R42139 VINP.n384 VINP.n142 4.5005
R42140 VINP.n223 VINP.n142 4.5005
R42141 VINP.n386 VINP.n142 4.5005
R42142 VINP.n222 VINP.n142 4.5005
R42143 VINP.n388 VINP.n142 4.5005
R42144 VINP.n221 VINP.n142 4.5005
R42145 VINP.n390 VINP.n142 4.5005
R42146 VINP.n220 VINP.n142 4.5005
R42147 VINP.n392 VINP.n142 4.5005
R42148 VINP.n219 VINP.n142 4.5005
R42149 VINP.n394 VINP.n142 4.5005
R42150 VINP.n218 VINP.n142 4.5005
R42151 VINP.n396 VINP.n142 4.5005
R42152 VINP.n217 VINP.n142 4.5005
R42153 VINP.n398 VINP.n142 4.5005
R42154 VINP.n216 VINP.n142 4.5005
R42155 VINP.n400 VINP.n142 4.5005
R42156 VINP.n215 VINP.n142 4.5005
R42157 VINP.n654 VINP.n142 4.5005
R42158 VINP.n656 VINP.n142 4.5005
R42159 VINP.n142 VINP.n0 4.5005
R42160 VINP.n278 VINP.n159 4.5005
R42161 VINP.n276 VINP.n159 4.5005
R42162 VINP.n280 VINP.n159 4.5005
R42163 VINP.n275 VINP.n159 4.5005
R42164 VINP.n282 VINP.n159 4.5005
R42165 VINP.n274 VINP.n159 4.5005
R42166 VINP.n284 VINP.n159 4.5005
R42167 VINP.n273 VINP.n159 4.5005
R42168 VINP.n286 VINP.n159 4.5005
R42169 VINP.n272 VINP.n159 4.5005
R42170 VINP.n288 VINP.n159 4.5005
R42171 VINP.n271 VINP.n159 4.5005
R42172 VINP.n290 VINP.n159 4.5005
R42173 VINP.n270 VINP.n159 4.5005
R42174 VINP.n292 VINP.n159 4.5005
R42175 VINP.n269 VINP.n159 4.5005
R42176 VINP.n294 VINP.n159 4.5005
R42177 VINP.n268 VINP.n159 4.5005
R42178 VINP.n296 VINP.n159 4.5005
R42179 VINP.n267 VINP.n159 4.5005
R42180 VINP.n298 VINP.n159 4.5005
R42181 VINP.n266 VINP.n159 4.5005
R42182 VINP.n300 VINP.n159 4.5005
R42183 VINP.n265 VINP.n159 4.5005
R42184 VINP.n302 VINP.n159 4.5005
R42185 VINP.n264 VINP.n159 4.5005
R42186 VINP.n304 VINP.n159 4.5005
R42187 VINP.n263 VINP.n159 4.5005
R42188 VINP.n306 VINP.n159 4.5005
R42189 VINP.n262 VINP.n159 4.5005
R42190 VINP.n308 VINP.n159 4.5005
R42191 VINP.n261 VINP.n159 4.5005
R42192 VINP.n310 VINP.n159 4.5005
R42193 VINP.n260 VINP.n159 4.5005
R42194 VINP.n312 VINP.n159 4.5005
R42195 VINP.n259 VINP.n159 4.5005
R42196 VINP.n314 VINP.n159 4.5005
R42197 VINP.n258 VINP.n159 4.5005
R42198 VINP.n316 VINP.n159 4.5005
R42199 VINP.n257 VINP.n159 4.5005
R42200 VINP.n318 VINP.n159 4.5005
R42201 VINP.n256 VINP.n159 4.5005
R42202 VINP.n320 VINP.n159 4.5005
R42203 VINP.n255 VINP.n159 4.5005
R42204 VINP.n322 VINP.n159 4.5005
R42205 VINP.n254 VINP.n159 4.5005
R42206 VINP.n324 VINP.n159 4.5005
R42207 VINP.n253 VINP.n159 4.5005
R42208 VINP.n326 VINP.n159 4.5005
R42209 VINP.n252 VINP.n159 4.5005
R42210 VINP.n328 VINP.n159 4.5005
R42211 VINP.n251 VINP.n159 4.5005
R42212 VINP.n330 VINP.n159 4.5005
R42213 VINP.n250 VINP.n159 4.5005
R42214 VINP.n332 VINP.n159 4.5005
R42215 VINP.n249 VINP.n159 4.5005
R42216 VINP.n334 VINP.n159 4.5005
R42217 VINP.n248 VINP.n159 4.5005
R42218 VINP.n336 VINP.n159 4.5005
R42219 VINP.n247 VINP.n159 4.5005
R42220 VINP.n338 VINP.n159 4.5005
R42221 VINP.n246 VINP.n159 4.5005
R42222 VINP.n340 VINP.n159 4.5005
R42223 VINP.n245 VINP.n159 4.5005
R42224 VINP.n342 VINP.n159 4.5005
R42225 VINP.n244 VINP.n159 4.5005
R42226 VINP.n344 VINP.n159 4.5005
R42227 VINP.n243 VINP.n159 4.5005
R42228 VINP.n346 VINP.n159 4.5005
R42229 VINP.n242 VINP.n159 4.5005
R42230 VINP.n348 VINP.n159 4.5005
R42231 VINP.n241 VINP.n159 4.5005
R42232 VINP.n350 VINP.n159 4.5005
R42233 VINP.n240 VINP.n159 4.5005
R42234 VINP.n352 VINP.n159 4.5005
R42235 VINP.n239 VINP.n159 4.5005
R42236 VINP.n354 VINP.n159 4.5005
R42237 VINP.n238 VINP.n159 4.5005
R42238 VINP.n356 VINP.n159 4.5005
R42239 VINP.n237 VINP.n159 4.5005
R42240 VINP.n358 VINP.n159 4.5005
R42241 VINP.n236 VINP.n159 4.5005
R42242 VINP.n360 VINP.n159 4.5005
R42243 VINP.n235 VINP.n159 4.5005
R42244 VINP.n362 VINP.n159 4.5005
R42245 VINP.n234 VINP.n159 4.5005
R42246 VINP.n364 VINP.n159 4.5005
R42247 VINP.n233 VINP.n159 4.5005
R42248 VINP.n366 VINP.n159 4.5005
R42249 VINP.n232 VINP.n159 4.5005
R42250 VINP.n368 VINP.n159 4.5005
R42251 VINP.n231 VINP.n159 4.5005
R42252 VINP.n370 VINP.n159 4.5005
R42253 VINP.n230 VINP.n159 4.5005
R42254 VINP.n372 VINP.n159 4.5005
R42255 VINP.n229 VINP.n159 4.5005
R42256 VINP.n374 VINP.n159 4.5005
R42257 VINP.n228 VINP.n159 4.5005
R42258 VINP.n376 VINP.n159 4.5005
R42259 VINP.n227 VINP.n159 4.5005
R42260 VINP.n378 VINP.n159 4.5005
R42261 VINP.n226 VINP.n159 4.5005
R42262 VINP.n380 VINP.n159 4.5005
R42263 VINP.n225 VINP.n159 4.5005
R42264 VINP.n382 VINP.n159 4.5005
R42265 VINP.n224 VINP.n159 4.5005
R42266 VINP.n384 VINP.n159 4.5005
R42267 VINP.n223 VINP.n159 4.5005
R42268 VINP.n386 VINP.n159 4.5005
R42269 VINP.n222 VINP.n159 4.5005
R42270 VINP.n388 VINP.n159 4.5005
R42271 VINP.n221 VINP.n159 4.5005
R42272 VINP.n390 VINP.n159 4.5005
R42273 VINP.n220 VINP.n159 4.5005
R42274 VINP.n392 VINP.n159 4.5005
R42275 VINP.n219 VINP.n159 4.5005
R42276 VINP.n394 VINP.n159 4.5005
R42277 VINP.n218 VINP.n159 4.5005
R42278 VINP.n396 VINP.n159 4.5005
R42279 VINP.n217 VINP.n159 4.5005
R42280 VINP.n398 VINP.n159 4.5005
R42281 VINP.n216 VINP.n159 4.5005
R42282 VINP.n400 VINP.n159 4.5005
R42283 VINP.n215 VINP.n159 4.5005
R42284 VINP.n654 VINP.n159 4.5005
R42285 VINP.n656 VINP.n159 4.5005
R42286 VINP.n159 VINP.n0 4.5005
R42287 VINP.n278 VINP.n141 4.5005
R42288 VINP.n276 VINP.n141 4.5005
R42289 VINP.n280 VINP.n141 4.5005
R42290 VINP.n275 VINP.n141 4.5005
R42291 VINP.n282 VINP.n141 4.5005
R42292 VINP.n274 VINP.n141 4.5005
R42293 VINP.n284 VINP.n141 4.5005
R42294 VINP.n273 VINP.n141 4.5005
R42295 VINP.n286 VINP.n141 4.5005
R42296 VINP.n272 VINP.n141 4.5005
R42297 VINP.n288 VINP.n141 4.5005
R42298 VINP.n271 VINP.n141 4.5005
R42299 VINP.n290 VINP.n141 4.5005
R42300 VINP.n270 VINP.n141 4.5005
R42301 VINP.n292 VINP.n141 4.5005
R42302 VINP.n269 VINP.n141 4.5005
R42303 VINP.n294 VINP.n141 4.5005
R42304 VINP.n268 VINP.n141 4.5005
R42305 VINP.n296 VINP.n141 4.5005
R42306 VINP.n267 VINP.n141 4.5005
R42307 VINP.n298 VINP.n141 4.5005
R42308 VINP.n266 VINP.n141 4.5005
R42309 VINP.n300 VINP.n141 4.5005
R42310 VINP.n265 VINP.n141 4.5005
R42311 VINP.n302 VINP.n141 4.5005
R42312 VINP.n264 VINP.n141 4.5005
R42313 VINP.n304 VINP.n141 4.5005
R42314 VINP.n263 VINP.n141 4.5005
R42315 VINP.n306 VINP.n141 4.5005
R42316 VINP.n262 VINP.n141 4.5005
R42317 VINP.n308 VINP.n141 4.5005
R42318 VINP.n261 VINP.n141 4.5005
R42319 VINP.n310 VINP.n141 4.5005
R42320 VINP.n260 VINP.n141 4.5005
R42321 VINP.n312 VINP.n141 4.5005
R42322 VINP.n259 VINP.n141 4.5005
R42323 VINP.n314 VINP.n141 4.5005
R42324 VINP.n258 VINP.n141 4.5005
R42325 VINP.n316 VINP.n141 4.5005
R42326 VINP.n257 VINP.n141 4.5005
R42327 VINP.n318 VINP.n141 4.5005
R42328 VINP.n256 VINP.n141 4.5005
R42329 VINP.n320 VINP.n141 4.5005
R42330 VINP.n255 VINP.n141 4.5005
R42331 VINP.n322 VINP.n141 4.5005
R42332 VINP.n254 VINP.n141 4.5005
R42333 VINP.n324 VINP.n141 4.5005
R42334 VINP.n253 VINP.n141 4.5005
R42335 VINP.n326 VINP.n141 4.5005
R42336 VINP.n252 VINP.n141 4.5005
R42337 VINP.n328 VINP.n141 4.5005
R42338 VINP.n251 VINP.n141 4.5005
R42339 VINP.n330 VINP.n141 4.5005
R42340 VINP.n250 VINP.n141 4.5005
R42341 VINP.n332 VINP.n141 4.5005
R42342 VINP.n249 VINP.n141 4.5005
R42343 VINP.n334 VINP.n141 4.5005
R42344 VINP.n248 VINP.n141 4.5005
R42345 VINP.n336 VINP.n141 4.5005
R42346 VINP.n247 VINP.n141 4.5005
R42347 VINP.n338 VINP.n141 4.5005
R42348 VINP.n246 VINP.n141 4.5005
R42349 VINP.n340 VINP.n141 4.5005
R42350 VINP.n245 VINP.n141 4.5005
R42351 VINP.n342 VINP.n141 4.5005
R42352 VINP.n244 VINP.n141 4.5005
R42353 VINP.n344 VINP.n141 4.5005
R42354 VINP.n243 VINP.n141 4.5005
R42355 VINP.n346 VINP.n141 4.5005
R42356 VINP.n242 VINP.n141 4.5005
R42357 VINP.n348 VINP.n141 4.5005
R42358 VINP.n241 VINP.n141 4.5005
R42359 VINP.n350 VINP.n141 4.5005
R42360 VINP.n240 VINP.n141 4.5005
R42361 VINP.n352 VINP.n141 4.5005
R42362 VINP.n239 VINP.n141 4.5005
R42363 VINP.n354 VINP.n141 4.5005
R42364 VINP.n238 VINP.n141 4.5005
R42365 VINP.n356 VINP.n141 4.5005
R42366 VINP.n237 VINP.n141 4.5005
R42367 VINP.n358 VINP.n141 4.5005
R42368 VINP.n236 VINP.n141 4.5005
R42369 VINP.n360 VINP.n141 4.5005
R42370 VINP.n235 VINP.n141 4.5005
R42371 VINP.n362 VINP.n141 4.5005
R42372 VINP.n234 VINP.n141 4.5005
R42373 VINP.n364 VINP.n141 4.5005
R42374 VINP.n233 VINP.n141 4.5005
R42375 VINP.n366 VINP.n141 4.5005
R42376 VINP.n232 VINP.n141 4.5005
R42377 VINP.n368 VINP.n141 4.5005
R42378 VINP.n231 VINP.n141 4.5005
R42379 VINP.n370 VINP.n141 4.5005
R42380 VINP.n230 VINP.n141 4.5005
R42381 VINP.n372 VINP.n141 4.5005
R42382 VINP.n229 VINP.n141 4.5005
R42383 VINP.n374 VINP.n141 4.5005
R42384 VINP.n228 VINP.n141 4.5005
R42385 VINP.n376 VINP.n141 4.5005
R42386 VINP.n227 VINP.n141 4.5005
R42387 VINP.n378 VINP.n141 4.5005
R42388 VINP.n226 VINP.n141 4.5005
R42389 VINP.n380 VINP.n141 4.5005
R42390 VINP.n225 VINP.n141 4.5005
R42391 VINP.n382 VINP.n141 4.5005
R42392 VINP.n224 VINP.n141 4.5005
R42393 VINP.n384 VINP.n141 4.5005
R42394 VINP.n223 VINP.n141 4.5005
R42395 VINP.n386 VINP.n141 4.5005
R42396 VINP.n222 VINP.n141 4.5005
R42397 VINP.n388 VINP.n141 4.5005
R42398 VINP.n221 VINP.n141 4.5005
R42399 VINP.n390 VINP.n141 4.5005
R42400 VINP.n220 VINP.n141 4.5005
R42401 VINP.n392 VINP.n141 4.5005
R42402 VINP.n219 VINP.n141 4.5005
R42403 VINP.n394 VINP.n141 4.5005
R42404 VINP.n218 VINP.n141 4.5005
R42405 VINP.n396 VINP.n141 4.5005
R42406 VINP.n217 VINP.n141 4.5005
R42407 VINP.n398 VINP.n141 4.5005
R42408 VINP.n216 VINP.n141 4.5005
R42409 VINP.n400 VINP.n141 4.5005
R42410 VINP.n215 VINP.n141 4.5005
R42411 VINP.n654 VINP.n141 4.5005
R42412 VINP.n656 VINP.n141 4.5005
R42413 VINP.n141 VINP.n0 4.5005
R42414 VINP.n278 VINP.n160 4.5005
R42415 VINP.n276 VINP.n160 4.5005
R42416 VINP.n280 VINP.n160 4.5005
R42417 VINP.n275 VINP.n160 4.5005
R42418 VINP.n282 VINP.n160 4.5005
R42419 VINP.n274 VINP.n160 4.5005
R42420 VINP.n284 VINP.n160 4.5005
R42421 VINP.n273 VINP.n160 4.5005
R42422 VINP.n286 VINP.n160 4.5005
R42423 VINP.n272 VINP.n160 4.5005
R42424 VINP.n288 VINP.n160 4.5005
R42425 VINP.n271 VINP.n160 4.5005
R42426 VINP.n290 VINP.n160 4.5005
R42427 VINP.n270 VINP.n160 4.5005
R42428 VINP.n292 VINP.n160 4.5005
R42429 VINP.n269 VINP.n160 4.5005
R42430 VINP.n294 VINP.n160 4.5005
R42431 VINP.n268 VINP.n160 4.5005
R42432 VINP.n296 VINP.n160 4.5005
R42433 VINP.n267 VINP.n160 4.5005
R42434 VINP.n298 VINP.n160 4.5005
R42435 VINP.n266 VINP.n160 4.5005
R42436 VINP.n300 VINP.n160 4.5005
R42437 VINP.n265 VINP.n160 4.5005
R42438 VINP.n302 VINP.n160 4.5005
R42439 VINP.n264 VINP.n160 4.5005
R42440 VINP.n304 VINP.n160 4.5005
R42441 VINP.n263 VINP.n160 4.5005
R42442 VINP.n306 VINP.n160 4.5005
R42443 VINP.n262 VINP.n160 4.5005
R42444 VINP.n308 VINP.n160 4.5005
R42445 VINP.n261 VINP.n160 4.5005
R42446 VINP.n310 VINP.n160 4.5005
R42447 VINP.n260 VINP.n160 4.5005
R42448 VINP.n312 VINP.n160 4.5005
R42449 VINP.n259 VINP.n160 4.5005
R42450 VINP.n314 VINP.n160 4.5005
R42451 VINP.n258 VINP.n160 4.5005
R42452 VINP.n316 VINP.n160 4.5005
R42453 VINP.n257 VINP.n160 4.5005
R42454 VINP.n318 VINP.n160 4.5005
R42455 VINP.n256 VINP.n160 4.5005
R42456 VINP.n320 VINP.n160 4.5005
R42457 VINP.n255 VINP.n160 4.5005
R42458 VINP.n322 VINP.n160 4.5005
R42459 VINP.n254 VINP.n160 4.5005
R42460 VINP.n324 VINP.n160 4.5005
R42461 VINP.n253 VINP.n160 4.5005
R42462 VINP.n326 VINP.n160 4.5005
R42463 VINP.n252 VINP.n160 4.5005
R42464 VINP.n328 VINP.n160 4.5005
R42465 VINP.n251 VINP.n160 4.5005
R42466 VINP.n330 VINP.n160 4.5005
R42467 VINP.n250 VINP.n160 4.5005
R42468 VINP.n332 VINP.n160 4.5005
R42469 VINP.n249 VINP.n160 4.5005
R42470 VINP.n334 VINP.n160 4.5005
R42471 VINP.n248 VINP.n160 4.5005
R42472 VINP.n336 VINP.n160 4.5005
R42473 VINP.n247 VINP.n160 4.5005
R42474 VINP.n338 VINP.n160 4.5005
R42475 VINP.n246 VINP.n160 4.5005
R42476 VINP.n340 VINP.n160 4.5005
R42477 VINP.n245 VINP.n160 4.5005
R42478 VINP.n342 VINP.n160 4.5005
R42479 VINP.n244 VINP.n160 4.5005
R42480 VINP.n344 VINP.n160 4.5005
R42481 VINP.n243 VINP.n160 4.5005
R42482 VINP.n346 VINP.n160 4.5005
R42483 VINP.n242 VINP.n160 4.5005
R42484 VINP.n348 VINP.n160 4.5005
R42485 VINP.n241 VINP.n160 4.5005
R42486 VINP.n350 VINP.n160 4.5005
R42487 VINP.n240 VINP.n160 4.5005
R42488 VINP.n352 VINP.n160 4.5005
R42489 VINP.n239 VINP.n160 4.5005
R42490 VINP.n354 VINP.n160 4.5005
R42491 VINP.n238 VINP.n160 4.5005
R42492 VINP.n356 VINP.n160 4.5005
R42493 VINP.n237 VINP.n160 4.5005
R42494 VINP.n358 VINP.n160 4.5005
R42495 VINP.n236 VINP.n160 4.5005
R42496 VINP.n360 VINP.n160 4.5005
R42497 VINP.n235 VINP.n160 4.5005
R42498 VINP.n362 VINP.n160 4.5005
R42499 VINP.n234 VINP.n160 4.5005
R42500 VINP.n364 VINP.n160 4.5005
R42501 VINP.n233 VINP.n160 4.5005
R42502 VINP.n366 VINP.n160 4.5005
R42503 VINP.n232 VINP.n160 4.5005
R42504 VINP.n368 VINP.n160 4.5005
R42505 VINP.n231 VINP.n160 4.5005
R42506 VINP.n370 VINP.n160 4.5005
R42507 VINP.n230 VINP.n160 4.5005
R42508 VINP.n372 VINP.n160 4.5005
R42509 VINP.n229 VINP.n160 4.5005
R42510 VINP.n374 VINP.n160 4.5005
R42511 VINP.n228 VINP.n160 4.5005
R42512 VINP.n376 VINP.n160 4.5005
R42513 VINP.n227 VINP.n160 4.5005
R42514 VINP.n378 VINP.n160 4.5005
R42515 VINP.n226 VINP.n160 4.5005
R42516 VINP.n380 VINP.n160 4.5005
R42517 VINP.n225 VINP.n160 4.5005
R42518 VINP.n382 VINP.n160 4.5005
R42519 VINP.n224 VINP.n160 4.5005
R42520 VINP.n384 VINP.n160 4.5005
R42521 VINP.n223 VINP.n160 4.5005
R42522 VINP.n386 VINP.n160 4.5005
R42523 VINP.n222 VINP.n160 4.5005
R42524 VINP.n388 VINP.n160 4.5005
R42525 VINP.n221 VINP.n160 4.5005
R42526 VINP.n390 VINP.n160 4.5005
R42527 VINP.n220 VINP.n160 4.5005
R42528 VINP.n392 VINP.n160 4.5005
R42529 VINP.n219 VINP.n160 4.5005
R42530 VINP.n394 VINP.n160 4.5005
R42531 VINP.n218 VINP.n160 4.5005
R42532 VINP.n396 VINP.n160 4.5005
R42533 VINP.n217 VINP.n160 4.5005
R42534 VINP.n398 VINP.n160 4.5005
R42535 VINP.n216 VINP.n160 4.5005
R42536 VINP.n400 VINP.n160 4.5005
R42537 VINP.n215 VINP.n160 4.5005
R42538 VINP.n654 VINP.n160 4.5005
R42539 VINP.n656 VINP.n160 4.5005
R42540 VINP.n160 VINP.n0 4.5005
R42541 VINP.n278 VINP.n140 4.5005
R42542 VINP.n276 VINP.n140 4.5005
R42543 VINP.n280 VINP.n140 4.5005
R42544 VINP.n275 VINP.n140 4.5005
R42545 VINP.n282 VINP.n140 4.5005
R42546 VINP.n274 VINP.n140 4.5005
R42547 VINP.n284 VINP.n140 4.5005
R42548 VINP.n273 VINP.n140 4.5005
R42549 VINP.n286 VINP.n140 4.5005
R42550 VINP.n272 VINP.n140 4.5005
R42551 VINP.n288 VINP.n140 4.5005
R42552 VINP.n271 VINP.n140 4.5005
R42553 VINP.n290 VINP.n140 4.5005
R42554 VINP.n270 VINP.n140 4.5005
R42555 VINP.n292 VINP.n140 4.5005
R42556 VINP.n269 VINP.n140 4.5005
R42557 VINP.n294 VINP.n140 4.5005
R42558 VINP.n268 VINP.n140 4.5005
R42559 VINP.n296 VINP.n140 4.5005
R42560 VINP.n267 VINP.n140 4.5005
R42561 VINP.n298 VINP.n140 4.5005
R42562 VINP.n266 VINP.n140 4.5005
R42563 VINP.n300 VINP.n140 4.5005
R42564 VINP.n265 VINP.n140 4.5005
R42565 VINP.n302 VINP.n140 4.5005
R42566 VINP.n264 VINP.n140 4.5005
R42567 VINP.n304 VINP.n140 4.5005
R42568 VINP.n263 VINP.n140 4.5005
R42569 VINP.n306 VINP.n140 4.5005
R42570 VINP.n262 VINP.n140 4.5005
R42571 VINP.n308 VINP.n140 4.5005
R42572 VINP.n261 VINP.n140 4.5005
R42573 VINP.n310 VINP.n140 4.5005
R42574 VINP.n260 VINP.n140 4.5005
R42575 VINP.n312 VINP.n140 4.5005
R42576 VINP.n259 VINP.n140 4.5005
R42577 VINP.n314 VINP.n140 4.5005
R42578 VINP.n258 VINP.n140 4.5005
R42579 VINP.n316 VINP.n140 4.5005
R42580 VINP.n257 VINP.n140 4.5005
R42581 VINP.n318 VINP.n140 4.5005
R42582 VINP.n256 VINP.n140 4.5005
R42583 VINP.n320 VINP.n140 4.5005
R42584 VINP.n255 VINP.n140 4.5005
R42585 VINP.n322 VINP.n140 4.5005
R42586 VINP.n254 VINP.n140 4.5005
R42587 VINP.n324 VINP.n140 4.5005
R42588 VINP.n253 VINP.n140 4.5005
R42589 VINP.n326 VINP.n140 4.5005
R42590 VINP.n252 VINP.n140 4.5005
R42591 VINP.n328 VINP.n140 4.5005
R42592 VINP.n251 VINP.n140 4.5005
R42593 VINP.n330 VINP.n140 4.5005
R42594 VINP.n250 VINP.n140 4.5005
R42595 VINP.n332 VINP.n140 4.5005
R42596 VINP.n249 VINP.n140 4.5005
R42597 VINP.n334 VINP.n140 4.5005
R42598 VINP.n248 VINP.n140 4.5005
R42599 VINP.n336 VINP.n140 4.5005
R42600 VINP.n247 VINP.n140 4.5005
R42601 VINP.n338 VINP.n140 4.5005
R42602 VINP.n246 VINP.n140 4.5005
R42603 VINP.n340 VINP.n140 4.5005
R42604 VINP.n245 VINP.n140 4.5005
R42605 VINP.n342 VINP.n140 4.5005
R42606 VINP.n244 VINP.n140 4.5005
R42607 VINP.n344 VINP.n140 4.5005
R42608 VINP.n243 VINP.n140 4.5005
R42609 VINP.n346 VINP.n140 4.5005
R42610 VINP.n242 VINP.n140 4.5005
R42611 VINP.n348 VINP.n140 4.5005
R42612 VINP.n241 VINP.n140 4.5005
R42613 VINP.n350 VINP.n140 4.5005
R42614 VINP.n240 VINP.n140 4.5005
R42615 VINP.n352 VINP.n140 4.5005
R42616 VINP.n239 VINP.n140 4.5005
R42617 VINP.n354 VINP.n140 4.5005
R42618 VINP.n238 VINP.n140 4.5005
R42619 VINP.n356 VINP.n140 4.5005
R42620 VINP.n237 VINP.n140 4.5005
R42621 VINP.n358 VINP.n140 4.5005
R42622 VINP.n236 VINP.n140 4.5005
R42623 VINP.n360 VINP.n140 4.5005
R42624 VINP.n235 VINP.n140 4.5005
R42625 VINP.n362 VINP.n140 4.5005
R42626 VINP.n234 VINP.n140 4.5005
R42627 VINP.n364 VINP.n140 4.5005
R42628 VINP.n233 VINP.n140 4.5005
R42629 VINP.n366 VINP.n140 4.5005
R42630 VINP.n232 VINP.n140 4.5005
R42631 VINP.n368 VINP.n140 4.5005
R42632 VINP.n231 VINP.n140 4.5005
R42633 VINP.n370 VINP.n140 4.5005
R42634 VINP.n230 VINP.n140 4.5005
R42635 VINP.n372 VINP.n140 4.5005
R42636 VINP.n229 VINP.n140 4.5005
R42637 VINP.n374 VINP.n140 4.5005
R42638 VINP.n228 VINP.n140 4.5005
R42639 VINP.n376 VINP.n140 4.5005
R42640 VINP.n227 VINP.n140 4.5005
R42641 VINP.n378 VINP.n140 4.5005
R42642 VINP.n226 VINP.n140 4.5005
R42643 VINP.n380 VINP.n140 4.5005
R42644 VINP.n225 VINP.n140 4.5005
R42645 VINP.n382 VINP.n140 4.5005
R42646 VINP.n224 VINP.n140 4.5005
R42647 VINP.n384 VINP.n140 4.5005
R42648 VINP.n223 VINP.n140 4.5005
R42649 VINP.n386 VINP.n140 4.5005
R42650 VINP.n222 VINP.n140 4.5005
R42651 VINP.n388 VINP.n140 4.5005
R42652 VINP.n221 VINP.n140 4.5005
R42653 VINP.n390 VINP.n140 4.5005
R42654 VINP.n220 VINP.n140 4.5005
R42655 VINP.n392 VINP.n140 4.5005
R42656 VINP.n219 VINP.n140 4.5005
R42657 VINP.n394 VINP.n140 4.5005
R42658 VINP.n218 VINP.n140 4.5005
R42659 VINP.n396 VINP.n140 4.5005
R42660 VINP.n217 VINP.n140 4.5005
R42661 VINP.n398 VINP.n140 4.5005
R42662 VINP.n216 VINP.n140 4.5005
R42663 VINP.n400 VINP.n140 4.5005
R42664 VINP.n215 VINP.n140 4.5005
R42665 VINP.n654 VINP.n140 4.5005
R42666 VINP.n656 VINP.n140 4.5005
R42667 VINP.n140 VINP.n0 4.5005
R42668 VINP.n278 VINP.n161 4.5005
R42669 VINP.n276 VINP.n161 4.5005
R42670 VINP.n280 VINP.n161 4.5005
R42671 VINP.n275 VINP.n161 4.5005
R42672 VINP.n282 VINP.n161 4.5005
R42673 VINP.n274 VINP.n161 4.5005
R42674 VINP.n284 VINP.n161 4.5005
R42675 VINP.n273 VINP.n161 4.5005
R42676 VINP.n286 VINP.n161 4.5005
R42677 VINP.n272 VINP.n161 4.5005
R42678 VINP.n288 VINP.n161 4.5005
R42679 VINP.n271 VINP.n161 4.5005
R42680 VINP.n290 VINP.n161 4.5005
R42681 VINP.n270 VINP.n161 4.5005
R42682 VINP.n292 VINP.n161 4.5005
R42683 VINP.n269 VINP.n161 4.5005
R42684 VINP.n294 VINP.n161 4.5005
R42685 VINP.n268 VINP.n161 4.5005
R42686 VINP.n296 VINP.n161 4.5005
R42687 VINP.n267 VINP.n161 4.5005
R42688 VINP.n298 VINP.n161 4.5005
R42689 VINP.n266 VINP.n161 4.5005
R42690 VINP.n300 VINP.n161 4.5005
R42691 VINP.n265 VINP.n161 4.5005
R42692 VINP.n302 VINP.n161 4.5005
R42693 VINP.n264 VINP.n161 4.5005
R42694 VINP.n304 VINP.n161 4.5005
R42695 VINP.n263 VINP.n161 4.5005
R42696 VINP.n306 VINP.n161 4.5005
R42697 VINP.n262 VINP.n161 4.5005
R42698 VINP.n308 VINP.n161 4.5005
R42699 VINP.n261 VINP.n161 4.5005
R42700 VINP.n310 VINP.n161 4.5005
R42701 VINP.n260 VINP.n161 4.5005
R42702 VINP.n312 VINP.n161 4.5005
R42703 VINP.n259 VINP.n161 4.5005
R42704 VINP.n314 VINP.n161 4.5005
R42705 VINP.n258 VINP.n161 4.5005
R42706 VINP.n316 VINP.n161 4.5005
R42707 VINP.n257 VINP.n161 4.5005
R42708 VINP.n318 VINP.n161 4.5005
R42709 VINP.n256 VINP.n161 4.5005
R42710 VINP.n320 VINP.n161 4.5005
R42711 VINP.n255 VINP.n161 4.5005
R42712 VINP.n322 VINP.n161 4.5005
R42713 VINP.n254 VINP.n161 4.5005
R42714 VINP.n324 VINP.n161 4.5005
R42715 VINP.n253 VINP.n161 4.5005
R42716 VINP.n326 VINP.n161 4.5005
R42717 VINP.n252 VINP.n161 4.5005
R42718 VINP.n328 VINP.n161 4.5005
R42719 VINP.n251 VINP.n161 4.5005
R42720 VINP.n330 VINP.n161 4.5005
R42721 VINP.n250 VINP.n161 4.5005
R42722 VINP.n332 VINP.n161 4.5005
R42723 VINP.n249 VINP.n161 4.5005
R42724 VINP.n334 VINP.n161 4.5005
R42725 VINP.n248 VINP.n161 4.5005
R42726 VINP.n336 VINP.n161 4.5005
R42727 VINP.n247 VINP.n161 4.5005
R42728 VINP.n338 VINP.n161 4.5005
R42729 VINP.n246 VINP.n161 4.5005
R42730 VINP.n340 VINP.n161 4.5005
R42731 VINP.n245 VINP.n161 4.5005
R42732 VINP.n342 VINP.n161 4.5005
R42733 VINP.n244 VINP.n161 4.5005
R42734 VINP.n344 VINP.n161 4.5005
R42735 VINP.n243 VINP.n161 4.5005
R42736 VINP.n346 VINP.n161 4.5005
R42737 VINP.n242 VINP.n161 4.5005
R42738 VINP.n348 VINP.n161 4.5005
R42739 VINP.n241 VINP.n161 4.5005
R42740 VINP.n350 VINP.n161 4.5005
R42741 VINP.n240 VINP.n161 4.5005
R42742 VINP.n352 VINP.n161 4.5005
R42743 VINP.n239 VINP.n161 4.5005
R42744 VINP.n354 VINP.n161 4.5005
R42745 VINP.n238 VINP.n161 4.5005
R42746 VINP.n356 VINP.n161 4.5005
R42747 VINP.n237 VINP.n161 4.5005
R42748 VINP.n358 VINP.n161 4.5005
R42749 VINP.n236 VINP.n161 4.5005
R42750 VINP.n360 VINP.n161 4.5005
R42751 VINP.n235 VINP.n161 4.5005
R42752 VINP.n362 VINP.n161 4.5005
R42753 VINP.n234 VINP.n161 4.5005
R42754 VINP.n364 VINP.n161 4.5005
R42755 VINP.n233 VINP.n161 4.5005
R42756 VINP.n366 VINP.n161 4.5005
R42757 VINP.n232 VINP.n161 4.5005
R42758 VINP.n368 VINP.n161 4.5005
R42759 VINP.n231 VINP.n161 4.5005
R42760 VINP.n370 VINP.n161 4.5005
R42761 VINP.n230 VINP.n161 4.5005
R42762 VINP.n372 VINP.n161 4.5005
R42763 VINP.n229 VINP.n161 4.5005
R42764 VINP.n374 VINP.n161 4.5005
R42765 VINP.n228 VINP.n161 4.5005
R42766 VINP.n376 VINP.n161 4.5005
R42767 VINP.n227 VINP.n161 4.5005
R42768 VINP.n378 VINP.n161 4.5005
R42769 VINP.n226 VINP.n161 4.5005
R42770 VINP.n380 VINP.n161 4.5005
R42771 VINP.n225 VINP.n161 4.5005
R42772 VINP.n382 VINP.n161 4.5005
R42773 VINP.n224 VINP.n161 4.5005
R42774 VINP.n384 VINP.n161 4.5005
R42775 VINP.n223 VINP.n161 4.5005
R42776 VINP.n386 VINP.n161 4.5005
R42777 VINP.n222 VINP.n161 4.5005
R42778 VINP.n388 VINP.n161 4.5005
R42779 VINP.n221 VINP.n161 4.5005
R42780 VINP.n390 VINP.n161 4.5005
R42781 VINP.n220 VINP.n161 4.5005
R42782 VINP.n392 VINP.n161 4.5005
R42783 VINP.n219 VINP.n161 4.5005
R42784 VINP.n394 VINP.n161 4.5005
R42785 VINP.n218 VINP.n161 4.5005
R42786 VINP.n396 VINP.n161 4.5005
R42787 VINP.n217 VINP.n161 4.5005
R42788 VINP.n398 VINP.n161 4.5005
R42789 VINP.n216 VINP.n161 4.5005
R42790 VINP.n400 VINP.n161 4.5005
R42791 VINP.n215 VINP.n161 4.5005
R42792 VINP.n654 VINP.n161 4.5005
R42793 VINP.n656 VINP.n161 4.5005
R42794 VINP.n161 VINP.n0 4.5005
R42795 VINP.n278 VINP.n139 4.5005
R42796 VINP.n276 VINP.n139 4.5005
R42797 VINP.n280 VINP.n139 4.5005
R42798 VINP.n275 VINP.n139 4.5005
R42799 VINP.n282 VINP.n139 4.5005
R42800 VINP.n274 VINP.n139 4.5005
R42801 VINP.n284 VINP.n139 4.5005
R42802 VINP.n273 VINP.n139 4.5005
R42803 VINP.n286 VINP.n139 4.5005
R42804 VINP.n272 VINP.n139 4.5005
R42805 VINP.n288 VINP.n139 4.5005
R42806 VINP.n271 VINP.n139 4.5005
R42807 VINP.n290 VINP.n139 4.5005
R42808 VINP.n270 VINP.n139 4.5005
R42809 VINP.n292 VINP.n139 4.5005
R42810 VINP.n269 VINP.n139 4.5005
R42811 VINP.n294 VINP.n139 4.5005
R42812 VINP.n268 VINP.n139 4.5005
R42813 VINP.n296 VINP.n139 4.5005
R42814 VINP.n267 VINP.n139 4.5005
R42815 VINP.n298 VINP.n139 4.5005
R42816 VINP.n266 VINP.n139 4.5005
R42817 VINP.n300 VINP.n139 4.5005
R42818 VINP.n265 VINP.n139 4.5005
R42819 VINP.n302 VINP.n139 4.5005
R42820 VINP.n264 VINP.n139 4.5005
R42821 VINP.n304 VINP.n139 4.5005
R42822 VINP.n263 VINP.n139 4.5005
R42823 VINP.n306 VINP.n139 4.5005
R42824 VINP.n262 VINP.n139 4.5005
R42825 VINP.n308 VINP.n139 4.5005
R42826 VINP.n261 VINP.n139 4.5005
R42827 VINP.n310 VINP.n139 4.5005
R42828 VINP.n260 VINP.n139 4.5005
R42829 VINP.n312 VINP.n139 4.5005
R42830 VINP.n259 VINP.n139 4.5005
R42831 VINP.n314 VINP.n139 4.5005
R42832 VINP.n258 VINP.n139 4.5005
R42833 VINP.n316 VINP.n139 4.5005
R42834 VINP.n257 VINP.n139 4.5005
R42835 VINP.n318 VINP.n139 4.5005
R42836 VINP.n256 VINP.n139 4.5005
R42837 VINP.n320 VINP.n139 4.5005
R42838 VINP.n255 VINP.n139 4.5005
R42839 VINP.n322 VINP.n139 4.5005
R42840 VINP.n254 VINP.n139 4.5005
R42841 VINP.n324 VINP.n139 4.5005
R42842 VINP.n253 VINP.n139 4.5005
R42843 VINP.n326 VINP.n139 4.5005
R42844 VINP.n252 VINP.n139 4.5005
R42845 VINP.n328 VINP.n139 4.5005
R42846 VINP.n251 VINP.n139 4.5005
R42847 VINP.n330 VINP.n139 4.5005
R42848 VINP.n250 VINP.n139 4.5005
R42849 VINP.n332 VINP.n139 4.5005
R42850 VINP.n249 VINP.n139 4.5005
R42851 VINP.n334 VINP.n139 4.5005
R42852 VINP.n248 VINP.n139 4.5005
R42853 VINP.n336 VINP.n139 4.5005
R42854 VINP.n247 VINP.n139 4.5005
R42855 VINP.n338 VINP.n139 4.5005
R42856 VINP.n246 VINP.n139 4.5005
R42857 VINP.n340 VINP.n139 4.5005
R42858 VINP.n245 VINP.n139 4.5005
R42859 VINP.n342 VINP.n139 4.5005
R42860 VINP.n244 VINP.n139 4.5005
R42861 VINP.n344 VINP.n139 4.5005
R42862 VINP.n243 VINP.n139 4.5005
R42863 VINP.n346 VINP.n139 4.5005
R42864 VINP.n242 VINP.n139 4.5005
R42865 VINP.n348 VINP.n139 4.5005
R42866 VINP.n241 VINP.n139 4.5005
R42867 VINP.n350 VINP.n139 4.5005
R42868 VINP.n240 VINP.n139 4.5005
R42869 VINP.n352 VINP.n139 4.5005
R42870 VINP.n239 VINP.n139 4.5005
R42871 VINP.n354 VINP.n139 4.5005
R42872 VINP.n238 VINP.n139 4.5005
R42873 VINP.n356 VINP.n139 4.5005
R42874 VINP.n237 VINP.n139 4.5005
R42875 VINP.n358 VINP.n139 4.5005
R42876 VINP.n236 VINP.n139 4.5005
R42877 VINP.n360 VINP.n139 4.5005
R42878 VINP.n235 VINP.n139 4.5005
R42879 VINP.n362 VINP.n139 4.5005
R42880 VINP.n234 VINP.n139 4.5005
R42881 VINP.n364 VINP.n139 4.5005
R42882 VINP.n233 VINP.n139 4.5005
R42883 VINP.n366 VINP.n139 4.5005
R42884 VINP.n232 VINP.n139 4.5005
R42885 VINP.n368 VINP.n139 4.5005
R42886 VINP.n231 VINP.n139 4.5005
R42887 VINP.n370 VINP.n139 4.5005
R42888 VINP.n230 VINP.n139 4.5005
R42889 VINP.n372 VINP.n139 4.5005
R42890 VINP.n229 VINP.n139 4.5005
R42891 VINP.n374 VINP.n139 4.5005
R42892 VINP.n228 VINP.n139 4.5005
R42893 VINP.n376 VINP.n139 4.5005
R42894 VINP.n227 VINP.n139 4.5005
R42895 VINP.n378 VINP.n139 4.5005
R42896 VINP.n226 VINP.n139 4.5005
R42897 VINP.n380 VINP.n139 4.5005
R42898 VINP.n225 VINP.n139 4.5005
R42899 VINP.n382 VINP.n139 4.5005
R42900 VINP.n224 VINP.n139 4.5005
R42901 VINP.n384 VINP.n139 4.5005
R42902 VINP.n223 VINP.n139 4.5005
R42903 VINP.n386 VINP.n139 4.5005
R42904 VINP.n222 VINP.n139 4.5005
R42905 VINP.n388 VINP.n139 4.5005
R42906 VINP.n221 VINP.n139 4.5005
R42907 VINP.n390 VINP.n139 4.5005
R42908 VINP.n220 VINP.n139 4.5005
R42909 VINP.n392 VINP.n139 4.5005
R42910 VINP.n219 VINP.n139 4.5005
R42911 VINP.n394 VINP.n139 4.5005
R42912 VINP.n218 VINP.n139 4.5005
R42913 VINP.n396 VINP.n139 4.5005
R42914 VINP.n217 VINP.n139 4.5005
R42915 VINP.n398 VINP.n139 4.5005
R42916 VINP.n216 VINP.n139 4.5005
R42917 VINP.n400 VINP.n139 4.5005
R42918 VINP.n215 VINP.n139 4.5005
R42919 VINP.n654 VINP.n139 4.5005
R42920 VINP.n656 VINP.n139 4.5005
R42921 VINP.n139 VINP.n0 4.5005
R42922 VINP.n278 VINP.n162 4.5005
R42923 VINP.n276 VINP.n162 4.5005
R42924 VINP.n280 VINP.n162 4.5005
R42925 VINP.n275 VINP.n162 4.5005
R42926 VINP.n282 VINP.n162 4.5005
R42927 VINP.n274 VINP.n162 4.5005
R42928 VINP.n284 VINP.n162 4.5005
R42929 VINP.n273 VINP.n162 4.5005
R42930 VINP.n286 VINP.n162 4.5005
R42931 VINP.n272 VINP.n162 4.5005
R42932 VINP.n288 VINP.n162 4.5005
R42933 VINP.n271 VINP.n162 4.5005
R42934 VINP.n290 VINP.n162 4.5005
R42935 VINP.n270 VINP.n162 4.5005
R42936 VINP.n292 VINP.n162 4.5005
R42937 VINP.n269 VINP.n162 4.5005
R42938 VINP.n294 VINP.n162 4.5005
R42939 VINP.n268 VINP.n162 4.5005
R42940 VINP.n296 VINP.n162 4.5005
R42941 VINP.n267 VINP.n162 4.5005
R42942 VINP.n298 VINP.n162 4.5005
R42943 VINP.n266 VINP.n162 4.5005
R42944 VINP.n300 VINP.n162 4.5005
R42945 VINP.n265 VINP.n162 4.5005
R42946 VINP.n302 VINP.n162 4.5005
R42947 VINP.n264 VINP.n162 4.5005
R42948 VINP.n304 VINP.n162 4.5005
R42949 VINP.n263 VINP.n162 4.5005
R42950 VINP.n306 VINP.n162 4.5005
R42951 VINP.n262 VINP.n162 4.5005
R42952 VINP.n308 VINP.n162 4.5005
R42953 VINP.n261 VINP.n162 4.5005
R42954 VINP.n310 VINP.n162 4.5005
R42955 VINP.n260 VINP.n162 4.5005
R42956 VINP.n312 VINP.n162 4.5005
R42957 VINP.n259 VINP.n162 4.5005
R42958 VINP.n314 VINP.n162 4.5005
R42959 VINP.n258 VINP.n162 4.5005
R42960 VINP.n316 VINP.n162 4.5005
R42961 VINP.n257 VINP.n162 4.5005
R42962 VINP.n318 VINP.n162 4.5005
R42963 VINP.n256 VINP.n162 4.5005
R42964 VINP.n320 VINP.n162 4.5005
R42965 VINP.n255 VINP.n162 4.5005
R42966 VINP.n322 VINP.n162 4.5005
R42967 VINP.n254 VINP.n162 4.5005
R42968 VINP.n324 VINP.n162 4.5005
R42969 VINP.n253 VINP.n162 4.5005
R42970 VINP.n326 VINP.n162 4.5005
R42971 VINP.n252 VINP.n162 4.5005
R42972 VINP.n328 VINP.n162 4.5005
R42973 VINP.n251 VINP.n162 4.5005
R42974 VINP.n330 VINP.n162 4.5005
R42975 VINP.n250 VINP.n162 4.5005
R42976 VINP.n332 VINP.n162 4.5005
R42977 VINP.n249 VINP.n162 4.5005
R42978 VINP.n334 VINP.n162 4.5005
R42979 VINP.n248 VINP.n162 4.5005
R42980 VINP.n336 VINP.n162 4.5005
R42981 VINP.n247 VINP.n162 4.5005
R42982 VINP.n338 VINP.n162 4.5005
R42983 VINP.n246 VINP.n162 4.5005
R42984 VINP.n340 VINP.n162 4.5005
R42985 VINP.n245 VINP.n162 4.5005
R42986 VINP.n342 VINP.n162 4.5005
R42987 VINP.n244 VINP.n162 4.5005
R42988 VINP.n344 VINP.n162 4.5005
R42989 VINP.n243 VINP.n162 4.5005
R42990 VINP.n346 VINP.n162 4.5005
R42991 VINP.n242 VINP.n162 4.5005
R42992 VINP.n348 VINP.n162 4.5005
R42993 VINP.n241 VINP.n162 4.5005
R42994 VINP.n350 VINP.n162 4.5005
R42995 VINP.n240 VINP.n162 4.5005
R42996 VINP.n352 VINP.n162 4.5005
R42997 VINP.n239 VINP.n162 4.5005
R42998 VINP.n354 VINP.n162 4.5005
R42999 VINP.n238 VINP.n162 4.5005
R43000 VINP.n356 VINP.n162 4.5005
R43001 VINP.n237 VINP.n162 4.5005
R43002 VINP.n358 VINP.n162 4.5005
R43003 VINP.n236 VINP.n162 4.5005
R43004 VINP.n360 VINP.n162 4.5005
R43005 VINP.n235 VINP.n162 4.5005
R43006 VINP.n362 VINP.n162 4.5005
R43007 VINP.n234 VINP.n162 4.5005
R43008 VINP.n364 VINP.n162 4.5005
R43009 VINP.n233 VINP.n162 4.5005
R43010 VINP.n366 VINP.n162 4.5005
R43011 VINP.n232 VINP.n162 4.5005
R43012 VINP.n368 VINP.n162 4.5005
R43013 VINP.n231 VINP.n162 4.5005
R43014 VINP.n370 VINP.n162 4.5005
R43015 VINP.n230 VINP.n162 4.5005
R43016 VINP.n372 VINP.n162 4.5005
R43017 VINP.n229 VINP.n162 4.5005
R43018 VINP.n374 VINP.n162 4.5005
R43019 VINP.n228 VINP.n162 4.5005
R43020 VINP.n376 VINP.n162 4.5005
R43021 VINP.n227 VINP.n162 4.5005
R43022 VINP.n378 VINP.n162 4.5005
R43023 VINP.n226 VINP.n162 4.5005
R43024 VINP.n380 VINP.n162 4.5005
R43025 VINP.n225 VINP.n162 4.5005
R43026 VINP.n382 VINP.n162 4.5005
R43027 VINP.n224 VINP.n162 4.5005
R43028 VINP.n384 VINP.n162 4.5005
R43029 VINP.n223 VINP.n162 4.5005
R43030 VINP.n386 VINP.n162 4.5005
R43031 VINP.n222 VINP.n162 4.5005
R43032 VINP.n388 VINP.n162 4.5005
R43033 VINP.n221 VINP.n162 4.5005
R43034 VINP.n390 VINP.n162 4.5005
R43035 VINP.n220 VINP.n162 4.5005
R43036 VINP.n392 VINP.n162 4.5005
R43037 VINP.n219 VINP.n162 4.5005
R43038 VINP.n394 VINP.n162 4.5005
R43039 VINP.n218 VINP.n162 4.5005
R43040 VINP.n396 VINP.n162 4.5005
R43041 VINP.n217 VINP.n162 4.5005
R43042 VINP.n398 VINP.n162 4.5005
R43043 VINP.n216 VINP.n162 4.5005
R43044 VINP.n400 VINP.n162 4.5005
R43045 VINP.n215 VINP.n162 4.5005
R43046 VINP.n654 VINP.n162 4.5005
R43047 VINP.n656 VINP.n162 4.5005
R43048 VINP.n162 VINP.n0 4.5005
R43049 VINP.n278 VINP.n138 4.5005
R43050 VINP.n276 VINP.n138 4.5005
R43051 VINP.n280 VINP.n138 4.5005
R43052 VINP.n275 VINP.n138 4.5005
R43053 VINP.n282 VINP.n138 4.5005
R43054 VINP.n274 VINP.n138 4.5005
R43055 VINP.n284 VINP.n138 4.5005
R43056 VINP.n273 VINP.n138 4.5005
R43057 VINP.n286 VINP.n138 4.5005
R43058 VINP.n272 VINP.n138 4.5005
R43059 VINP.n288 VINP.n138 4.5005
R43060 VINP.n271 VINP.n138 4.5005
R43061 VINP.n290 VINP.n138 4.5005
R43062 VINP.n270 VINP.n138 4.5005
R43063 VINP.n292 VINP.n138 4.5005
R43064 VINP.n269 VINP.n138 4.5005
R43065 VINP.n294 VINP.n138 4.5005
R43066 VINP.n268 VINP.n138 4.5005
R43067 VINP.n296 VINP.n138 4.5005
R43068 VINP.n267 VINP.n138 4.5005
R43069 VINP.n298 VINP.n138 4.5005
R43070 VINP.n266 VINP.n138 4.5005
R43071 VINP.n300 VINP.n138 4.5005
R43072 VINP.n265 VINP.n138 4.5005
R43073 VINP.n302 VINP.n138 4.5005
R43074 VINP.n264 VINP.n138 4.5005
R43075 VINP.n304 VINP.n138 4.5005
R43076 VINP.n263 VINP.n138 4.5005
R43077 VINP.n306 VINP.n138 4.5005
R43078 VINP.n262 VINP.n138 4.5005
R43079 VINP.n308 VINP.n138 4.5005
R43080 VINP.n261 VINP.n138 4.5005
R43081 VINP.n310 VINP.n138 4.5005
R43082 VINP.n260 VINP.n138 4.5005
R43083 VINP.n312 VINP.n138 4.5005
R43084 VINP.n259 VINP.n138 4.5005
R43085 VINP.n314 VINP.n138 4.5005
R43086 VINP.n258 VINP.n138 4.5005
R43087 VINP.n316 VINP.n138 4.5005
R43088 VINP.n257 VINP.n138 4.5005
R43089 VINP.n318 VINP.n138 4.5005
R43090 VINP.n256 VINP.n138 4.5005
R43091 VINP.n320 VINP.n138 4.5005
R43092 VINP.n255 VINP.n138 4.5005
R43093 VINP.n322 VINP.n138 4.5005
R43094 VINP.n254 VINP.n138 4.5005
R43095 VINP.n324 VINP.n138 4.5005
R43096 VINP.n253 VINP.n138 4.5005
R43097 VINP.n326 VINP.n138 4.5005
R43098 VINP.n252 VINP.n138 4.5005
R43099 VINP.n328 VINP.n138 4.5005
R43100 VINP.n251 VINP.n138 4.5005
R43101 VINP.n330 VINP.n138 4.5005
R43102 VINP.n250 VINP.n138 4.5005
R43103 VINP.n332 VINP.n138 4.5005
R43104 VINP.n249 VINP.n138 4.5005
R43105 VINP.n334 VINP.n138 4.5005
R43106 VINP.n248 VINP.n138 4.5005
R43107 VINP.n336 VINP.n138 4.5005
R43108 VINP.n247 VINP.n138 4.5005
R43109 VINP.n338 VINP.n138 4.5005
R43110 VINP.n246 VINP.n138 4.5005
R43111 VINP.n340 VINP.n138 4.5005
R43112 VINP.n245 VINP.n138 4.5005
R43113 VINP.n342 VINP.n138 4.5005
R43114 VINP.n244 VINP.n138 4.5005
R43115 VINP.n344 VINP.n138 4.5005
R43116 VINP.n243 VINP.n138 4.5005
R43117 VINP.n346 VINP.n138 4.5005
R43118 VINP.n242 VINP.n138 4.5005
R43119 VINP.n348 VINP.n138 4.5005
R43120 VINP.n241 VINP.n138 4.5005
R43121 VINP.n350 VINP.n138 4.5005
R43122 VINP.n240 VINP.n138 4.5005
R43123 VINP.n352 VINP.n138 4.5005
R43124 VINP.n239 VINP.n138 4.5005
R43125 VINP.n354 VINP.n138 4.5005
R43126 VINP.n238 VINP.n138 4.5005
R43127 VINP.n356 VINP.n138 4.5005
R43128 VINP.n237 VINP.n138 4.5005
R43129 VINP.n358 VINP.n138 4.5005
R43130 VINP.n236 VINP.n138 4.5005
R43131 VINP.n360 VINP.n138 4.5005
R43132 VINP.n235 VINP.n138 4.5005
R43133 VINP.n362 VINP.n138 4.5005
R43134 VINP.n234 VINP.n138 4.5005
R43135 VINP.n364 VINP.n138 4.5005
R43136 VINP.n233 VINP.n138 4.5005
R43137 VINP.n366 VINP.n138 4.5005
R43138 VINP.n232 VINP.n138 4.5005
R43139 VINP.n368 VINP.n138 4.5005
R43140 VINP.n231 VINP.n138 4.5005
R43141 VINP.n370 VINP.n138 4.5005
R43142 VINP.n230 VINP.n138 4.5005
R43143 VINP.n372 VINP.n138 4.5005
R43144 VINP.n229 VINP.n138 4.5005
R43145 VINP.n374 VINP.n138 4.5005
R43146 VINP.n228 VINP.n138 4.5005
R43147 VINP.n376 VINP.n138 4.5005
R43148 VINP.n227 VINP.n138 4.5005
R43149 VINP.n378 VINP.n138 4.5005
R43150 VINP.n226 VINP.n138 4.5005
R43151 VINP.n380 VINP.n138 4.5005
R43152 VINP.n225 VINP.n138 4.5005
R43153 VINP.n382 VINP.n138 4.5005
R43154 VINP.n224 VINP.n138 4.5005
R43155 VINP.n384 VINP.n138 4.5005
R43156 VINP.n223 VINP.n138 4.5005
R43157 VINP.n386 VINP.n138 4.5005
R43158 VINP.n222 VINP.n138 4.5005
R43159 VINP.n388 VINP.n138 4.5005
R43160 VINP.n221 VINP.n138 4.5005
R43161 VINP.n390 VINP.n138 4.5005
R43162 VINP.n220 VINP.n138 4.5005
R43163 VINP.n392 VINP.n138 4.5005
R43164 VINP.n219 VINP.n138 4.5005
R43165 VINP.n394 VINP.n138 4.5005
R43166 VINP.n218 VINP.n138 4.5005
R43167 VINP.n396 VINP.n138 4.5005
R43168 VINP.n217 VINP.n138 4.5005
R43169 VINP.n398 VINP.n138 4.5005
R43170 VINP.n216 VINP.n138 4.5005
R43171 VINP.n400 VINP.n138 4.5005
R43172 VINP.n215 VINP.n138 4.5005
R43173 VINP.n654 VINP.n138 4.5005
R43174 VINP.n656 VINP.n138 4.5005
R43175 VINP.n138 VINP.n0 4.5005
R43176 VINP.n278 VINP.n163 4.5005
R43177 VINP.n276 VINP.n163 4.5005
R43178 VINP.n280 VINP.n163 4.5005
R43179 VINP.n275 VINP.n163 4.5005
R43180 VINP.n282 VINP.n163 4.5005
R43181 VINP.n274 VINP.n163 4.5005
R43182 VINP.n284 VINP.n163 4.5005
R43183 VINP.n273 VINP.n163 4.5005
R43184 VINP.n286 VINP.n163 4.5005
R43185 VINP.n272 VINP.n163 4.5005
R43186 VINP.n288 VINP.n163 4.5005
R43187 VINP.n271 VINP.n163 4.5005
R43188 VINP.n290 VINP.n163 4.5005
R43189 VINP.n270 VINP.n163 4.5005
R43190 VINP.n292 VINP.n163 4.5005
R43191 VINP.n269 VINP.n163 4.5005
R43192 VINP.n294 VINP.n163 4.5005
R43193 VINP.n268 VINP.n163 4.5005
R43194 VINP.n296 VINP.n163 4.5005
R43195 VINP.n267 VINP.n163 4.5005
R43196 VINP.n298 VINP.n163 4.5005
R43197 VINP.n266 VINP.n163 4.5005
R43198 VINP.n300 VINP.n163 4.5005
R43199 VINP.n265 VINP.n163 4.5005
R43200 VINP.n302 VINP.n163 4.5005
R43201 VINP.n264 VINP.n163 4.5005
R43202 VINP.n304 VINP.n163 4.5005
R43203 VINP.n263 VINP.n163 4.5005
R43204 VINP.n306 VINP.n163 4.5005
R43205 VINP.n262 VINP.n163 4.5005
R43206 VINP.n308 VINP.n163 4.5005
R43207 VINP.n261 VINP.n163 4.5005
R43208 VINP.n310 VINP.n163 4.5005
R43209 VINP.n260 VINP.n163 4.5005
R43210 VINP.n312 VINP.n163 4.5005
R43211 VINP.n259 VINP.n163 4.5005
R43212 VINP.n314 VINP.n163 4.5005
R43213 VINP.n258 VINP.n163 4.5005
R43214 VINP.n316 VINP.n163 4.5005
R43215 VINP.n257 VINP.n163 4.5005
R43216 VINP.n318 VINP.n163 4.5005
R43217 VINP.n256 VINP.n163 4.5005
R43218 VINP.n320 VINP.n163 4.5005
R43219 VINP.n255 VINP.n163 4.5005
R43220 VINP.n322 VINP.n163 4.5005
R43221 VINP.n254 VINP.n163 4.5005
R43222 VINP.n324 VINP.n163 4.5005
R43223 VINP.n253 VINP.n163 4.5005
R43224 VINP.n326 VINP.n163 4.5005
R43225 VINP.n252 VINP.n163 4.5005
R43226 VINP.n328 VINP.n163 4.5005
R43227 VINP.n251 VINP.n163 4.5005
R43228 VINP.n330 VINP.n163 4.5005
R43229 VINP.n250 VINP.n163 4.5005
R43230 VINP.n332 VINP.n163 4.5005
R43231 VINP.n249 VINP.n163 4.5005
R43232 VINP.n334 VINP.n163 4.5005
R43233 VINP.n248 VINP.n163 4.5005
R43234 VINP.n336 VINP.n163 4.5005
R43235 VINP.n247 VINP.n163 4.5005
R43236 VINP.n338 VINP.n163 4.5005
R43237 VINP.n246 VINP.n163 4.5005
R43238 VINP.n340 VINP.n163 4.5005
R43239 VINP.n245 VINP.n163 4.5005
R43240 VINP.n342 VINP.n163 4.5005
R43241 VINP.n244 VINP.n163 4.5005
R43242 VINP.n344 VINP.n163 4.5005
R43243 VINP.n243 VINP.n163 4.5005
R43244 VINP.n346 VINP.n163 4.5005
R43245 VINP.n242 VINP.n163 4.5005
R43246 VINP.n348 VINP.n163 4.5005
R43247 VINP.n241 VINP.n163 4.5005
R43248 VINP.n350 VINP.n163 4.5005
R43249 VINP.n240 VINP.n163 4.5005
R43250 VINP.n352 VINP.n163 4.5005
R43251 VINP.n239 VINP.n163 4.5005
R43252 VINP.n354 VINP.n163 4.5005
R43253 VINP.n238 VINP.n163 4.5005
R43254 VINP.n356 VINP.n163 4.5005
R43255 VINP.n237 VINP.n163 4.5005
R43256 VINP.n358 VINP.n163 4.5005
R43257 VINP.n236 VINP.n163 4.5005
R43258 VINP.n360 VINP.n163 4.5005
R43259 VINP.n235 VINP.n163 4.5005
R43260 VINP.n362 VINP.n163 4.5005
R43261 VINP.n234 VINP.n163 4.5005
R43262 VINP.n364 VINP.n163 4.5005
R43263 VINP.n233 VINP.n163 4.5005
R43264 VINP.n366 VINP.n163 4.5005
R43265 VINP.n232 VINP.n163 4.5005
R43266 VINP.n368 VINP.n163 4.5005
R43267 VINP.n231 VINP.n163 4.5005
R43268 VINP.n370 VINP.n163 4.5005
R43269 VINP.n230 VINP.n163 4.5005
R43270 VINP.n372 VINP.n163 4.5005
R43271 VINP.n229 VINP.n163 4.5005
R43272 VINP.n374 VINP.n163 4.5005
R43273 VINP.n228 VINP.n163 4.5005
R43274 VINP.n376 VINP.n163 4.5005
R43275 VINP.n227 VINP.n163 4.5005
R43276 VINP.n378 VINP.n163 4.5005
R43277 VINP.n226 VINP.n163 4.5005
R43278 VINP.n380 VINP.n163 4.5005
R43279 VINP.n225 VINP.n163 4.5005
R43280 VINP.n382 VINP.n163 4.5005
R43281 VINP.n224 VINP.n163 4.5005
R43282 VINP.n384 VINP.n163 4.5005
R43283 VINP.n223 VINP.n163 4.5005
R43284 VINP.n386 VINP.n163 4.5005
R43285 VINP.n222 VINP.n163 4.5005
R43286 VINP.n388 VINP.n163 4.5005
R43287 VINP.n221 VINP.n163 4.5005
R43288 VINP.n390 VINP.n163 4.5005
R43289 VINP.n220 VINP.n163 4.5005
R43290 VINP.n392 VINP.n163 4.5005
R43291 VINP.n219 VINP.n163 4.5005
R43292 VINP.n394 VINP.n163 4.5005
R43293 VINP.n218 VINP.n163 4.5005
R43294 VINP.n396 VINP.n163 4.5005
R43295 VINP.n217 VINP.n163 4.5005
R43296 VINP.n398 VINP.n163 4.5005
R43297 VINP.n216 VINP.n163 4.5005
R43298 VINP.n400 VINP.n163 4.5005
R43299 VINP.n215 VINP.n163 4.5005
R43300 VINP.n654 VINP.n163 4.5005
R43301 VINP.n656 VINP.n163 4.5005
R43302 VINP.n163 VINP.n0 4.5005
R43303 VINP.n278 VINP.n137 4.5005
R43304 VINP.n276 VINP.n137 4.5005
R43305 VINP.n280 VINP.n137 4.5005
R43306 VINP.n275 VINP.n137 4.5005
R43307 VINP.n282 VINP.n137 4.5005
R43308 VINP.n274 VINP.n137 4.5005
R43309 VINP.n284 VINP.n137 4.5005
R43310 VINP.n273 VINP.n137 4.5005
R43311 VINP.n286 VINP.n137 4.5005
R43312 VINP.n272 VINP.n137 4.5005
R43313 VINP.n288 VINP.n137 4.5005
R43314 VINP.n271 VINP.n137 4.5005
R43315 VINP.n290 VINP.n137 4.5005
R43316 VINP.n270 VINP.n137 4.5005
R43317 VINP.n292 VINP.n137 4.5005
R43318 VINP.n269 VINP.n137 4.5005
R43319 VINP.n294 VINP.n137 4.5005
R43320 VINP.n268 VINP.n137 4.5005
R43321 VINP.n296 VINP.n137 4.5005
R43322 VINP.n267 VINP.n137 4.5005
R43323 VINP.n298 VINP.n137 4.5005
R43324 VINP.n266 VINP.n137 4.5005
R43325 VINP.n300 VINP.n137 4.5005
R43326 VINP.n265 VINP.n137 4.5005
R43327 VINP.n302 VINP.n137 4.5005
R43328 VINP.n264 VINP.n137 4.5005
R43329 VINP.n304 VINP.n137 4.5005
R43330 VINP.n263 VINP.n137 4.5005
R43331 VINP.n306 VINP.n137 4.5005
R43332 VINP.n262 VINP.n137 4.5005
R43333 VINP.n308 VINP.n137 4.5005
R43334 VINP.n261 VINP.n137 4.5005
R43335 VINP.n310 VINP.n137 4.5005
R43336 VINP.n260 VINP.n137 4.5005
R43337 VINP.n312 VINP.n137 4.5005
R43338 VINP.n259 VINP.n137 4.5005
R43339 VINP.n314 VINP.n137 4.5005
R43340 VINP.n258 VINP.n137 4.5005
R43341 VINP.n316 VINP.n137 4.5005
R43342 VINP.n257 VINP.n137 4.5005
R43343 VINP.n318 VINP.n137 4.5005
R43344 VINP.n256 VINP.n137 4.5005
R43345 VINP.n320 VINP.n137 4.5005
R43346 VINP.n255 VINP.n137 4.5005
R43347 VINP.n322 VINP.n137 4.5005
R43348 VINP.n254 VINP.n137 4.5005
R43349 VINP.n324 VINP.n137 4.5005
R43350 VINP.n253 VINP.n137 4.5005
R43351 VINP.n326 VINP.n137 4.5005
R43352 VINP.n252 VINP.n137 4.5005
R43353 VINP.n328 VINP.n137 4.5005
R43354 VINP.n251 VINP.n137 4.5005
R43355 VINP.n330 VINP.n137 4.5005
R43356 VINP.n250 VINP.n137 4.5005
R43357 VINP.n332 VINP.n137 4.5005
R43358 VINP.n249 VINP.n137 4.5005
R43359 VINP.n334 VINP.n137 4.5005
R43360 VINP.n248 VINP.n137 4.5005
R43361 VINP.n336 VINP.n137 4.5005
R43362 VINP.n247 VINP.n137 4.5005
R43363 VINP.n338 VINP.n137 4.5005
R43364 VINP.n246 VINP.n137 4.5005
R43365 VINP.n340 VINP.n137 4.5005
R43366 VINP.n245 VINP.n137 4.5005
R43367 VINP.n342 VINP.n137 4.5005
R43368 VINP.n244 VINP.n137 4.5005
R43369 VINP.n344 VINP.n137 4.5005
R43370 VINP.n243 VINP.n137 4.5005
R43371 VINP.n346 VINP.n137 4.5005
R43372 VINP.n242 VINP.n137 4.5005
R43373 VINP.n348 VINP.n137 4.5005
R43374 VINP.n241 VINP.n137 4.5005
R43375 VINP.n350 VINP.n137 4.5005
R43376 VINP.n240 VINP.n137 4.5005
R43377 VINP.n352 VINP.n137 4.5005
R43378 VINP.n239 VINP.n137 4.5005
R43379 VINP.n354 VINP.n137 4.5005
R43380 VINP.n238 VINP.n137 4.5005
R43381 VINP.n356 VINP.n137 4.5005
R43382 VINP.n237 VINP.n137 4.5005
R43383 VINP.n358 VINP.n137 4.5005
R43384 VINP.n236 VINP.n137 4.5005
R43385 VINP.n360 VINP.n137 4.5005
R43386 VINP.n235 VINP.n137 4.5005
R43387 VINP.n362 VINP.n137 4.5005
R43388 VINP.n234 VINP.n137 4.5005
R43389 VINP.n364 VINP.n137 4.5005
R43390 VINP.n233 VINP.n137 4.5005
R43391 VINP.n366 VINP.n137 4.5005
R43392 VINP.n232 VINP.n137 4.5005
R43393 VINP.n368 VINP.n137 4.5005
R43394 VINP.n231 VINP.n137 4.5005
R43395 VINP.n370 VINP.n137 4.5005
R43396 VINP.n230 VINP.n137 4.5005
R43397 VINP.n372 VINP.n137 4.5005
R43398 VINP.n229 VINP.n137 4.5005
R43399 VINP.n374 VINP.n137 4.5005
R43400 VINP.n228 VINP.n137 4.5005
R43401 VINP.n376 VINP.n137 4.5005
R43402 VINP.n227 VINP.n137 4.5005
R43403 VINP.n378 VINP.n137 4.5005
R43404 VINP.n226 VINP.n137 4.5005
R43405 VINP.n380 VINP.n137 4.5005
R43406 VINP.n225 VINP.n137 4.5005
R43407 VINP.n382 VINP.n137 4.5005
R43408 VINP.n224 VINP.n137 4.5005
R43409 VINP.n384 VINP.n137 4.5005
R43410 VINP.n223 VINP.n137 4.5005
R43411 VINP.n386 VINP.n137 4.5005
R43412 VINP.n222 VINP.n137 4.5005
R43413 VINP.n388 VINP.n137 4.5005
R43414 VINP.n221 VINP.n137 4.5005
R43415 VINP.n390 VINP.n137 4.5005
R43416 VINP.n220 VINP.n137 4.5005
R43417 VINP.n392 VINP.n137 4.5005
R43418 VINP.n219 VINP.n137 4.5005
R43419 VINP.n394 VINP.n137 4.5005
R43420 VINP.n218 VINP.n137 4.5005
R43421 VINP.n396 VINP.n137 4.5005
R43422 VINP.n217 VINP.n137 4.5005
R43423 VINP.n398 VINP.n137 4.5005
R43424 VINP.n216 VINP.n137 4.5005
R43425 VINP.n400 VINP.n137 4.5005
R43426 VINP.n215 VINP.n137 4.5005
R43427 VINP.n654 VINP.n137 4.5005
R43428 VINP.n656 VINP.n137 4.5005
R43429 VINP.n137 VINP.n0 4.5005
R43430 VINP.n278 VINP.n164 4.5005
R43431 VINP.n276 VINP.n164 4.5005
R43432 VINP.n280 VINP.n164 4.5005
R43433 VINP.n275 VINP.n164 4.5005
R43434 VINP.n282 VINP.n164 4.5005
R43435 VINP.n274 VINP.n164 4.5005
R43436 VINP.n284 VINP.n164 4.5005
R43437 VINP.n273 VINP.n164 4.5005
R43438 VINP.n286 VINP.n164 4.5005
R43439 VINP.n272 VINP.n164 4.5005
R43440 VINP.n288 VINP.n164 4.5005
R43441 VINP.n271 VINP.n164 4.5005
R43442 VINP.n290 VINP.n164 4.5005
R43443 VINP.n270 VINP.n164 4.5005
R43444 VINP.n292 VINP.n164 4.5005
R43445 VINP.n269 VINP.n164 4.5005
R43446 VINP.n294 VINP.n164 4.5005
R43447 VINP.n268 VINP.n164 4.5005
R43448 VINP.n296 VINP.n164 4.5005
R43449 VINP.n267 VINP.n164 4.5005
R43450 VINP.n298 VINP.n164 4.5005
R43451 VINP.n266 VINP.n164 4.5005
R43452 VINP.n300 VINP.n164 4.5005
R43453 VINP.n265 VINP.n164 4.5005
R43454 VINP.n302 VINP.n164 4.5005
R43455 VINP.n264 VINP.n164 4.5005
R43456 VINP.n304 VINP.n164 4.5005
R43457 VINP.n263 VINP.n164 4.5005
R43458 VINP.n306 VINP.n164 4.5005
R43459 VINP.n262 VINP.n164 4.5005
R43460 VINP.n308 VINP.n164 4.5005
R43461 VINP.n261 VINP.n164 4.5005
R43462 VINP.n310 VINP.n164 4.5005
R43463 VINP.n260 VINP.n164 4.5005
R43464 VINP.n312 VINP.n164 4.5005
R43465 VINP.n259 VINP.n164 4.5005
R43466 VINP.n314 VINP.n164 4.5005
R43467 VINP.n258 VINP.n164 4.5005
R43468 VINP.n316 VINP.n164 4.5005
R43469 VINP.n257 VINP.n164 4.5005
R43470 VINP.n318 VINP.n164 4.5005
R43471 VINP.n256 VINP.n164 4.5005
R43472 VINP.n320 VINP.n164 4.5005
R43473 VINP.n255 VINP.n164 4.5005
R43474 VINP.n322 VINP.n164 4.5005
R43475 VINP.n254 VINP.n164 4.5005
R43476 VINP.n324 VINP.n164 4.5005
R43477 VINP.n253 VINP.n164 4.5005
R43478 VINP.n326 VINP.n164 4.5005
R43479 VINP.n252 VINP.n164 4.5005
R43480 VINP.n328 VINP.n164 4.5005
R43481 VINP.n251 VINP.n164 4.5005
R43482 VINP.n330 VINP.n164 4.5005
R43483 VINP.n250 VINP.n164 4.5005
R43484 VINP.n332 VINP.n164 4.5005
R43485 VINP.n249 VINP.n164 4.5005
R43486 VINP.n334 VINP.n164 4.5005
R43487 VINP.n248 VINP.n164 4.5005
R43488 VINP.n336 VINP.n164 4.5005
R43489 VINP.n247 VINP.n164 4.5005
R43490 VINP.n338 VINP.n164 4.5005
R43491 VINP.n246 VINP.n164 4.5005
R43492 VINP.n340 VINP.n164 4.5005
R43493 VINP.n245 VINP.n164 4.5005
R43494 VINP.n342 VINP.n164 4.5005
R43495 VINP.n244 VINP.n164 4.5005
R43496 VINP.n344 VINP.n164 4.5005
R43497 VINP.n243 VINP.n164 4.5005
R43498 VINP.n346 VINP.n164 4.5005
R43499 VINP.n242 VINP.n164 4.5005
R43500 VINP.n348 VINP.n164 4.5005
R43501 VINP.n241 VINP.n164 4.5005
R43502 VINP.n350 VINP.n164 4.5005
R43503 VINP.n240 VINP.n164 4.5005
R43504 VINP.n352 VINP.n164 4.5005
R43505 VINP.n239 VINP.n164 4.5005
R43506 VINP.n354 VINP.n164 4.5005
R43507 VINP.n238 VINP.n164 4.5005
R43508 VINP.n356 VINP.n164 4.5005
R43509 VINP.n237 VINP.n164 4.5005
R43510 VINP.n358 VINP.n164 4.5005
R43511 VINP.n236 VINP.n164 4.5005
R43512 VINP.n360 VINP.n164 4.5005
R43513 VINP.n235 VINP.n164 4.5005
R43514 VINP.n362 VINP.n164 4.5005
R43515 VINP.n234 VINP.n164 4.5005
R43516 VINP.n364 VINP.n164 4.5005
R43517 VINP.n233 VINP.n164 4.5005
R43518 VINP.n366 VINP.n164 4.5005
R43519 VINP.n232 VINP.n164 4.5005
R43520 VINP.n368 VINP.n164 4.5005
R43521 VINP.n231 VINP.n164 4.5005
R43522 VINP.n370 VINP.n164 4.5005
R43523 VINP.n230 VINP.n164 4.5005
R43524 VINP.n372 VINP.n164 4.5005
R43525 VINP.n229 VINP.n164 4.5005
R43526 VINP.n374 VINP.n164 4.5005
R43527 VINP.n228 VINP.n164 4.5005
R43528 VINP.n376 VINP.n164 4.5005
R43529 VINP.n227 VINP.n164 4.5005
R43530 VINP.n378 VINP.n164 4.5005
R43531 VINP.n226 VINP.n164 4.5005
R43532 VINP.n380 VINP.n164 4.5005
R43533 VINP.n225 VINP.n164 4.5005
R43534 VINP.n382 VINP.n164 4.5005
R43535 VINP.n224 VINP.n164 4.5005
R43536 VINP.n384 VINP.n164 4.5005
R43537 VINP.n223 VINP.n164 4.5005
R43538 VINP.n386 VINP.n164 4.5005
R43539 VINP.n222 VINP.n164 4.5005
R43540 VINP.n388 VINP.n164 4.5005
R43541 VINP.n221 VINP.n164 4.5005
R43542 VINP.n390 VINP.n164 4.5005
R43543 VINP.n220 VINP.n164 4.5005
R43544 VINP.n392 VINP.n164 4.5005
R43545 VINP.n219 VINP.n164 4.5005
R43546 VINP.n394 VINP.n164 4.5005
R43547 VINP.n218 VINP.n164 4.5005
R43548 VINP.n396 VINP.n164 4.5005
R43549 VINP.n217 VINP.n164 4.5005
R43550 VINP.n398 VINP.n164 4.5005
R43551 VINP.n216 VINP.n164 4.5005
R43552 VINP.n400 VINP.n164 4.5005
R43553 VINP.n215 VINP.n164 4.5005
R43554 VINP.n654 VINP.n164 4.5005
R43555 VINP.n656 VINP.n164 4.5005
R43556 VINP.n164 VINP.n0 4.5005
R43557 VINP.n278 VINP.n136 4.5005
R43558 VINP.n276 VINP.n136 4.5005
R43559 VINP.n280 VINP.n136 4.5005
R43560 VINP.n275 VINP.n136 4.5005
R43561 VINP.n282 VINP.n136 4.5005
R43562 VINP.n274 VINP.n136 4.5005
R43563 VINP.n284 VINP.n136 4.5005
R43564 VINP.n273 VINP.n136 4.5005
R43565 VINP.n286 VINP.n136 4.5005
R43566 VINP.n272 VINP.n136 4.5005
R43567 VINP.n288 VINP.n136 4.5005
R43568 VINP.n271 VINP.n136 4.5005
R43569 VINP.n290 VINP.n136 4.5005
R43570 VINP.n270 VINP.n136 4.5005
R43571 VINP.n292 VINP.n136 4.5005
R43572 VINP.n269 VINP.n136 4.5005
R43573 VINP.n294 VINP.n136 4.5005
R43574 VINP.n268 VINP.n136 4.5005
R43575 VINP.n296 VINP.n136 4.5005
R43576 VINP.n267 VINP.n136 4.5005
R43577 VINP.n298 VINP.n136 4.5005
R43578 VINP.n266 VINP.n136 4.5005
R43579 VINP.n300 VINP.n136 4.5005
R43580 VINP.n265 VINP.n136 4.5005
R43581 VINP.n302 VINP.n136 4.5005
R43582 VINP.n264 VINP.n136 4.5005
R43583 VINP.n304 VINP.n136 4.5005
R43584 VINP.n263 VINP.n136 4.5005
R43585 VINP.n306 VINP.n136 4.5005
R43586 VINP.n262 VINP.n136 4.5005
R43587 VINP.n308 VINP.n136 4.5005
R43588 VINP.n261 VINP.n136 4.5005
R43589 VINP.n310 VINP.n136 4.5005
R43590 VINP.n260 VINP.n136 4.5005
R43591 VINP.n312 VINP.n136 4.5005
R43592 VINP.n259 VINP.n136 4.5005
R43593 VINP.n314 VINP.n136 4.5005
R43594 VINP.n258 VINP.n136 4.5005
R43595 VINP.n316 VINP.n136 4.5005
R43596 VINP.n257 VINP.n136 4.5005
R43597 VINP.n318 VINP.n136 4.5005
R43598 VINP.n256 VINP.n136 4.5005
R43599 VINP.n320 VINP.n136 4.5005
R43600 VINP.n255 VINP.n136 4.5005
R43601 VINP.n322 VINP.n136 4.5005
R43602 VINP.n254 VINP.n136 4.5005
R43603 VINP.n324 VINP.n136 4.5005
R43604 VINP.n253 VINP.n136 4.5005
R43605 VINP.n326 VINP.n136 4.5005
R43606 VINP.n252 VINP.n136 4.5005
R43607 VINP.n328 VINP.n136 4.5005
R43608 VINP.n251 VINP.n136 4.5005
R43609 VINP.n330 VINP.n136 4.5005
R43610 VINP.n250 VINP.n136 4.5005
R43611 VINP.n332 VINP.n136 4.5005
R43612 VINP.n249 VINP.n136 4.5005
R43613 VINP.n334 VINP.n136 4.5005
R43614 VINP.n248 VINP.n136 4.5005
R43615 VINP.n336 VINP.n136 4.5005
R43616 VINP.n247 VINP.n136 4.5005
R43617 VINP.n338 VINP.n136 4.5005
R43618 VINP.n246 VINP.n136 4.5005
R43619 VINP.n340 VINP.n136 4.5005
R43620 VINP.n245 VINP.n136 4.5005
R43621 VINP.n342 VINP.n136 4.5005
R43622 VINP.n244 VINP.n136 4.5005
R43623 VINP.n344 VINP.n136 4.5005
R43624 VINP.n243 VINP.n136 4.5005
R43625 VINP.n346 VINP.n136 4.5005
R43626 VINP.n242 VINP.n136 4.5005
R43627 VINP.n348 VINP.n136 4.5005
R43628 VINP.n241 VINP.n136 4.5005
R43629 VINP.n350 VINP.n136 4.5005
R43630 VINP.n240 VINP.n136 4.5005
R43631 VINP.n352 VINP.n136 4.5005
R43632 VINP.n239 VINP.n136 4.5005
R43633 VINP.n354 VINP.n136 4.5005
R43634 VINP.n238 VINP.n136 4.5005
R43635 VINP.n356 VINP.n136 4.5005
R43636 VINP.n237 VINP.n136 4.5005
R43637 VINP.n358 VINP.n136 4.5005
R43638 VINP.n236 VINP.n136 4.5005
R43639 VINP.n360 VINP.n136 4.5005
R43640 VINP.n235 VINP.n136 4.5005
R43641 VINP.n362 VINP.n136 4.5005
R43642 VINP.n234 VINP.n136 4.5005
R43643 VINP.n364 VINP.n136 4.5005
R43644 VINP.n233 VINP.n136 4.5005
R43645 VINP.n366 VINP.n136 4.5005
R43646 VINP.n232 VINP.n136 4.5005
R43647 VINP.n368 VINP.n136 4.5005
R43648 VINP.n231 VINP.n136 4.5005
R43649 VINP.n370 VINP.n136 4.5005
R43650 VINP.n230 VINP.n136 4.5005
R43651 VINP.n372 VINP.n136 4.5005
R43652 VINP.n229 VINP.n136 4.5005
R43653 VINP.n374 VINP.n136 4.5005
R43654 VINP.n228 VINP.n136 4.5005
R43655 VINP.n376 VINP.n136 4.5005
R43656 VINP.n227 VINP.n136 4.5005
R43657 VINP.n378 VINP.n136 4.5005
R43658 VINP.n226 VINP.n136 4.5005
R43659 VINP.n380 VINP.n136 4.5005
R43660 VINP.n225 VINP.n136 4.5005
R43661 VINP.n382 VINP.n136 4.5005
R43662 VINP.n224 VINP.n136 4.5005
R43663 VINP.n384 VINP.n136 4.5005
R43664 VINP.n223 VINP.n136 4.5005
R43665 VINP.n386 VINP.n136 4.5005
R43666 VINP.n222 VINP.n136 4.5005
R43667 VINP.n388 VINP.n136 4.5005
R43668 VINP.n221 VINP.n136 4.5005
R43669 VINP.n390 VINP.n136 4.5005
R43670 VINP.n220 VINP.n136 4.5005
R43671 VINP.n392 VINP.n136 4.5005
R43672 VINP.n219 VINP.n136 4.5005
R43673 VINP.n394 VINP.n136 4.5005
R43674 VINP.n218 VINP.n136 4.5005
R43675 VINP.n396 VINP.n136 4.5005
R43676 VINP.n217 VINP.n136 4.5005
R43677 VINP.n398 VINP.n136 4.5005
R43678 VINP.n216 VINP.n136 4.5005
R43679 VINP.n400 VINP.n136 4.5005
R43680 VINP.n215 VINP.n136 4.5005
R43681 VINP.n654 VINP.n136 4.5005
R43682 VINP.n656 VINP.n136 4.5005
R43683 VINP.n136 VINP.n0 4.5005
R43684 VINP.n278 VINP.n165 4.5005
R43685 VINP.n276 VINP.n165 4.5005
R43686 VINP.n280 VINP.n165 4.5005
R43687 VINP.n275 VINP.n165 4.5005
R43688 VINP.n282 VINP.n165 4.5005
R43689 VINP.n274 VINP.n165 4.5005
R43690 VINP.n284 VINP.n165 4.5005
R43691 VINP.n273 VINP.n165 4.5005
R43692 VINP.n286 VINP.n165 4.5005
R43693 VINP.n272 VINP.n165 4.5005
R43694 VINP.n288 VINP.n165 4.5005
R43695 VINP.n271 VINP.n165 4.5005
R43696 VINP.n290 VINP.n165 4.5005
R43697 VINP.n270 VINP.n165 4.5005
R43698 VINP.n292 VINP.n165 4.5005
R43699 VINP.n269 VINP.n165 4.5005
R43700 VINP.n294 VINP.n165 4.5005
R43701 VINP.n268 VINP.n165 4.5005
R43702 VINP.n296 VINP.n165 4.5005
R43703 VINP.n267 VINP.n165 4.5005
R43704 VINP.n298 VINP.n165 4.5005
R43705 VINP.n266 VINP.n165 4.5005
R43706 VINP.n300 VINP.n165 4.5005
R43707 VINP.n265 VINP.n165 4.5005
R43708 VINP.n302 VINP.n165 4.5005
R43709 VINP.n264 VINP.n165 4.5005
R43710 VINP.n304 VINP.n165 4.5005
R43711 VINP.n263 VINP.n165 4.5005
R43712 VINP.n306 VINP.n165 4.5005
R43713 VINP.n262 VINP.n165 4.5005
R43714 VINP.n308 VINP.n165 4.5005
R43715 VINP.n261 VINP.n165 4.5005
R43716 VINP.n310 VINP.n165 4.5005
R43717 VINP.n260 VINP.n165 4.5005
R43718 VINP.n312 VINP.n165 4.5005
R43719 VINP.n259 VINP.n165 4.5005
R43720 VINP.n314 VINP.n165 4.5005
R43721 VINP.n258 VINP.n165 4.5005
R43722 VINP.n316 VINP.n165 4.5005
R43723 VINP.n257 VINP.n165 4.5005
R43724 VINP.n318 VINP.n165 4.5005
R43725 VINP.n256 VINP.n165 4.5005
R43726 VINP.n320 VINP.n165 4.5005
R43727 VINP.n255 VINP.n165 4.5005
R43728 VINP.n322 VINP.n165 4.5005
R43729 VINP.n254 VINP.n165 4.5005
R43730 VINP.n324 VINP.n165 4.5005
R43731 VINP.n253 VINP.n165 4.5005
R43732 VINP.n326 VINP.n165 4.5005
R43733 VINP.n252 VINP.n165 4.5005
R43734 VINP.n328 VINP.n165 4.5005
R43735 VINP.n251 VINP.n165 4.5005
R43736 VINP.n330 VINP.n165 4.5005
R43737 VINP.n250 VINP.n165 4.5005
R43738 VINP.n332 VINP.n165 4.5005
R43739 VINP.n249 VINP.n165 4.5005
R43740 VINP.n334 VINP.n165 4.5005
R43741 VINP.n248 VINP.n165 4.5005
R43742 VINP.n336 VINP.n165 4.5005
R43743 VINP.n247 VINP.n165 4.5005
R43744 VINP.n338 VINP.n165 4.5005
R43745 VINP.n246 VINP.n165 4.5005
R43746 VINP.n340 VINP.n165 4.5005
R43747 VINP.n245 VINP.n165 4.5005
R43748 VINP.n342 VINP.n165 4.5005
R43749 VINP.n244 VINP.n165 4.5005
R43750 VINP.n344 VINP.n165 4.5005
R43751 VINP.n243 VINP.n165 4.5005
R43752 VINP.n346 VINP.n165 4.5005
R43753 VINP.n242 VINP.n165 4.5005
R43754 VINP.n348 VINP.n165 4.5005
R43755 VINP.n241 VINP.n165 4.5005
R43756 VINP.n350 VINP.n165 4.5005
R43757 VINP.n240 VINP.n165 4.5005
R43758 VINP.n352 VINP.n165 4.5005
R43759 VINP.n239 VINP.n165 4.5005
R43760 VINP.n354 VINP.n165 4.5005
R43761 VINP.n238 VINP.n165 4.5005
R43762 VINP.n356 VINP.n165 4.5005
R43763 VINP.n237 VINP.n165 4.5005
R43764 VINP.n358 VINP.n165 4.5005
R43765 VINP.n236 VINP.n165 4.5005
R43766 VINP.n360 VINP.n165 4.5005
R43767 VINP.n235 VINP.n165 4.5005
R43768 VINP.n362 VINP.n165 4.5005
R43769 VINP.n234 VINP.n165 4.5005
R43770 VINP.n364 VINP.n165 4.5005
R43771 VINP.n233 VINP.n165 4.5005
R43772 VINP.n366 VINP.n165 4.5005
R43773 VINP.n232 VINP.n165 4.5005
R43774 VINP.n368 VINP.n165 4.5005
R43775 VINP.n231 VINP.n165 4.5005
R43776 VINP.n370 VINP.n165 4.5005
R43777 VINP.n230 VINP.n165 4.5005
R43778 VINP.n372 VINP.n165 4.5005
R43779 VINP.n229 VINP.n165 4.5005
R43780 VINP.n374 VINP.n165 4.5005
R43781 VINP.n228 VINP.n165 4.5005
R43782 VINP.n376 VINP.n165 4.5005
R43783 VINP.n227 VINP.n165 4.5005
R43784 VINP.n378 VINP.n165 4.5005
R43785 VINP.n226 VINP.n165 4.5005
R43786 VINP.n380 VINP.n165 4.5005
R43787 VINP.n225 VINP.n165 4.5005
R43788 VINP.n382 VINP.n165 4.5005
R43789 VINP.n224 VINP.n165 4.5005
R43790 VINP.n384 VINP.n165 4.5005
R43791 VINP.n223 VINP.n165 4.5005
R43792 VINP.n386 VINP.n165 4.5005
R43793 VINP.n222 VINP.n165 4.5005
R43794 VINP.n388 VINP.n165 4.5005
R43795 VINP.n221 VINP.n165 4.5005
R43796 VINP.n390 VINP.n165 4.5005
R43797 VINP.n220 VINP.n165 4.5005
R43798 VINP.n392 VINP.n165 4.5005
R43799 VINP.n219 VINP.n165 4.5005
R43800 VINP.n394 VINP.n165 4.5005
R43801 VINP.n218 VINP.n165 4.5005
R43802 VINP.n396 VINP.n165 4.5005
R43803 VINP.n217 VINP.n165 4.5005
R43804 VINP.n398 VINP.n165 4.5005
R43805 VINP.n216 VINP.n165 4.5005
R43806 VINP.n400 VINP.n165 4.5005
R43807 VINP.n215 VINP.n165 4.5005
R43808 VINP.n654 VINP.n165 4.5005
R43809 VINP.n656 VINP.n165 4.5005
R43810 VINP.n165 VINP.n0 4.5005
R43811 VINP.n278 VINP.n135 4.5005
R43812 VINP.n276 VINP.n135 4.5005
R43813 VINP.n280 VINP.n135 4.5005
R43814 VINP.n275 VINP.n135 4.5005
R43815 VINP.n282 VINP.n135 4.5005
R43816 VINP.n274 VINP.n135 4.5005
R43817 VINP.n284 VINP.n135 4.5005
R43818 VINP.n273 VINP.n135 4.5005
R43819 VINP.n286 VINP.n135 4.5005
R43820 VINP.n272 VINP.n135 4.5005
R43821 VINP.n288 VINP.n135 4.5005
R43822 VINP.n271 VINP.n135 4.5005
R43823 VINP.n290 VINP.n135 4.5005
R43824 VINP.n270 VINP.n135 4.5005
R43825 VINP.n292 VINP.n135 4.5005
R43826 VINP.n269 VINP.n135 4.5005
R43827 VINP.n294 VINP.n135 4.5005
R43828 VINP.n268 VINP.n135 4.5005
R43829 VINP.n296 VINP.n135 4.5005
R43830 VINP.n267 VINP.n135 4.5005
R43831 VINP.n298 VINP.n135 4.5005
R43832 VINP.n266 VINP.n135 4.5005
R43833 VINP.n300 VINP.n135 4.5005
R43834 VINP.n265 VINP.n135 4.5005
R43835 VINP.n302 VINP.n135 4.5005
R43836 VINP.n264 VINP.n135 4.5005
R43837 VINP.n304 VINP.n135 4.5005
R43838 VINP.n263 VINP.n135 4.5005
R43839 VINP.n306 VINP.n135 4.5005
R43840 VINP.n262 VINP.n135 4.5005
R43841 VINP.n308 VINP.n135 4.5005
R43842 VINP.n261 VINP.n135 4.5005
R43843 VINP.n310 VINP.n135 4.5005
R43844 VINP.n260 VINP.n135 4.5005
R43845 VINP.n312 VINP.n135 4.5005
R43846 VINP.n259 VINP.n135 4.5005
R43847 VINP.n314 VINP.n135 4.5005
R43848 VINP.n258 VINP.n135 4.5005
R43849 VINP.n316 VINP.n135 4.5005
R43850 VINP.n257 VINP.n135 4.5005
R43851 VINP.n318 VINP.n135 4.5005
R43852 VINP.n256 VINP.n135 4.5005
R43853 VINP.n320 VINP.n135 4.5005
R43854 VINP.n255 VINP.n135 4.5005
R43855 VINP.n322 VINP.n135 4.5005
R43856 VINP.n254 VINP.n135 4.5005
R43857 VINP.n324 VINP.n135 4.5005
R43858 VINP.n253 VINP.n135 4.5005
R43859 VINP.n326 VINP.n135 4.5005
R43860 VINP.n252 VINP.n135 4.5005
R43861 VINP.n328 VINP.n135 4.5005
R43862 VINP.n251 VINP.n135 4.5005
R43863 VINP.n330 VINP.n135 4.5005
R43864 VINP.n250 VINP.n135 4.5005
R43865 VINP.n332 VINP.n135 4.5005
R43866 VINP.n249 VINP.n135 4.5005
R43867 VINP.n334 VINP.n135 4.5005
R43868 VINP.n248 VINP.n135 4.5005
R43869 VINP.n336 VINP.n135 4.5005
R43870 VINP.n247 VINP.n135 4.5005
R43871 VINP.n338 VINP.n135 4.5005
R43872 VINP.n246 VINP.n135 4.5005
R43873 VINP.n340 VINP.n135 4.5005
R43874 VINP.n245 VINP.n135 4.5005
R43875 VINP.n342 VINP.n135 4.5005
R43876 VINP.n244 VINP.n135 4.5005
R43877 VINP.n344 VINP.n135 4.5005
R43878 VINP.n243 VINP.n135 4.5005
R43879 VINP.n346 VINP.n135 4.5005
R43880 VINP.n242 VINP.n135 4.5005
R43881 VINP.n348 VINP.n135 4.5005
R43882 VINP.n241 VINP.n135 4.5005
R43883 VINP.n350 VINP.n135 4.5005
R43884 VINP.n240 VINP.n135 4.5005
R43885 VINP.n352 VINP.n135 4.5005
R43886 VINP.n239 VINP.n135 4.5005
R43887 VINP.n354 VINP.n135 4.5005
R43888 VINP.n238 VINP.n135 4.5005
R43889 VINP.n356 VINP.n135 4.5005
R43890 VINP.n237 VINP.n135 4.5005
R43891 VINP.n358 VINP.n135 4.5005
R43892 VINP.n236 VINP.n135 4.5005
R43893 VINP.n360 VINP.n135 4.5005
R43894 VINP.n235 VINP.n135 4.5005
R43895 VINP.n362 VINP.n135 4.5005
R43896 VINP.n234 VINP.n135 4.5005
R43897 VINP.n364 VINP.n135 4.5005
R43898 VINP.n233 VINP.n135 4.5005
R43899 VINP.n366 VINP.n135 4.5005
R43900 VINP.n232 VINP.n135 4.5005
R43901 VINP.n368 VINP.n135 4.5005
R43902 VINP.n231 VINP.n135 4.5005
R43903 VINP.n370 VINP.n135 4.5005
R43904 VINP.n230 VINP.n135 4.5005
R43905 VINP.n372 VINP.n135 4.5005
R43906 VINP.n229 VINP.n135 4.5005
R43907 VINP.n374 VINP.n135 4.5005
R43908 VINP.n228 VINP.n135 4.5005
R43909 VINP.n376 VINP.n135 4.5005
R43910 VINP.n227 VINP.n135 4.5005
R43911 VINP.n378 VINP.n135 4.5005
R43912 VINP.n226 VINP.n135 4.5005
R43913 VINP.n380 VINP.n135 4.5005
R43914 VINP.n225 VINP.n135 4.5005
R43915 VINP.n382 VINP.n135 4.5005
R43916 VINP.n224 VINP.n135 4.5005
R43917 VINP.n384 VINP.n135 4.5005
R43918 VINP.n223 VINP.n135 4.5005
R43919 VINP.n386 VINP.n135 4.5005
R43920 VINP.n222 VINP.n135 4.5005
R43921 VINP.n388 VINP.n135 4.5005
R43922 VINP.n221 VINP.n135 4.5005
R43923 VINP.n390 VINP.n135 4.5005
R43924 VINP.n220 VINP.n135 4.5005
R43925 VINP.n392 VINP.n135 4.5005
R43926 VINP.n219 VINP.n135 4.5005
R43927 VINP.n394 VINP.n135 4.5005
R43928 VINP.n218 VINP.n135 4.5005
R43929 VINP.n396 VINP.n135 4.5005
R43930 VINP.n217 VINP.n135 4.5005
R43931 VINP.n398 VINP.n135 4.5005
R43932 VINP.n216 VINP.n135 4.5005
R43933 VINP.n400 VINP.n135 4.5005
R43934 VINP.n215 VINP.n135 4.5005
R43935 VINP.n654 VINP.n135 4.5005
R43936 VINP.n656 VINP.n135 4.5005
R43937 VINP.n135 VINP.n0 4.5005
R43938 VINP.n278 VINP.n166 4.5005
R43939 VINP.n276 VINP.n166 4.5005
R43940 VINP.n280 VINP.n166 4.5005
R43941 VINP.n275 VINP.n166 4.5005
R43942 VINP.n282 VINP.n166 4.5005
R43943 VINP.n274 VINP.n166 4.5005
R43944 VINP.n284 VINP.n166 4.5005
R43945 VINP.n273 VINP.n166 4.5005
R43946 VINP.n286 VINP.n166 4.5005
R43947 VINP.n272 VINP.n166 4.5005
R43948 VINP.n288 VINP.n166 4.5005
R43949 VINP.n271 VINP.n166 4.5005
R43950 VINP.n290 VINP.n166 4.5005
R43951 VINP.n270 VINP.n166 4.5005
R43952 VINP.n292 VINP.n166 4.5005
R43953 VINP.n269 VINP.n166 4.5005
R43954 VINP.n294 VINP.n166 4.5005
R43955 VINP.n268 VINP.n166 4.5005
R43956 VINP.n296 VINP.n166 4.5005
R43957 VINP.n267 VINP.n166 4.5005
R43958 VINP.n298 VINP.n166 4.5005
R43959 VINP.n266 VINP.n166 4.5005
R43960 VINP.n300 VINP.n166 4.5005
R43961 VINP.n265 VINP.n166 4.5005
R43962 VINP.n302 VINP.n166 4.5005
R43963 VINP.n264 VINP.n166 4.5005
R43964 VINP.n304 VINP.n166 4.5005
R43965 VINP.n263 VINP.n166 4.5005
R43966 VINP.n306 VINP.n166 4.5005
R43967 VINP.n262 VINP.n166 4.5005
R43968 VINP.n308 VINP.n166 4.5005
R43969 VINP.n261 VINP.n166 4.5005
R43970 VINP.n310 VINP.n166 4.5005
R43971 VINP.n260 VINP.n166 4.5005
R43972 VINP.n312 VINP.n166 4.5005
R43973 VINP.n259 VINP.n166 4.5005
R43974 VINP.n314 VINP.n166 4.5005
R43975 VINP.n258 VINP.n166 4.5005
R43976 VINP.n316 VINP.n166 4.5005
R43977 VINP.n257 VINP.n166 4.5005
R43978 VINP.n318 VINP.n166 4.5005
R43979 VINP.n256 VINP.n166 4.5005
R43980 VINP.n320 VINP.n166 4.5005
R43981 VINP.n255 VINP.n166 4.5005
R43982 VINP.n322 VINP.n166 4.5005
R43983 VINP.n254 VINP.n166 4.5005
R43984 VINP.n324 VINP.n166 4.5005
R43985 VINP.n253 VINP.n166 4.5005
R43986 VINP.n326 VINP.n166 4.5005
R43987 VINP.n252 VINP.n166 4.5005
R43988 VINP.n328 VINP.n166 4.5005
R43989 VINP.n251 VINP.n166 4.5005
R43990 VINP.n330 VINP.n166 4.5005
R43991 VINP.n250 VINP.n166 4.5005
R43992 VINP.n332 VINP.n166 4.5005
R43993 VINP.n249 VINP.n166 4.5005
R43994 VINP.n334 VINP.n166 4.5005
R43995 VINP.n248 VINP.n166 4.5005
R43996 VINP.n336 VINP.n166 4.5005
R43997 VINP.n247 VINP.n166 4.5005
R43998 VINP.n338 VINP.n166 4.5005
R43999 VINP.n246 VINP.n166 4.5005
R44000 VINP.n340 VINP.n166 4.5005
R44001 VINP.n245 VINP.n166 4.5005
R44002 VINP.n342 VINP.n166 4.5005
R44003 VINP.n244 VINP.n166 4.5005
R44004 VINP.n344 VINP.n166 4.5005
R44005 VINP.n243 VINP.n166 4.5005
R44006 VINP.n346 VINP.n166 4.5005
R44007 VINP.n242 VINP.n166 4.5005
R44008 VINP.n348 VINP.n166 4.5005
R44009 VINP.n241 VINP.n166 4.5005
R44010 VINP.n350 VINP.n166 4.5005
R44011 VINP.n240 VINP.n166 4.5005
R44012 VINP.n352 VINP.n166 4.5005
R44013 VINP.n239 VINP.n166 4.5005
R44014 VINP.n354 VINP.n166 4.5005
R44015 VINP.n238 VINP.n166 4.5005
R44016 VINP.n356 VINP.n166 4.5005
R44017 VINP.n237 VINP.n166 4.5005
R44018 VINP.n358 VINP.n166 4.5005
R44019 VINP.n236 VINP.n166 4.5005
R44020 VINP.n360 VINP.n166 4.5005
R44021 VINP.n235 VINP.n166 4.5005
R44022 VINP.n362 VINP.n166 4.5005
R44023 VINP.n234 VINP.n166 4.5005
R44024 VINP.n364 VINP.n166 4.5005
R44025 VINP.n233 VINP.n166 4.5005
R44026 VINP.n366 VINP.n166 4.5005
R44027 VINP.n232 VINP.n166 4.5005
R44028 VINP.n368 VINP.n166 4.5005
R44029 VINP.n231 VINP.n166 4.5005
R44030 VINP.n370 VINP.n166 4.5005
R44031 VINP.n230 VINP.n166 4.5005
R44032 VINP.n372 VINP.n166 4.5005
R44033 VINP.n229 VINP.n166 4.5005
R44034 VINP.n374 VINP.n166 4.5005
R44035 VINP.n228 VINP.n166 4.5005
R44036 VINP.n376 VINP.n166 4.5005
R44037 VINP.n227 VINP.n166 4.5005
R44038 VINP.n378 VINP.n166 4.5005
R44039 VINP.n226 VINP.n166 4.5005
R44040 VINP.n380 VINP.n166 4.5005
R44041 VINP.n225 VINP.n166 4.5005
R44042 VINP.n382 VINP.n166 4.5005
R44043 VINP.n224 VINP.n166 4.5005
R44044 VINP.n384 VINP.n166 4.5005
R44045 VINP.n223 VINP.n166 4.5005
R44046 VINP.n386 VINP.n166 4.5005
R44047 VINP.n222 VINP.n166 4.5005
R44048 VINP.n388 VINP.n166 4.5005
R44049 VINP.n221 VINP.n166 4.5005
R44050 VINP.n390 VINP.n166 4.5005
R44051 VINP.n220 VINP.n166 4.5005
R44052 VINP.n392 VINP.n166 4.5005
R44053 VINP.n219 VINP.n166 4.5005
R44054 VINP.n394 VINP.n166 4.5005
R44055 VINP.n218 VINP.n166 4.5005
R44056 VINP.n396 VINP.n166 4.5005
R44057 VINP.n217 VINP.n166 4.5005
R44058 VINP.n398 VINP.n166 4.5005
R44059 VINP.n216 VINP.n166 4.5005
R44060 VINP.n400 VINP.n166 4.5005
R44061 VINP.n215 VINP.n166 4.5005
R44062 VINP.n654 VINP.n166 4.5005
R44063 VINP.n656 VINP.n166 4.5005
R44064 VINP.n166 VINP.n0 4.5005
R44065 VINP.n278 VINP.n134 4.5005
R44066 VINP.n276 VINP.n134 4.5005
R44067 VINP.n280 VINP.n134 4.5005
R44068 VINP.n275 VINP.n134 4.5005
R44069 VINP.n282 VINP.n134 4.5005
R44070 VINP.n274 VINP.n134 4.5005
R44071 VINP.n284 VINP.n134 4.5005
R44072 VINP.n273 VINP.n134 4.5005
R44073 VINP.n286 VINP.n134 4.5005
R44074 VINP.n272 VINP.n134 4.5005
R44075 VINP.n288 VINP.n134 4.5005
R44076 VINP.n271 VINP.n134 4.5005
R44077 VINP.n290 VINP.n134 4.5005
R44078 VINP.n270 VINP.n134 4.5005
R44079 VINP.n292 VINP.n134 4.5005
R44080 VINP.n269 VINP.n134 4.5005
R44081 VINP.n294 VINP.n134 4.5005
R44082 VINP.n268 VINP.n134 4.5005
R44083 VINP.n296 VINP.n134 4.5005
R44084 VINP.n267 VINP.n134 4.5005
R44085 VINP.n298 VINP.n134 4.5005
R44086 VINP.n266 VINP.n134 4.5005
R44087 VINP.n300 VINP.n134 4.5005
R44088 VINP.n265 VINP.n134 4.5005
R44089 VINP.n302 VINP.n134 4.5005
R44090 VINP.n264 VINP.n134 4.5005
R44091 VINP.n304 VINP.n134 4.5005
R44092 VINP.n263 VINP.n134 4.5005
R44093 VINP.n306 VINP.n134 4.5005
R44094 VINP.n262 VINP.n134 4.5005
R44095 VINP.n308 VINP.n134 4.5005
R44096 VINP.n261 VINP.n134 4.5005
R44097 VINP.n310 VINP.n134 4.5005
R44098 VINP.n260 VINP.n134 4.5005
R44099 VINP.n312 VINP.n134 4.5005
R44100 VINP.n259 VINP.n134 4.5005
R44101 VINP.n314 VINP.n134 4.5005
R44102 VINP.n258 VINP.n134 4.5005
R44103 VINP.n316 VINP.n134 4.5005
R44104 VINP.n257 VINP.n134 4.5005
R44105 VINP.n318 VINP.n134 4.5005
R44106 VINP.n256 VINP.n134 4.5005
R44107 VINP.n320 VINP.n134 4.5005
R44108 VINP.n255 VINP.n134 4.5005
R44109 VINP.n322 VINP.n134 4.5005
R44110 VINP.n254 VINP.n134 4.5005
R44111 VINP.n324 VINP.n134 4.5005
R44112 VINP.n253 VINP.n134 4.5005
R44113 VINP.n326 VINP.n134 4.5005
R44114 VINP.n252 VINP.n134 4.5005
R44115 VINP.n328 VINP.n134 4.5005
R44116 VINP.n251 VINP.n134 4.5005
R44117 VINP.n330 VINP.n134 4.5005
R44118 VINP.n250 VINP.n134 4.5005
R44119 VINP.n332 VINP.n134 4.5005
R44120 VINP.n249 VINP.n134 4.5005
R44121 VINP.n334 VINP.n134 4.5005
R44122 VINP.n248 VINP.n134 4.5005
R44123 VINP.n336 VINP.n134 4.5005
R44124 VINP.n247 VINP.n134 4.5005
R44125 VINP.n338 VINP.n134 4.5005
R44126 VINP.n246 VINP.n134 4.5005
R44127 VINP.n340 VINP.n134 4.5005
R44128 VINP.n245 VINP.n134 4.5005
R44129 VINP.n342 VINP.n134 4.5005
R44130 VINP.n244 VINP.n134 4.5005
R44131 VINP.n344 VINP.n134 4.5005
R44132 VINP.n243 VINP.n134 4.5005
R44133 VINP.n346 VINP.n134 4.5005
R44134 VINP.n242 VINP.n134 4.5005
R44135 VINP.n348 VINP.n134 4.5005
R44136 VINP.n241 VINP.n134 4.5005
R44137 VINP.n350 VINP.n134 4.5005
R44138 VINP.n240 VINP.n134 4.5005
R44139 VINP.n352 VINP.n134 4.5005
R44140 VINP.n239 VINP.n134 4.5005
R44141 VINP.n354 VINP.n134 4.5005
R44142 VINP.n238 VINP.n134 4.5005
R44143 VINP.n356 VINP.n134 4.5005
R44144 VINP.n237 VINP.n134 4.5005
R44145 VINP.n358 VINP.n134 4.5005
R44146 VINP.n236 VINP.n134 4.5005
R44147 VINP.n360 VINP.n134 4.5005
R44148 VINP.n235 VINP.n134 4.5005
R44149 VINP.n362 VINP.n134 4.5005
R44150 VINP.n234 VINP.n134 4.5005
R44151 VINP.n364 VINP.n134 4.5005
R44152 VINP.n233 VINP.n134 4.5005
R44153 VINP.n366 VINP.n134 4.5005
R44154 VINP.n232 VINP.n134 4.5005
R44155 VINP.n368 VINP.n134 4.5005
R44156 VINP.n231 VINP.n134 4.5005
R44157 VINP.n370 VINP.n134 4.5005
R44158 VINP.n230 VINP.n134 4.5005
R44159 VINP.n372 VINP.n134 4.5005
R44160 VINP.n229 VINP.n134 4.5005
R44161 VINP.n374 VINP.n134 4.5005
R44162 VINP.n228 VINP.n134 4.5005
R44163 VINP.n376 VINP.n134 4.5005
R44164 VINP.n227 VINP.n134 4.5005
R44165 VINP.n378 VINP.n134 4.5005
R44166 VINP.n226 VINP.n134 4.5005
R44167 VINP.n380 VINP.n134 4.5005
R44168 VINP.n225 VINP.n134 4.5005
R44169 VINP.n382 VINP.n134 4.5005
R44170 VINP.n224 VINP.n134 4.5005
R44171 VINP.n384 VINP.n134 4.5005
R44172 VINP.n223 VINP.n134 4.5005
R44173 VINP.n386 VINP.n134 4.5005
R44174 VINP.n222 VINP.n134 4.5005
R44175 VINP.n388 VINP.n134 4.5005
R44176 VINP.n221 VINP.n134 4.5005
R44177 VINP.n390 VINP.n134 4.5005
R44178 VINP.n220 VINP.n134 4.5005
R44179 VINP.n392 VINP.n134 4.5005
R44180 VINP.n219 VINP.n134 4.5005
R44181 VINP.n394 VINP.n134 4.5005
R44182 VINP.n218 VINP.n134 4.5005
R44183 VINP.n396 VINP.n134 4.5005
R44184 VINP.n217 VINP.n134 4.5005
R44185 VINP.n398 VINP.n134 4.5005
R44186 VINP.n216 VINP.n134 4.5005
R44187 VINP.n400 VINP.n134 4.5005
R44188 VINP.n215 VINP.n134 4.5005
R44189 VINP.n654 VINP.n134 4.5005
R44190 VINP.n656 VINP.n134 4.5005
R44191 VINP.n134 VINP.n0 4.5005
R44192 VINP.n278 VINP.n167 4.5005
R44193 VINP.n276 VINP.n167 4.5005
R44194 VINP.n280 VINP.n167 4.5005
R44195 VINP.n275 VINP.n167 4.5005
R44196 VINP.n282 VINP.n167 4.5005
R44197 VINP.n274 VINP.n167 4.5005
R44198 VINP.n284 VINP.n167 4.5005
R44199 VINP.n273 VINP.n167 4.5005
R44200 VINP.n286 VINP.n167 4.5005
R44201 VINP.n272 VINP.n167 4.5005
R44202 VINP.n288 VINP.n167 4.5005
R44203 VINP.n271 VINP.n167 4.5005
R44204 VINP.n290 VINP.n167 4.5005
R44205 VINP.n270 VINP.n167 4.5005
R44206 VINP.n292 VINP.n167 4.5005
R44207 VINP.n269 VINP.n167 4.5005
R44208 VINP.n294 VINP.n167 4.5005
R44209 VINP.n268 VINP.n167 4.5005
R44210 VINP.n296 VINP.n167 4.5005
R44211 VINP.n267 VINP.n167 4.5005
R44212 VINP.n298 VINP.n167 4.5005
R44213 VINP.n266 VINP.n167 4.5005
R44214 VINP.n300 VINP.n167 4.5005
R44215 VINP.n265 VINP.n167 4.5005
R44216 VINP.n302 VINP.n167 4.5005
R44217 VINP.n264 VINP.n167 4.5005
R44218 VINP.n304 VINP.n167 4.5005
R44219 VINP.n263 VINP.n167 4.5005
R44220 VINP.n306 VINP.n167 4.5005
R44221 VINP.n262 VINP.n167 4.5005
R44222 VINP.n308 VINP.n167 4.5005
R44223 VINP.n261 VINP.n167 4.5005
R44224 VINP.n310 VINP.n167 4.5005
R44225 VINP.n260 VINP.n167 4.5005
R44226 VINP.n312 VINP.n167 4.5005
R44227 VINP.n259 VINP.n167 4.5005
R44228 VINP.n314 VINP.n167 4.5005
R44229 VINP.n258 VINP.n167 4.5005
R44230 VINP.n316 VINP.n167 4.5005
R44231 VINP.n257 VINP.n167 4.5005
R44232 VINP.n318 VINP.n167 4.5005
R44233 VINP.n256 VINP.n167 4.5005
R44234 VINP.n320 VINP.n167 4.5005
R44235 VINP.n255 VINP.n167 4.5005
R44236 VINP.n322 VINP.n167 4.5005
R44237 VINP.n254 VINP.n167 4.5005
R44238 VINP.n324 VINP.n167 4.5005
R44239 VINP.n253 VINP.n167 4.5005
R44240 VINP.n326 VINP.n167 4.5005
R44241 VINP.n252 VINP.n167 4.5005
R44242 VINP.n328 VINP.n167 4.5005
R44243 VINP.n251 VINP.n167 4.5005
R44244 VINP.n330 VINP.n167 4.5005
R44245 VINP.n250 VINP.n167 4.5005
R44246 VINP.n332 VINP.n167 4.5005
R44247 VINP.n249 VINP.n167 4.5005
R44248 VINP.n334 VINP.n167 4.5005
R44249 VINP.n248 VINP.n167 4.5005
R44250 VINP.n336 VINP.n167 4.5005
R44251 VINP.n247 VINP.n167 4.5005
R44252 VINP.n338 VINP.n167 4.5005
R44253 VINP.n246 VINP.n167 4.5005
R44254 VINP.n340 VINP.n167 4.5005
R44255 VINP.n245 VINP.n167 4.5005
R44256 VINP.n342 VINP.n167 4.5005
R44257 VINP.n244 VINP.n167 4.5005
R44258 VINP.n344 VINP.n167 4.5005
R44259 VINP.n243 VINP.n167 4.5005
R44260 VINP.n346 VINP.n167 4.5005
R44261 VINP.n242 VINP.n167 4.5005
R44262 VINP.n348 VINP.n167 4.5005
R44263 VINP.n241 VINP.n167 4.5005
R44264 VINP.n350 VINP.n167 4.5005
R44265 VINP.n240 VINP.n167 4.5005
R44266 VINP.n352 VINP.n167 4.5005
R44267 VINP.n239 VINP.n167 4.5005
R44268 VINP.n354 VINP.n167 4.5005
R44269 VINP.n238 VINP.n167 4.5005
R44270 VINP.n356 VINP.n167 4.5005
R44271 VINP.n237 VINP.n167 4.5005
R44272 VINP.n358 VINP.n167 4.5005
R44273 VINP.n236 VINP.n167 4.5005
R44274 VINP.n360 VINP.n167 4.5005
R44275 VINP.n235 VINP.n167 4.5005
R44276 VINP.n362 VINP.n167 4.5005
R44277 VINP.n234 VINP.n167 4.5005
R44278 VINP.n364 VINP.n167 4.5005
R44279 VINP.n233 VINP.n167 4.5005
R44280 VINP.n366 VINP.n167 4.5005
R44281 VINP.n232 VINP.n167 4.5005
R44282 VINP.n368 VINP.n167 4.5005
R44283 VINP.n231 VINP.n167 4.5005
R44284 VINP.n370 VINP.n167 4.5005
R44285 VINP.n230 VINP.n167 4.5005
R44286 VINP.n372 VINP.n167 4.5005
R44287 VINP.n229 VINP.n167 4.5005
R44288 VINP.n374 VINP.n167 4.5005
R44289 VINP.n228 VINP.n167 4.5005
R44290 VINP.n376 VINP.n167 4.5005
R44291 VINP.n227 VINP.n167 4.5005
R44292 VINP.n378 VINP.n167 4.5005
R44293 VINP.n226 VINP.n167 4.5005
R44294 VINP.n380 VINP.n167 4.5005
R44295 VINP.n225 VINP.n167 4.5005
R44296 VINP.n382 VINP.n167 4.5005
R44297 VINP.n224 VINP.n167 4.5005
R44298 VINP.n384 VINP.n167 4.5005
R44299 VINP.n223 VINP.n167 4.5005
R44300 VINP.n386 VINP.n167 4.5005
R44301 VINP.n222 VINP.n167 4.5005
R44302 VINP.n388 VINP.n167 4.5005
R44303 VINP.n221 VINP.n167 4.5005
R44304 VINP.n390 VINP.n167 4.5005
R44305 VINP.n220 VINP.n167 4.5005
R44306 VINP.n392 VINP.n167 4.5005
R44307 VINP.n219 VINP.n167 4.5005
R44308 VINP.n394 VINP.n167 4.5005
R44309 VINP.n218 VINP.n167 4.5005
R44310 VINP.n396 VINP.n167 4.5005
R44311 VINP.n217 VINP.n167 4.5005
R44312 VINP.n398 VINP.n167 4.5005
R44313 VINP.n216 VINP.n167 4.5005
R44314 VINP.n400 VINP.n167 4.5005
R44315 VINP.n215 VINP.n167 4.5005
R44316 VINP.n654 VINP.n167 4.5005
R44317 VINP.n656 VINP.n167 4.5005
R44318 VINP.n167 VINP.n0 4.5005
R44319 VINP.n278 VINP.n133 4.5005
R44320 VINP.n276 VINP.n133 4.5005
R44321 VINP.n280 VINP.n133 4.5005
R44322 VINP.n275 VINP.n133 4.5005
R44323 VINP.n282 VINP.n133 4.5005
R44324 VINP.n274 VINP.n133 4.5005
R44325 VINP.n284 VINP.n133 4.5005
R44326 VINP.n273 VINP.n133 4.5005
R44327 VINP.n286 VINP.n133 4.5005
R44328 VINP.n272 VINP.n133 4.5005
R44329 VINP.n288 VINP.n133 4.5005
R44330 VINP.n271 VINP.n133 4.5005
R44331 VINP.n290 VINP.n133 4.5005
R44332 VINP.n270 VINP.n133 4.5005
R44333 VINP.n292 VINP.n133 4.5005
R44334 VINP.n269 VINP.n133 4.5005
R44335 VINP.n294 VINP.n133 4.5005
R44336 VINP.n268 VINP.n133 4.5005
R44337 VINP.n296 VINP.n133 4.5005
R44338 VINP.n267 VINP.n133 4.5005
R44339 VINP.n298 VINP.n133 4.5005
R44340 VINP.n266 VINP.n133 4.5005
R44341 VINP.n300 VINP.n133 4.5005
R44342 VINP.n265 VINP.n133 4.5005
R44343 VINP.n302 VINP.n133 4.5005
R44344 VINP.n264 VINP.n133 4.5005
R44345 VINP.n304 VINP.n133 4.5005
R44346 VINP.n263 VINP.n133 4.5005
R44347 VINP.n306 VINP.n133 4.5005
R44348 VINP.n262 VINP.n133 4.5005
R44349 VINP.n308 VINP.n133 4.5005
R44350 VINP.n261 VINP.n133 4.5005
R44351 VINP.n310 VINP.n133 4.5005
R44352 VINP.n260 VINP.n133 4.5005
R44353 VINP.n312 VINP.n133 4.5005
R44354 VINP.n259 VINP.n133 4.5005
R44355 VINP.n314 VINP.n133 4.5005
R44356 VINP.n258 VINP.n133 4.5005
R44357 VINP.n316 VINP.n133 4.5005
R44358 VINP.n257 VINP.n133 4.5005
R44359 VINP.n318 VINP.n133 4.5005
R44360 VINP.n256 VINP.n133 4.5005
R44361 VINP.n320 VINP.n133 4.5005
R44362 VINP.n255 VINP.n133 4.5005
R44363 VINP.n322 VINP.n133 4.5005
R44364 VINP.n254 VINP.n133 4.5005
R44365 VINP.n324 VINP.n133 4.5005
R44366 VINP.n253 VINP.n133 4.5005
R44367 VINP.n326 VINP.n133 4.5005
R44368 VINP.n252 VINP.n133 4.5005
R44369 VINP.n328 VINP.n133 4.5005
R44370 VINP.n251 VINP.n133 4.5005
R44371 VINP.n330 VINP.n133 4.5005
R44372 VINP.n250 VINP.n133 4.5005
R44373 VINP.n332 VINP.n133 4.5005
R44374 VINP.n249 VINP.n133 4.5005
R44375 VINP.n334 VINP.n133 4.5005
R44376 VINP.n248 VINP.n133 4.5005
R44377 VINP.n336 VINP.n133 4.5005
R44378 VINP.n247 VINP.n133 4.5005
R44379 VINP.n338 VINP.n133 4.5005
R44380 VINP.n246 VINP.n133 4.5005
R44381 VINP.n340 VINP.n133 4.5005
R44382 VINP.n245 VINP.n133 4.5005
R44383 VINP.n342 VINP.n133 4.5005
R44384 VINP.n244 VINP.n133 4.5005
R44385 VINP.n344 VINP.n133 4.5005
R44386 VINP.n243 VINP.n133 4.5005
R44387 VINP.n346 VINP.n133 4.5005
R44388 VINP.n242 VINP.n133 4.5005
R44389 VINP.n348 VINP.n133 4.5005
R44390 VINP.n241 VINP.n133 4.5005
R44391 VINP.n350 VINP.n133 4.5005
R44392 VINP.n240 VINP.n133 4.5005
R44393 VINP.n352 VINP.n133 4.5005
R44394 VINP.n239 VINP.n133 4.5005
R44395 VINP.n354 VINP.n133 4.5005
R44396 VINP.n238 VINP.n133 4.5005
R44397 VINP.n356 VINP.n133 4.5005
R44398 VINP.n237 VINP.n133 4.5005
R44399 VINP.n358 VINP.n133 4.5005
R44400 VINP.n236 VINP.n133 4.5005
R44401 VINP.n360 VINP.n133 4.5005
R44402 VINP.n235 VINP.n133 4.5005
R44403 VINP.n362 VINP.n133 4.5005
R44404 VINP.n234 VINP.n133 4.5005
R44405 VINP.n364 VINP.n133 4.5005
R44406 VINP.n233 VINP.n133 4.5005
R44407 VINP.n366 VINP.n133 4.5005
R44408 VINP.n232 VINP.n133 4.5005
R44409 VINP.n368 VINP.n133 4.5005
R44410 VINP.n231 VINP.n133 4.5005
R44411 VINP.n370 VINP.n133 4.5005
R44412 VINP.n230 VINP.n133 4.5005
R44413 VINP.n372 VINP.n133 4.5005
R44414 VINP.n229 VINP.n133 4.5005
R44415 VINP.n374 VINP.n133 4.5005
R44416 VINP.n228 VINP.n133 4.5005
R44417 VINP.n376 VINP.n133 4.5005
R44418 VINP.n227 VINP.n133 4.5005
R44419 VINP.n378 VINP.n133 4.5005
R44420 VINP.n226 VINP.n133 4.5005
R44421 VINP.n380 VINP.n133 4.5005
R44422 VINP.n225 VINP.n133 4.5005
R44423 VINP.n382 VINP.n133 4.5005
R44424 VINP.n224 VINP.n133 4.5005
R44425 VINP.n384 VINP.n133 4.5005
R44426 VINP.n223 VINP.n133 4.5005
R44427 VINP.n386 VINP.n133 4.5005
R44428 VINP.n222 VINP.n133 4.5005
R44429 VINP.n388 VINP.n133 4.5005
R44430 VINP.n221 VINP.n133 4.5005
R44431 VINP.n390 VINP.n133 4.5005
R44432 VINP.n220 VINP.n133 4.5005
R44433 VINP.n392 VINP.n133 4.5005
R44434 VINP.n219 VINP.n133 4.5005
R44435 VINP.n394 VINP.n133 4.5005
R44436 VINP.n218 VINP.n133 4.5005
R44437 VINP.n396 VINP.n133 4.5005
R44438 VINP.n217 VINP.n133 4.5005
R44439 VINP.n398 VINP.n133 4.5005
R44440 VINP.n216 VINP.n133 4.5005
R44441 VINP.n400 VINP.n133 4.5005
R44442 VINP.n215 VINP.n133 4.5005
R44443 VINP.n654 VINP.n133 4.5005
R44444 VINP.n656 VINP.n133 4.5005
R44445 VINP.n133 VINP.n0 4.5005
R44446 VINP.n278 VINP.n168 4.5005
R44447 VINP.n276 VINP.n168 4.5005
R44448 VINP.n280 VINP.n168 4.5005
R44449 VINP.n275 VINP.n168 4.5005
R44450 VINP.n282 VINP.n168 4.5005
R44451 VINP.n274 VINP.n168 4.5005
R44452 VINP.n284 VINP.n168 4.5005
R44453 VINP.n273 VINP.n168 4.5005
R44454 VINP.n286 VINP.n168 4.5005
R44455 VINP.n272 VINP.n168 4.5005
R44456 VINP.n288 VINP.n168 4.5005
R44457 VINP.n271 VINP.n168 4.5005
R44458 VINP.n290 VINP.n168 4.5005
R44459 VINP.n270 VINP.n168 4.5005
R44460 VINP.n292 VINP.n168 4.5005
R44461 VINP.n269 VINP.n168 4.5005
R44462 VINP.n294 VINP.n168 4.5005
R44463 VINP.n268 VINP.n168 4.5005
R44464 VINP.n296 VINP.n168 4.5005
R44465 VINP.n267 VINP.n168 4.5005
R44466 VINP.n298 VINP.n168 4.5005
R44467 VINP.n266 VINP.n168 4.5005
R44468 VINP.n300 VINP.n168 4.5005
R44469 VINP.n265 VINP.n168 4.5005
R44470 VINP.n302 VINP.n168 4.5005
R44471 VINP.n264 VINP.n168 4.5005
R44472 VINP.n304 VINP.n168 4.5005
R44473 VINP.n263 VINP.n168 4.5005
R44474 VINP.n306 VINP.n168 4.5005
R44475 VINP.n262 VINP.n168 4.5005
R44476 VINP.n308 VINP.n168 4.5005
R44477 VINP.n261 VINP.n168 4.5005
R44478 VINP.n310 VINP.n168 4.5005
R44479 VINP.n260 VINP.n168 4.5005
R44480 VINP.n312 VINP.n168 4.5005
R44481 VINP.n259 VINP.n168 4.5005
R44482 VINP.n314 VINP.n168 4.5005
R44483 VINP.n258 VINP.n168 4.5005
R44484 VINP.n316 VINP.n168 4.5005
R44485 VINP.n257 VINP.n168 4.5005
R44486 VINP.n318 VINP.n168 4.5005
R44487 VINP.n256 VINP.n168 4.5005
R44488 VINP.n320 VINP.n168 4.5005
R44489 VINP.n255 VINP.n168 4.5005
R44490 VINP.n322 VINP.n168 4.5005
R44491 VINP.n254 VINP.n168 4.5005
R44492 VINP.n324 VINP.n168 4.5005
R44493 VINP.n253 VINP.n168 4.5005
R44494 VINP.n326 VINP.n168 4.5005
R44495 VINP.n252 VINP.n168 4.5005
R44496 VINP.n328 VINP.n168 4.5005
R44497 VINP.n251 VINP.n168 4.5005
R44498 VINP.n330 VINP.n168 4.5005
R44499 VINP.n250 VINP.n168 4.5005
R44500 VINP.n332 VINP.n168 4.5005
R44501 VINP.n249 VINP.n168 4.5005
R44502 VINP.n334 VINP.n168 4.5005
R44503 VINP.n248 VINP.n168 4.5005
R44504 VINP.n336 VINP.n168 4.5005
R44505 VINP.n247 VINP.n168 4.5005
R44506 VINP.n338 VINP.n168 4.5005
R44507 VINP.n246 VINP.n168 4.5005
R44508 VINP.n340 VINP.n168 4.5005
R44509 VINP.n245 VINP.n168 4.5005
R44510 VINP.n342 VINP.n168 4.5005
R44511 VINP.n244 VINP.n168 4.5005
R44512 VINP.n344 VINP.n168 4.5005
R44513 VINP.n243 VINP.n168 4.5005
R44514 VINP.n346 VINP.n168 4.5005
R44515 VINP.n242 VINP.n168 4.5005
R44516 VINP.n348 VINP.n168 4.5005
R44517 VINP.n241 VINP.n168 4.5005
R44518 VINP.n350 VINP.n168 4.5005
R44519 VINP.n240 VINP.n168 4.5005
R44520 VINP.n352 VINP.n168 4.5005
R44521 VINP.n239 VINP.n168 4.5005
R44522 VINP.n354 VINP.n168 4.5005
R44523 VINP.n238 VINP.n168 4.5005
R44524 VINP.n356 VINP.n168 4.5005
R44525 VINP.n237 VINP.n168 4.5005
R44526 VINP.n358 VINP.n168 4.5005
R44527 VINP.n236 VINP.n168 4.5005
R44528 VINP.n360 VINP.n168 4.5005
R44529 VINP.n235 VINP.n168 4.5005
R44530 VINP.n362 VINP.n168 4.5005
R44531 VINP.n234 VINP.n168 4.5005
R44532 VINP.n364 VINP.n168 4.5005
R44533 VINP.n233 VINP.n168 4.5005
R44534 VINP.n366 VINP.n168 4.5005
R44535 VINP.n232 VINP.n168 4.5005
R44536 VINP.n368 VINP.n168 4.5005
R44537 VINP.n231 VINP.n168 4.5005
R44538 VINP.n370 VINP.n168 4.5005
R44539 VINP.n230 VINP.n168 4.5005
R44540 VINP.n372 VINP.n168 4.5005
R44541 VINP.n229 VINP.n168 4.5005
R44542 VINP.n374 VINP.n168 4.5005
R44543 VINP.n228 VINP.n168 4.5005
R44544 VINP.n376 VINP.n168 4.5005
R44545 VINP.n227 VINP.n168 4.5005
R44546 VINP.n378 VINP.n168 4.5005
R44547 VINP.n226 VINP.n168 4.5005
R44548 VINP.n380 VINP.n168 4.5005
R44549 VINP.n225 VINP.n168 4.5005
R44550 VINP.n382 VINP.n168 4.5005
R44551 VINP.n224 VINP.n168 4.5005
R44552 VINP.n384 VINP.n168 4.5005
R44553 VINP.n223 VINP.n168 4.5005
R44554 VINP.n386 VINP.n168 4.5005
R44555 VINP.n222 VINP.n168 4.5005
R44556 VINP.n388 VINP.n168 4.5005
R44557 VINP.n221 VINP.n168 4.5005
R44558 VINP.n390 VINP.n168 4.5005
R44559 VINP.n220 VINP.n168 4.5005
R44560 VINP.n392 VINP.n168 4.5005
R44561 VINP.n219 VINP.n168 4.5005
R44562 VINP.n394 VINP.n168 4.5005
R44563 VINP.n218 VINP.n168 4.5005
R44564 VINP.n396 VINP.n168 4.5005
R44565 VINP.n217 VINP.n168 4.5005
R44566 VINP.n398 VINP.n168 4.5005
R44567 VINP.n216 VINP.n168 4.5005
R44568 VINP.n400 VINP.n168 4.5005
R44569 VINP.n215 VINP.n168 4.5005
R44570 VINP.n654 VINP.n168 4.5005
R44571 VINP.n656 VINP.n168 4.5005
R44572 VINP.n168 VINP.n0 4.5005
R44573 VINP.n278 VINP.n132 4.5005
R44574 VINP.n276 VINP.n132 4.5005
R44575 VINP.n280 VINP.n132 4.5005
R44576 VINP.n275 VINP.n132 4.5005
R44577 VINP.n282 VINP.n132 4.5005
R44578 VINP.n274 VINP.n132 4.5005
R44579 VINP.n284 VINP.n132 4.5005
R44580 VINP.n273 VINP.n132 4.5005
R44581 VINP.n286 VINP.n132 4.5005
R44582 VINP.n272 VINP.n132 4.5005
R44583 VINP.n288 VINP.n132 4.5005
R44584 VINP.n271 VINP.n132 4.5005
R44585 VINP.n290 VINP.n132 4.5005
R44586 VINP.n270 VINP.n132 4.5005
R44587 VINP.n292 VINP.n132 4.5005
R44588 VINP.n269 VINP.n132 4.5005
R44589 VINP.n294 VINP.n132 4.5005
R44590 VINP.n268 VINP.n132 4.5005
R44591 VINP.n296 VINP.n132 4.5005
R44592 VINP.n267 VINP.n132 4.5005
R44593 VINP.n298 VINP.n132 4.5005
R44594 VINP.n266 VINP.n132 4.5005
R44595 VINP.n300 VINP.n132 4.5005
R44596 VINP.n265 VINP.n132 4.5005
R44597 VINP.n302 VINP.n132 4.5005
R44598 VINP.n264 VINP.n132 4.5005
R44599 VINP.n304 VINP.n132 4.5005
R44600 VINP.n263 VINP.n132 4.5005
R44601 VINP.n306 VINP.n132 4.5005
R44602 VINP.n262 VINP.n132 4.5005
R44603 VINP.n308 VINP.n132 4.5005
R44604 VINP.n261 VINP.n132 4.5005
R44605 VINP.n310 VINP.n132 4.5005
R44606 VINP.n260 VINP.n132 4.5005
R44607 VINP.n312 VINP.n132 4.5005
R44608 VINP.n259 VINP.n132 4.5005
R44609 VINP.n314 VINP.n132 4.5005
R44610 VINP.n258 VINP.n132 4.5005
R44611 VINP.n316 VINP.n132 4.5005
R44612 VINP.n257 VINP.n132 4.5005
R44613 VINP.n318 VINP.n132 4.5005
R44614 VINP.n256 VINP.n132 4.5005
R44615 VINP.n320 VINP.n132 4.5005
R44616 VINP.n255 VINP.n132 4.5005
R44617 VINP.n322 VINP.n132 4.5005
R44618 VINP.n254 VINP.n132 4.5005
R44619 VINP.n324 VINP.n132 4.5005
R44620 VINP.n253 VINP.n132 4.5005
R44621 VINP.n326 VINP.n132 4.5005
R44622 VINP.n252 VINP.n132 4.5005
R44623 VINP.n328 VINP.n132 4.5005
R44624 VINP.n251 VINP.n132 4.5005
R44625 VINP.n330 VINP.n132 4.5005
R44626 VINP.n250 VINP.n132 4.5005
R44627 VINP.n332 VINP.n132 4.5005
R44628 VINP.n249 VINP.n132 4.5005
R44629 VINP.n334 VINP.n132 4.5005
R44630 VINP.n248 VINP.n132 4.5005
R44631 VINP.n336 VINP.n132 4.5005
R44632 VINP.n247 VINP.n132 4.5005
R44633 VINP.n338 VINP.n132 4.5005
R44634 VINP.n246 VINP.n132 4.5005
R44635 VINP.n340 VINP.n132 4.5005
R44636 VINP.n245 VINP.n132 4.5005
R44637 VINP.n342 VINP.n132 4.5005
R44638 VINP.n244 VINP.n132 4.5005
R44639 VINP.n344 VINP.n132 4.5005
R44640 VINP.n243 VINP.n132 4.5005
R44641 VINP.n346 VINP.n132 4.5005
R44642 VINP.n242 VINP.n132 4.5005
R44643 VINP.n348 VINP.n132 4.5005
R44644 VINP.n241 VINP.n132 4.5005
R44645 VINP.n350 VINP.n132 4.5005
R44646 VINP.n240 VINP.n132 4.5005
R44647 VINP.n352 VINP.n132 4.5005
R44648 VINP.n239 VINP.n132 4.5005
R44649 VINP.n354 VINP.n132 4.5005
R44650 VINP.n238 VINP.n132 4.5005
R44651 VINP.n356 VINP.n132 4.5005
R44652 VINP.n237 VINP.n132 4.5005
R44653 VINP.n358 VINP.n132 4.5005
R44654 VINP.n236 VINP.n132 4.5005
R44655 VINP.n360 VINP.n132 4.5005
R44656 VINP.n235 VINP.n132 4.5005
R44657 VINP.n362 VINP.n132 4.5005
R44658 VINP.n234 VINP.n132 4.5005
R44659 VINP.n364 VINP.n132 4.5005
R44660 VINP.n233 VINP.n132 4.5005
R44661 VINP.n366 VINP.n132 4.5005
R44662 VINP.n232 VINP.n132 4.5005
R44663 VINP.n368 VINP.n132 4.5005
R44664 VINP.n231 VINP.n132 4.5005
R44665 VINP.n370 VINP.n132 4.5005
R44666 VINP.n230 VINP.n132 4.5005
R44667 VINP.n372 VINP.n132 4.5005
R44668 VINP.n229 VINP.n132 4.5005
R44669 VINP.n374 VINP.n132 4.5005
R44670 VINP.n228 VINP.n132 4.5005
R44671 VINP.n376 VINP.n132 4.5005
R44672 VINP.n227 VINP.n132 4.5005
R44673 VINP.n378 VINP.n132 4.5005
R44674 VINP.n226 VINP.n132 4.5005
R44675 VINP.n380 VINP.n132 4.5005
R44676 VINP.n225 VINP.n132 4.5005
R44677 VINP.n382 VINP.n132 4.5005
R44678 VINP.n224 VINP.n132 4.5005
R44679 VINP.n384 VINP.n132 4.5005
R44680 VINP.n223 VINP.n132 4.5005
R44681 VINP.n386 VINP.n132 4.5005
R44682 VINP.n222 VINP.n132 4.5005
R44683 VINP.n388 VINP.n132 4.5005
R44684 VINP.n221 VINP.n132 4.5005
R44685 VINP.n390 VINP.n132 4.5005
R44686 VINP.n220 VINP.n132 4.5005
R44687 VINP.n392 VINP.n132 4.5005
R44688 VINP.n219 VINP.n132 4.5005
R44689 VINP.n394 VINP.n132 4.5005
R44690 VINP.n218 VINP.n132 4.5005
R44691 VINP.n396 VINP.n132 4.5005
R44692 VINP.n217 VINP.n132 4.5005
R44693 VINP.n398 VINP.n132 4.5005
R44694 VINP.n216 VINP.n132 4.5005
R44695 VINP.n400 VINP.n132 4.5005
R44696 VINP.n215 VINP.n132 4.5005
R44697 VINP.n654 VINP.n132 4.5005
R44698 VINP.n656 VINP.n132 4.5005
R44699 VINP.n132 VINP.n0 4.5005
R44700 VINP.n278 VINP.n169 4.5005
R44701 VINP.n276 VINP.n169 4.5005
R44702 VINP.n280 VINP.n169 4.5005
R44703 VINP.n275 VINP.n169 4.5005
R44704 VINP.n282 VINP.n169 4.5005
R44705 VINP.n274 VINP.n169 4.5005
R44706 VINP.n284 VINP.n169 4.5005
R44707 VINP.n273 VINP.n169 4.5005
R44708 VINP.n286 VINP.n169 4.5005
R44709 VINP.n272 VINP.n169 4.5005
R44710 VINP.n288 VINP.n169 4.5005
R44711 VINP.n271 VINP.n169 4.5005
R44712 VINP.n290 VINP.n169 4.5005
R44713 VINP.n270 VINP.n169 4.5005
R44714 VINP.n292 VINP.n169 4.5005
R44715 VINP.n269 VINP.n169 4.5005
R44716 VINP.n294 VINP.n169 4.5005
R44717 VINP.n268 VINP.n169 4.5005
R44718 VINP.n296 VINP.n169 4.5005
R44719 VINP.n267 VINP.n169 4.5005
R44720 VINP.n298 VINP.n169 4.5005
R44721 VINP.n266 VINP.n169 4.5005
R44722 VINP.n300 VINP.n169 4.5005
R44723 VINP.n265 VINP.n169 4.5005
R44724 VINP.n302 VINP.n169 4.5005
R44725 VINP.n264 VINP.n169 4.5005
R44726 VINP.n304 VINP.n169 4.5005
R44727 VINP.n263 VINP.n169 4.5005
R44728 VINP.n306 VINP.n169 4.5005
R44729 VINP.n262 VINP.n169 4.5005
R44730 VINP.n308 VINP.n169 4.5005
R44731 VINP.n261 VINP.n169 4.5005
R44732 VINP.n310 VINP.n169 4.5005
R44733 VINP.n260 VINP.n169 4.5005
R44734 VINP.n312 VINP.n169 4.5005
R44735 VINP.n259 VINP.n169 4.5005
R44736 VINP.n314 VINP.n169 4.5005
R44737 VINP.n258 VINP.n169 4.5005
R44738 VINP.n316 VINP.n169 4.5005
R44739 VINP.n257 VINP.n169 4.5005
R44740 VINP.n318 VINP.n169 4.5005
R44741 VINP.n256 VINP.n169 4.5005
R44742 VINP.n320 VINP.n169 4.5005
R44743 VINP.n255 VINP.n169 4.5005
R44744 VINP.n322 VINP.n169 4.5005
R44745 VINP.n254 VINP.n169 4.5005
R44746 VINP.n324 VINP.n169 4.5005
R44747 VINP.n253 VINP.n169 4.5005
R44748 VINP.n326 VINP.n169 4.5005
R44749 VINP.n252 VINP.n169 4.5005
R44750 VINP.n328 VINP.n169 4.5005
R44751 VINP.n251 VINP.n169 4.5005
R44752 VINP.n330 VINP.n169 4.5005
R44753 VINP.n250 VINP.n169 4.5005
R44754 VINP.n332 VINP.n169 4.5005
R44755 VINP.n249 VINP.n169 4.5005
R44756 VINP.n334 VINP.n169 4.5005
R44757 VINP.n248 VINP.n169 4.5005
R44758 VINP.n336 VINP.n169 4.5005
R44759 VINP.n247 VINP.n169 4.5005
R44760 VINP.n338 VINP.n169 4.5005
R44761 VINP.n246 VINP.n169 4.5005
R44762 VINP.n340 VINP.n169 4.5005
R44763 VINP.n245 VINP.n169 4.5005
R44764 VINP.n342 VINP.n169 4.5005
R44765 VINP.n244 VINP.n169 4.5005
R44766 VINP.n344 VINP.n169 4.5005
R44767 VINP.n243 VINP.n169 4.5005
R44768 VINP.n346 VINP.n169 4.5005
R44769 VINP.n242 VINP.n169 4.5005
R44770 VINP.n348 VINP.n169 4.5005
R44771 VINP.n241 VINP.n169 4.5005
R44772 VINP.n350 VINP.n169 4.5005
R44773 VINP.n240 VINP.n169 4.5005
R44774 VINP.n352 VINP.n169 4.5005
R44775 VINP.n239 VINP.n169 4.5005
R44776 VINP.n354 VINP.n169 4.5005
R44777 VINP.n238 VINP.n169 4.5005
R44778 VINP.n356 VINP.n169 4.5005
R44779 VINP.n237 VINP.n169 4.5005
R44780 VINP.n358 VINP.n169 4.5005
R44781 VINP.n236 VINP.n169 4.5005
R44782 VINP.n360 VINP.n169 4.5005
R44783 VINP.n235 VINP.n169 4.5005
R44784 VINP.n362 VINP.n169 4.5005
R44785 VINP.n234 VINP.n169 4.5005
R44786 VINP.n364 VINP.n169 4.5005
R44787 VINP.n233 VINP.n169 4.5005
R44788 VINP.n366 VINP.n169 4.5005
R44789 VINP.n232 VINP.n169 4.5005
R44790 VINP.n368 VINP.n169 4.5005
R44791 VINP.n231 VINP.n169 4.5005
R44792 VINP.n370 VINP.n169 4.5005
R44793 VINP.n230 VINP.n169 4.5005
R44794 VINP.n372 VINP.n169 4.5005
R44795 VINP.n229 VINP.n169 4.5005
R44796 VINP.n374 VINP.n169 4.5005
R44797 VINP.n228 VINP.n169 4.5005
R44798 VINP.n376 VINP.n169 4.5005
R44799 VINP.n227 VINP.n169 4.5005
R44800 VINP.n378 VINP.n169 4.5005
R44801 VINP.n226 VINP.n169 4.5005
R44802 VINP.n380 VINP.n169 4.5005
R44803 VINP.n225 VINP.n169 4.5005
R44804 VINP.n382 VINP.n169 4.5005
R44805 VINP.n224 VINP.n169 4.5005
R44806 VINP.n384 VINP.n169 4.5005
R44807 VINP.n223 VINP.n169 4.5005
R44808 VINP.n386 VINP.n169 4.5005
R44809 VINP.n222 VINP.n169 4.5005
R44810 VINP.n388 VINP.n169 4.5005
R44811 VINP.n221 VINP.n169 4.5005
R44812 VINP.n390 VINP.n169 4.5005
R44813 VINP.n220 VINP.n169 4.5005
R44814 VINP.n392 VINP.n169 4.5005
R44815 VINP.n219 VINP.n169 4.5005
R44816 VINP.n394 VINP.n169 4.5005
R44817 VINP.n218 VINP.n169 4.5005
R44818 VINP.n396 VINP.n169 4.5005
R44819 VINP.n217 VINP.n169 4.5005
R44820 VINP.n398 VINP.n169 4.5005
R44821 VINP.n216 VINP.n169 4.5005
R44822 VINP.n400 VINP.n169 4.5005
R44823 VINP.n215 VINP.n169 4.5005
R44824 VINP.n654 VINP.n169 4.5005
R44825 VINP.n656 VINP.n169 4.5005
R44826 VINP.n169 VINP.n0 4.5005
R44827 VINP.n278 VINP.n131 4.5005
R44828 VINP.n276 VINP.n131 4.5005
R44829 VINP.n280 VINP.n131 4.5005
R44830 VINP.n275 VINP.n131 4.5005
R44831 VINP.n282 VINP.n131 4.5005
R44832 VINP.n274 VINP.n131 4.5005
R44833 VINP.n284 VINP.n131 4.5005
R44834 VINP.n273 VINP.n131 4.5005
R44835 VINP.n286 VINP.n131 4.5005
R44836 VINP.n272 VINP.n131 4.5005
R44837 VINP.n288 VINP.n131 4.5005
R44838 VINP.n271 VINP.n131 4.5005
R44839 VINP.n290 VINP.n131 4.5005
R44840 VINP.n270 VINP.n131 4.5005
R44841 VINP.n292 VINP.n131 4.5005
R44842 VINP.n269 VINP.n131 4.5005
R44843 VINP.n294 VINP.n131 4.5005
R44844 VINP.n268 VINP.n131 4.5005
R44845 VINP.n296 VINP.n131 4.5005
R44846 VINP.n267 VINP.n131 4.5005
R44847 VINP.n298 VINP.n131 4.5005
R44848 VINP.n266 VINP.n131 4.5005
R44849 VINP.n300 VINP.n131 4.5005
R44850 VINP.n265 VINP.n131 4.5005
R44851 VINP.n302 VINP.n131 4.5005
R44852 VINP.n264 VINP.n131 4.5005
R44853 VINP.n304 VINP.n131 4.5005
R44854 VINP.n263 VINP.n131 4.5005
R44855 VINP.n306 VINP.n131 4.5005
R44856 VINP.n262 VINP.n131 4.5005
R44857 VINP.n308 VINP.n131 4.5005
R44858 VINP.n261 VINP.n131 4.5005
R44859 VINP.n310 VINP.n131 4.5005
R44860 VINP.n260 VINP.n131 4.5005
R44861 VINP.n312 VINP.n131 4.5005
R44862 VINP.n259 VINP.n131 4.5005
R44863 VINP.n314 VINP.n131 4.5005
R44864 VINP.n258 VINP.n131 4.5005
R44865 VINP.n316 VINP.n131 4.5005
R44866 VINP.n257 VINP.n131 4.5005
R44867 VINP.n318 VINP.n131 4.5005
R44868 VINP.n256 VINP.n131 4.5005
R44869 VINP.n320 VINP.n131 4.5005
R44870 VINP.n255 VINP.n131 4.5005
R44871 VINP.n322 VINP.n131 4.5005
R44872 VINP.n254 VINP.n131 4.5005
R44873 VINP.n324 VINP.n131 4.5005
R44874 VINP.n253 VINP.n131 4.5005
R44875 VINP.n326 VINP.n131 4.5005
R44876 VINP.n252 VINP.n131 4.5005
R44877 VINP.n328 VINP.n131 4.5005
R44878 VINP.n251 VINP.n131 4.5005
R44879 VINP.n330 VINP.n131 4.5005
R44880 VINP.n250 VINP.n131 4.5005
R44881 VINP.n332 VINP.n131 4.5005
R44882 VINP.n249 VINP.n131 4.5005
R44883 VINP.n334 VINP.n131 4.5005
R44884 VINP.n248 VINP.n131 4.5005
R44885 VINP.n336 VINP.n131 4.5005
R44886 VINP.n247 VINP.n131 4.5005
R44887 VINP.n338 VINP.n131 4.5005
R44888 VINP.n246 VINP.n131 4.5005
R44889 VINP.n340 VINP.n131 4.5005
R44890 VINP.n245 VINP.n131 4.5005
R44891 VINP.n342 VINP.n131 4.5005
R44892 VINP.n244 VINP.n131 4.5005
R44893 VINP.n344 VINP.n131 4.5005
R44894 VINP.n243 VINP.n131 4.5005
R44895 VINP.n346 VINP.n131 4.5005
R44896 VINP.n242 VINP.n131 4.5005
R44897 VINP.n348 VINP.n131 4.5005
R44898 VINP.n241 VINP.n131 4.5005
R44899 VINP.n350 VINP.n131 4.5005
R44900 VINP.n240 VINP.n131 4.5005
R44901 VINP.n352 VINP.n131 4.5005
R44902 VINP.n239 VINP.n131 4.5005
R44903 VINP.n354 VINP.n131 4.5005
R44904 VINP.n238 VINP.n131 4.5005
R44905 VINP.n356 VINP.n131 4.5005
R44906 VINP.n237 VINP.n131 4.5005
R44907 VINP.n358 VINP.n131 4.5005
R44908 VINP.n236 VINP.n131 4.5005
R44909 VINP.n360 VINP.n131 4.5005
R44910 VINP.n235 VINP.n131 4.5005
R44911 VINP.n362 VINP.n131 4.5005
R44912 VINP.n234 VINP.n131 4.5005
R44913 VINP.n364 VINP.n131 4.5005
R44914 VINP.n233 VINP.n131 4.5005
R44915 VINP.n366 VINP.n131 4.5005
R44916 VINP.n232 VINP.n131 4.5005
R44917 VINP.n368 VINP.n131 4.5005
R44918 VINP.n231 VINP.n131 4.5005
R44919 VINP.n370 VINP.n131 4.5005
R44920 VINP.n230 VINP.n131 4.5005
R44921 VINP.n372 VINP.n131 4.5005
R44922 VINP.n229 VINP.n131 4.5005
R44923 VINP.n374 VINP.n131 4.5005
R44924 VINP.n228 VINP.n131 4.5005
R44925 VINP.n376 VINP.n131 4.5005
R44926 VINP.n227 VINP.n131 4.5005
R44927 VINP.n378 VINP.n131 4.5005
R44928 VINP.n226 VINP.n131 4.5005
R44929 VINP.n380 VINP.n131 4.5005
R44930 VINP.n225 VINP.n131 4.5005
R44931 VINP.n382 VINP.n131 4.5005
R44932 VINP.n224 VINP.n131 4.5005
R44933 VINP.n384 VINP.n131 4.5005
R44934 VINP.n223 VINP.n131 4.5005
R44935 VINP.n386 VINP.n131 4.5005
R44936 VINP.n222 VINP.n131 4.5005
R44937 VINP.n388 VINP.n131 4.5005
R44938 VINP.n221 VINP.n131 4.5005
R44939 VINP.n390 VINP.n131 4.5005
R44940 VINP.n220 VINP.n131 4.5005
R44941 VINP.n392 VINP.n131 4.5005
R44942 VINP.n219 VINP.n131 4.5005
R44943 VINP.n394 VINP.n131 4.5005
R44944 VINP.n218 VINP.n131 4.5005
R44945 VINP.n396 VINP.n131 4.5005
R44946 VINP.n217 VINP.n131 4.5005
R44947 VINP.n398 VINP.n131 4.5005
R44948 VINP.n216 VINP.n131 4.5005
R44949 VINP.n400 VINP.n131 4.5005
R44950 VINP.n215 VINP.n131 4.5005
R44951 VINP.n654 VINP.n131 4.5005
R44952 VINP.n656 VINP.n131 4.5005
R44953 VINP.n131 VINP.n0 4.5005
R44954 VINP.n278 VINP.n170 4.5005
R44955 VINP.n276 VINP.n170 4.5005
R44956 VINP.n280 VINP.n170 4.5005
R44957 VINP.n275 VINP.n170 4.5005
R44958 VINP.n282 VINP.n170 4.5005
R44959 VINP.n274 VINP.n170 4.5005
R44960 VINP.n284 VINP.n170 4.5005
R44961 VINP.n273 VINP.n170 4.5005
R44962 VINP.n286 VINP.n170 4.5005
R44963 VINP.n272 VINP.n170 4.5005
R44964 VINP.n288 VINP.n170 4.5005
R44965 VINP.n271 VINP.n170 4.5005
R44966 VINP.n290 VINP.n170 4.5005
R44967 VINP.n270 VINP.n170 4.5005
R44968 VINP.n292 VINP.n170 4.5005
R44969 VINP.n269 VINP.n170 4.5005
R44970 VINP.n294 VINP.n170 4.5005
R44971 VINP.n268 VINP.n170 4.5005
R44972 VINP.n296 VINP.n170 4.5005
R44973 VINP.n267 VINP.n170 4.5005
R44974 VINP.n298 VINP.n170 4.5005
R44975 VINP.n266 VINP.n170 4.5005
R44976 VINP.n300 VINP.n170 4.5005
R44977 VINP.n265 VINP.n170 4.5005
R44978 VINP.n302 VINP.n170 4.5005
R44979 VINP.n264 VINP.n170 4.5005
R44980 VINP.n304 VINP.n170 4.5005
R44981 VINP.n263 VINP.n170 4.5005
R44982 VINP.n306 VINP.n170 4.5005
R44983 VINP.n262 VINP.n170 4.5005
R44984 VINP.n308 VINP.n170 4.5005
R44985 VINP.n261 VINP.n170 4.5005
R44986 VINP.n310 VINP.n170 4.5005
R44987 VINP.n260 VINP.n170 4.5005
R44988 VINP.n312 VINP.n170 4.5005
R44989 VINP.n259 VINP.n170 4.5005
R44990 VINP.n314 VINP.n170 4.5005
R44991 VINP.n258 VINP.n170 4.5005
R44992 VINP.n316 VINP.n170 4.5005
R44993 VINP.n257 VINP.n170 4.5005
R44994 VINP.n318 VINP.n170 4.5005
R44995 VINP.n256 VINP.n170 4.5005
R44996 VINP.n320 VINP.n170 4.5005
R44997 VINP.n255 VINP.n170 4.5005
R44998 VINP.n322 VINP.n170 4.5005
R44999 VINP.n254 VINP.n170 4.5005
R45000 VINP.n324 VINP.n170 4.5005
R45001 VINP.n253 VINP.n170 4.5005
R45002 VINP.n326 VINP.n170 4.5005
R45003 VINP.n252 VINP.n170 4.5005
R45004 VINP.n328 VINP.n170 4.5005
R45005 VINP.n251 VINP.n170 4.5005
R45006 VINP.n330 VINP.n170 4.5005
R45007 VINP.n250 VINP.n170 4.5005
R45008 VINP.n332 VINP.n170 4.5005
R45009 VINP.n249 VINP.n170 4.5005
R45010 VINP.n334 VINP.n170 4.5005
R45011 VINP.n248 VINP.n170 4.5005
R45012 VINP.n336 VINP.n170 4.5005
R45013 VINP.n247 VINP.n170 4.5005
R45014 VINP.n338 VINP.n170 4.5005
R45015 VINP.n246 VINP.n170 4.5005
R45016 VINP.n340 VINP.n170 4.5005
R45017 VINP.n245 VINP.n170 4.5005
R45018 VINP.n342 VINP.n170 4.5005
R45019 VINP.n244 VINP.n170 4.5005
R45020 VINP.n344 VINP.n170 4.5005
R45021 VINP.n243 VINP.n170 4.5005
R45022 VINP.n346 VINP.n170 4.5005
R45023 VINP.n242 VINP.n170 4.5005
R45024 VINP.n348 VINP.n170 4.5005
R45025 VINP.n241 VINP.n170 4.5005
R45026 VINP.n350 VINP.n170 4.5005
R45027 VINP.n240 VINP.n170 4.5005
R45028 VINP.n352 VINP.n170 4.5005
R45029 VINP.n239 VINP.n170 4.5005
R45030 VINP.n354 VINP.n170 4.5005
R45031 VINP.n238 VINP.n170 4.5005
R45032 VINP.n356 VINP.n170 4.5005
R45033 VINP.n237 VINP.n170 4.5005
R45034 VINP.n358 VINP.n170 4.5005
R45035 VINP.n236 VINP.n170 4.5005
R45036 VINP.n360 VINP.n170 4.5005
R45037 VINP.n235 VINP.n170 4.5005
R45038 VINP.n362 VINP.n170 4.5005
R45039 VINP.n234 VINP.n170 4.5005
R45040 VINP.n364 VINP.n170 4.5005
R45041 VINP.n233 VINP.n170 4.5005
R45042 VINP.n366 VINP.n170 4.5005
R45043 VINP.n232 VINP.n170 4.5005
R45044 VINP.n368 VINP.n170 4.5005
R45045 VINP.n231 VINP.n170 4.5005
R45046 VINP.n370 VINP.n170 4.5005
R45047 VINP.n230 VINP.n170 4.5005
R45048 VINP.n372 VINP.n170 4.5005
R45049 VINP.n229 VINP.n170 4.5005
R45050 VINP.n374 VINP.n170 4.5005
R45051 VINP.n228 VINP.n170 4.5005
R45052 VINP.n376 VINP.n170 4.5005
R45053 VINP.n227 VINP.n170 4.5005
R45054 VINP.n378 VINP.n170 4.5005
R45055 VINP.n226 VINP.n170 4.5005
R45056 VINP.n380 VINP.n170 4.5005
R45057 VINP.n225 VINP.n170 4.5005
R45058 VINP.n382 VINP.n170 4.5005
R45059 VINP.n224 VINP.n170 4.5005
R45060 VINP.n384 VINP.n170 4.5005
R45061 VINP.n223 VINP.n170 4.5005
R45062 VINP.n386 VINP.n170 4.5005
R45063 VINP.n222 VINP.n170 4.5005
R45064 VINP.n388 VINP.n170 4.5005
R45065 VINP.n221 VINP.n170 4.5005
R45066 VINP.n390 VINP.n170 4.5005
R45067 VINP.n220 VINP.n170 4.5005
R45068 VINP.n392 VINP.n170 4.5005
R45069 VINP.n219 VINP.n170 4.5005
R45070 VINP.n394 VINP.n170 4.5005
R45071 VINP.n218 VINP.n170 4.5005
R45072 VINP.n396 VINP.n170 4.5005
R45073 VINP.n217 VINP.n170 4.5005
R45074 VINP.n398 VINP.n170 4.5005
R45075 VINP.n216 VINP.n170 4.5005
R45076 VINP.n400 VINP.n170 4.5005
R45077 VINP.n215 VINP.n170 4.5005
R45078 VINP.n654 VINP.n170 4.5005
R45079 VINP.n656 VINP.n170 4.5005
R45080 VINP.n170 VINP.n0 4.5005
R45081 VINP.n278 VINP.n130 4.5005
R45082 VINP.n276 VINP.n130 4.5005
R45083 VINP.n280 VINP.n130 4.5005
R45084 VINP.n275 VINP.n130 4.5005
R45085 VINP.n282 VINP.n130 4.5005
R45086 VINP.n274 VINP.n130 4.5005
R45087 VINP.n284 VINP.n130 4.5005
R45088 VINP.n273 VINP.n130 4.5005
R45089 VINP.n286 VINP.n130 4.5005
R45090 VINP.n272 VINP.n130 4.5005
R45091 VINP.n288 VINP.n130 4.5005
R45092 VINP.n271 VINP.n130 4.5005
R45093 VINP.n290 VINP.n130 4.5005
R45094 VINP.n270 VINP.n130 4.5005
R45095 VINP.n292 VINP.n130 4.5005
R45096 VINP.n269 VINP.n130 4.5005
R45097 VINP.n294 VINP.n130 4.5005
R45098 VINP.n268 VINP.n130 4.5005
R45099 VINP.n296 VINP.n130 4.5005
R45100 VINP.n267 VINP.n130 4.5005
R45101 VINP.n298 VINP.n130 4.5005
R45102 VINP.n266 VINP.n130 4.5005
R45103 VINP.n300 VINP.n130 4.5005
R45104 VINP.n265 VINP.n130 4.5005
R45105 VINP.n302 VINP.n130 4.5005
R45106 VINP.n264 VINP.n130 4.5005
R45107 VINP.n304 VINP.n130 4.5005
R45108 VINP.n263 VINP.n130 4.5005
R45109 VINP.n306 VINP.n130 4.5005
R45110 VINP.n262 VINP.n130 4.5005
R45111 VINP.n308 VINP.n130 4.5005
R45112 VINP.n261 VINP.n130 4.5005
R45113 VINP.n310 VINP.n130 4.5005
R45114 VINP.n260 VINP.n130 4.5005
R45115 VINP.n312 VINP.n130 4.5005
R45116 VINP.n259 VINP.n130 4.5005
R45117 VINP.n314 VINP.n130 4.5005
R45118 VINP.n258 VINP.n130 4.5005
R45119 VINP.n316 VINP.n130 4.5005
R45120 VINP.n257 VINP.n130 4.5005
R45121 VINP.n318 VINP.n130 4.5005
R45122 VINP.n256 VINP.n130 4.5005
R45123 VINP.n320 VINP.n130 4.5005
R45124 VINP.n255 VINP.n130 4.5005
R45125 VINP.n322 VINP.n130 4.5005
R45126 VINP.n254 VINP.n130 4.5005
R45127 VINP.n324 VINP.n130 4.5005
R45128 VINP.n253 VINP.n130 4.5005
R45129 VINP.n326 VINP.n130 4.5005
R45130 VINP.n252 VINP.n130 4.5005
R45131 VINP.n328 VINP.n130 4.5005
R45132 VINP.n251 VINP.n130 4.5005
R45133 VINP.n330 VINP.n130 4.5005
R45134 VINP.n250 VINP.n130 4.5005
R45135 VINP.n332 VINP.n130 4.5005
R45136 VINP.n249 VINP.n130 4.5005
R45137 VINP.n334 VINP.n130 4.5005
R45138 VINP.n248 VINP.n130 4.5005
R45139 VINP.n336 VINP.n130 4.5005
R45140 VINP.n247 VINP.n130 4.5005
R45141 VINP.n338 VINP.n130 4.5005
R45142 VINP.n246 VINP.n130 4.5005
R45143 VINP.n340 VINP.n130 4.5005
R45144 VINP.n245 VINP.n130 4.5005
R45145 VINP.n342 VINP.n130 4.5005
R45146 VINP.n244 VINP.n130 4.5005
R45147 VINP.n344 VINP.n130 4.5005
R45148 VINP.n243 VINP.n130 4.5005
R45149 VINP.n346 VINP.n130 4.5005
R45150 VINP.n242 VINP.n130 4.5005
R45151 VINP.n348 VINP.n130 4.5005
R45152 VINP.n241 VINP.n130 4.5005
R45153 VINP.n350 VINP.n130 4.5005
R45154 VINP.n240 VINP.n130 4.5005
R45155 VINP.n352 VINP.n130 4.5005
R45156 VINP.n239 VINP.n130 4.5005
R45157 VINP.n354 VINP.n130 4.5005
R45158 VINP.n238 VINP.n130 4.5005
R45159 VINP.n356 VINP.n130 4.5005
R45160 VINP.n237 VINP.n130 4.5005
R45161 VINP.n358 VINP.n130 4.5005
R45162 VINP.n236 VINP.n130 4.5005
R45163 VINP.n360 VINP.n130 4.5005
R45164 VINP.n235 VINP.n130 4.5005
R45165 VINP.n362 VINP.n130 4.5005
R45166 VINP.n234 VINP.n130 4.5005
R45167 VINP.n364 VINP.n130 4.5005
R45168 VINP.n233 VINP.n130 4.5005
R45169 VINP.n366 VINP.n130 4.5005
R45170 VINP.n232 VINP.n130 4.5005
R45171 VINP.n368 VINP.n130 4.5005
R45172 VINP.n231 VINP.n130 4.5005
R45173 VINP.n370 VINP.n130 4.5005
R45174 VINP.n230 VINP.n130 4.5005
R45175 VINP.n372 VINP.n130 4.5005
R45176 VINP.n229 VINP.n130 4.5005
R45177 VINP.n374 VINP.n130 4.5005
R45178 VINP.n228 VINP.n130 4.5005
R45179 VINP.n376 VINP.n130 4.5005
R45180 VINP.n227 VINP.n130 4.5005
R45181 VINP.n378 VINP.n130 4.5005
R45182 VINP.n226 VINP.n130 4.5005
R45183 VINP.n380 VINP.n130 4.5005
R45184 VINP.n225 VINP.n130 4.5005
R45185 VINP.n382 VINP.n130 4.5005
R45186 VINP.n224 VINP.n130 4.5005
R45187 VINP.n384 VINP.n130 4.5005
R45188 VINP.n223 VINP.n130 4.5005
R45189 VINP.n386 VINP.n130 4.5005
R45190 VINP.n222 VINP.n130 4.5005
R45191 VINP.n388 VINP.n130 4.5005
R45192 VINP.n221 VINP.n130 4.5005
R45193 VINP.n390 VINP.n130 4.5005
R45194 VINP.n220 VINP.n130 4.5005
R45195 VINP.n392 VINP.n130 4.5005
R45196 VINP.n219 VINP.n130 4.5005
R45197 VINP.n394 VINP.n130 4.5005
R45198 VINP.n218 VINP.n130 4.5005
R45199 VINP.n396 VINP.n130 4.5005
R45200 VINP.n217 VINP.n130 4.5005
R45201 VINP.n398 VINP.n130 4.5005
R45202 VINP.n216 VINP.n130 4.5005
R45203 VINP.n400 VINP.n130 4.5005
R45204 VINP.n215 VINP.n130 4.5005
R45205 VINP.n654 VINP.n130 4.5005
R45206 VINP.n656 VINP.n130 4.5005
R45207 VINP.n130 VINP.n0 4.5005
R45208 VINP.n278 VINP.n171 4.5005
R45209 VINP.n276 VINP.n171 4.5005
R45210 VINP.n280 VINP.n171 4.5005
R45211 VINP.n275 VINP.n171 4.5005
R45212 VINP.n282 VINP.n171 4.5005
R45213 VINP.n274 VINP.n171 4.5005
R45214 VINP.n284 VINP.n171 4.5005
R45215 VINP.n273 VINP.n171 4.5005
R45216 VINP.n286 VINP.n171 4.5005
R45217 VINP.n272 VINP.n171 4.5005
R45218 VINP.n288 VINP.n171 4.5005
R45219 VINP.n271 VINP.n171 4.5005
R45220 VINP.n290 VINP.n171 4.5005
R45221 VINP.n270 VINP.n171 4.5005
R45222 VINP.n292 VINP.n171 4.5005
R45223 VINP.n269 VINP.n171 4.5005
R45224 VINP.n294 VINP.n171 4.5005
R45225 VINP.n268 VINP.n171 4.5005
R45226 VINP.n296 VINP.n171 4.5005
R45227 VINP.n267 VINP.n171 4.5005
R45228 VINP.n298 VINP.n171 4.5005
R45229 VINP.n266 VINP.n171 4.5005
R45230 VINP.n300 VINP.n171 4.5005
R45231 VINP.n265 VINP.n171 4.5005
R45232 VINP.n302 VINP.n171 4.5005
R45233 VINP.n264 VINP.n171 4.5005
R45234 VINP.n304 VINP.n171 4.5005
R45235 VINP.n263 VINP.n171 4.5005
R45236 VINP.n306 VINP.n171 4.5005
R45237 VINP.n262 VINP.n171 4.5005
R45238 VINP.n308 VINP.n171 4.5005
R45239 VINP.n261 VINP.n171 4.5005
R45240 VINP.n310 VINP.n171 4.5005
R45241 VINP.n260 VINP.n171 4.5005
R45242 VINP.n312 VINP.n171 4.5005
R45243 VINP.n259 VINP.n171 4.5005
R45244 VINP.n314 VINP.n171 4.5005
R45245 VINP.n258 VINP.n171 4.5005
R45246 VINP.n316 VINP.n171 4.5005
R45247 VINP.n257 VINP.n171 4.5005
R45248 VINP.n318 VINP.n171 4.5005
R45249 VINP.n256 VINP.n171 4.5005
R45250 VINP.n320 VINP.n171 4.5005
R45251 VINP.n255 VINP.n171 4.5005
R45252 VINP.n322 VINP.n171 4.5005
R45253 VINP.n254 VINP.n171 4.5005
R45254 VINP.n324 VINP.n171 4.5005
R45255 VINP.n253 VINP.n171 4.5005
R45256 VINP.n326 VINP.n171 4.5005
R45257 VINP.n252 VINP.n171 4.5005
R45258 VINP.n328 VINP.n171 4.5005
R45259 VINP.n251 VINP.n171 4.5005
R45260 VINP.n330 VINP.n171 4.5005
R45261 VINP.n250 VINP.n171 4.5005
R45262 VINP.n332 VINP.n171 4.5005
R45263 VINP.n249 VINP.n171 4.5005
R45264 VINP.n334 VINP.n171 4.5005
R45265 VINP.n248 VINP.n171 4.5005
R45266 VINP.n336 VINP.n171 4.5005
R45267 VINP.n247 VINP.n171 4.5005
R45268 VINP.n338 VINP.n171 4.5005
R45269 VINP.n246 VINP.n171 4.5005
R45270 VINP.n340 VINP.n171 4.5005
R45271 VINP.n245 VINP.n171 4.5005
R45272 VINP.n342 VINP.n171 4.5005
R45273 VINP.n244 VINP.n171 4.5005
R45274 VINP.n344 VINP.n171 4.5005
R45275 VINP.n243 VINP.n171 4.5005
R45276 VINP.n346 VINP.n171 4.5005
R45277 VINP.n242 VINP.n171 4.5005
R45278 VINP.n348 VINP.n171 4.5005
R45279 VINP.n241 VINP.n171 4.5005
R45280 VINP.n350 VINP.n171 4.5005
R45281 VINP.n240 VINP.n171 4.5005
R45282 VINP.n352 VINP.n171 4.5005
R45283 VINP.n239 VINP.n171 4.5005
R45284 VINP.n354 VINP.n171 4.5005
R45285 VINP.n238 VINP.n171 4.5005
R45286 VINP.n356 VINP.n171 4.5005
R45287 VINP.n237 VINP.n171 4.5005
R45288 VINP.n358 VINP.n171 4.5005
R45289 VINP.n236 VINP.n171 4.5005
R45290 VINP.n360 VINP.n171 4.5005
R45291 VINP.n235 VINP.n171 4.5005
R45292 VINP.n362 VINP.n171 4.5005
R45293 VINP.n234 VINP.n171 4.5005
R45294 VINP.n364 VINP.n171 4.5005
R45295 VINP.n233 VINP.n171 4.5005
R45296 VINP.n366 VINP.n171 4.5005
R45297 VINP.n232 VINP.n171 4.5005
R45298 VINP.n368 VINP.n171 4.5005
R45299 VINP.n231 VINP.n171 4.5005
R45300 VINP.n370 VINP.n171 4.5005
R45301 VINP.n230 VINP.n171 4.5005
R45302 VINP.n372 VINP.n171 4.5005
R45303 VINP.n229 VINP.n171 4.5005
R45304 VINP.n374 VINP.n171 4.5005
R45305 VINP.n228 VINP.n171 4.5005
R45306 VINP.n376 VINP.n171 4.5005
R45307 VINP.n227 VINP.n171 4.5005
R45308 VINP.n378 VINP.n171 4.5005
R45309 VINP.n226 VINP.n171 4.5005
R45310 VINP.n380 VINP.n171 4.5005
R45311 VINP.n225 VINP.n171 4.5005
R45312 VINP.n382 VINP.n171 4.5005
R45313 VINP.n224 VINP.n171 4.5005
R45314 VINP.n384 VINP.n171 4.5005
R45315 VINP.n223 VINP.n171 4.5005
R45316 VINP.n386 VINP.n171 4.5005
R45317 VINP.n222 VINP.n171 4.5005
R45318 VINP.n388 VINP.n171 4.5005
R45319 VINP.n221 VINP.n171 4.5005
R45320 VINP.n390 VINP.n171 4.5005
R45321 VINP.n220 VINP.n171 4.5005
R45322 VINP.n392 VINP.n171 4.5005
R45323 VINP.n219 VINP.n171 4.5005
R45324 VINP.n394 VINP.n171 4.5005
R45325 VINP.n218 VINP.n171 4.5005
R45326 VINP.n396 VINP.n171 4.5005
R45327 VINP.n217 VINP.n171 4.5005
R45328 VINP.n398 VINP.n171 4.5005
R45329 VINP.n216 VINP.n171 4.5005
R45330 VINP.n400 VINP.n171 4.5005
R45331 VINP.n215 VINP.n171 4.5005
R45332 VINP.n654 VINP.n171 4.5005
R45333 VINP.n656 VINP.n171 4.5005
R45334 VINP.n171 VINP.n0 4.5005
R45335 VINP.n278 VINP.n129 4.5005
R45336 VINP.n276 VINP.n129 4.5005
R45337 VINP.n280 VINP.n129 4.5005
R45338 VINP.n275 VINP.n129 4.5005
R45339 VINP.n282 VINP.n129 4.5005
R45340 VINP.n274 VINP.n129 4.5005
R45341 VINP.n284 VINP.n129 4.5005
R45342 VINP.n273 VINP.n129 4.5005
R45343 VINP.n286 VINP.n129 4.5005
R45344 VINP.n272 VINP.n129 4.5005
R45345 VINP.n288 VINP.n129 4.5005
R45346 VINP.n271 VINP.n129 4.5005
R45347 VINP.n290 VINP.n129 4.5005
R45348 VINP.n270 VINP.n129 4.5005
R45349 VINP.n292 VINP.n129 4.5005
R45350 VINP.n269 VINP.n129 4.5005
R45351 VINP.n294 VINP.n129 4.5005
R45352 VINP.n268 VINP.n129 4.5005
R45353 VINP.n296 VINP.n129 4.5005
R45354 VINP.n267 VINP.n129 4.5005
R45355 VINP.n298 VINP.n129 4.5005
R45356 VINP.n266 VINP.n129 4.5005
R45357 VINP.n300 VINP.n129 4.5005
R45358 VINP.n265 VINP.n129 4.5005
R45359 VINP.n302 VINP.n129 4.5005
R45360 VINP.n264 VINP.n129 4.5005
R45361 VINP.n304 VINP.n129 4.5005
R45362 VINP.n263 VINP.n129 4.5005
R45363 VINP.n306 VINP.n129 4.5005
R45364 VINP.n262 VINP.n129 4.5005
R45365 VINP.n308 VINP.n129 4.5005
R45366 VINP.n261 VINP.n129 4.5005
R45367 VINP.n310 VINP.n129 4.5005
R45368 VINP.n260 VINP.n129 4.5005
R45369 VINP.n312 VINP.n129 4.5005
R45370 VINP.n259 VINP.n129 4.5005
R45371 VINP.n314 VINP.n129 4.5005
R45372 VINP.n258 VINP.n129 4.5005
R45373 VINP.n316 VINP.n129 4.5005
R45374 VINP.n257 VINP.n129 4.5005
R45375 VINP.n318 VINP.n129 4.5005
R45376 VINP.n256 VINP.n129 4.5005
R45377 VINP.n320 VINP.n129 4.5005
R45378 VINP.n255 VINP.n129 4.5005
R45379 VINP.n322 VINP.n129 4.5005
R45380 VINP.n254 VINP.n129 4.5005
R45381 VINP.n324 VINP.n129 4.5005
R45382 VINP.n253 VINP.n129 4.5005
R45383 VINP.n326 VINP.n129 4.5005
R45384 VINP.n252 VINP.n129 4.5005
R45385 VINP.n328 VINP.n129 4.5005
R45386 VINP.n251 VINP.n129 4.5005
R45387 VINP.n330 VINP.n129 4.5005
R45388 VINP.n250 VINP.n129 4.5005
R45389 VINP.n332 VINP.n129 4.5005
R45390 VINP.n249 VINP.n129 4.5005
R45391 VINP.n334 VINP.n129 4.5005
R45392 VINP.n248 VINP.n129 4.5005
R45393 VINP.n336 VINP.n129 4.5005
R45394 VINP.n247 VINP.n129 4.5005
R45395 VINP.n338 VINP.n129 4.5005
R45396 VINP.n246 VINP.n129 4.5005
R45397 VINP.n340 VINP.n129 4.5005
R45398 VINP.n245 VINP.n129 4.5005
R45399 VINP.n342 VINP.n129 4.5005
R45400 VINP.n244 VINP.n129 4.5005
R45401 VINP.n344 VINP.n129 4.5005
R45402 VINP.n243 VINP.n129 4.5005
R45403 VINP.n346 VINP.n129 4.5005
R45404 VINP.n242 VINP.n129 4.5005
R45405 VINP.n348 VINP.n129 4.5005
R45406 VINP.n241 VINP.n129 4.5005
R45407 VINP.n350 VINP.n129 4.5005
R45408 VINP.n240 VINP.n129 4.5005
R45409 VINP.n352 VINP.n129 4.5005
R45410 VINP.n239 VINP.n129 4.5005
R45411 VINP.n354 VINP.n129 4.5005
R45412 VINP.n238 VINP.n129 4.5005
R45413 VINP.n356 VINP.n129 4.5005
R45414 VINP.n237 VINP.n129 4.5005
R45415 VINP.n358 VINP.n129 4.5005
R45416 VINP.n236 VINP.n129 4.5005
R45417 VINP.n360 VINP.n129 4.5005
R45418 VINP.n235 VINP.n129 4.5005
R45419 VINP.n362 VINP.n129 4.5005
R45420 VINP.n234 VINP.n129 4.5005
R45421 VINP.n364 VINP.n129 4.5005
R45422 VINP.n233 VINP.n129 4.5005
R45423 VINP.n366 VINP.n129 4.5005
R45424 VINP.n232 VINP.n129 4.5005
R45425 VINP.n368 VINP.n129 4.5005
R45426 VINP.n231 VINP.n129 4.5005
R45427 VINP.n370 VINP.n129 4.5005
R45428 VINP.n230 VINP.n129 4.5005
R45429 VINP.n372 VINP.n129 4.5005
R45430 VINP.n229 VINP.n129 4.5005
R45431 VINP.n374 VINP.n129 4.5005
R45432 VINP.n228 VINP.n129 4.5005
R45433 VINP.n376 VINP.n129 4.5005
R45434 VINP.n227 VINP.n129 4.5005
R45435 VINP.n378 VINP.n129 4.5005
R45436 VINP.n226 VINP.n129 4.5005
R45437 VINP.n380 VINP.n129 4.5005
R45438 VINP.n225 VINP.n129 4.5005
R45439 VINP.n382 VINP.n129 4.5005
R45440 VINP.n224 VINP.n129 4.5005
R45441 VINP.n384 VINP.n129 4.5005
R45442 VINP.n223 VINP.n129 4.5005
R45443 VINP.n386 VINP.n129 4.5005
R45444 VINP.n222 VINP.n129 4.5005
R45445 VINP.n388 VINP.n129 4.5005
R45446 VINP.n221 VINP.n129 4.5005
R45447 VINP.n390 VINP.n129 4.5005
R45448 VINP.n220 VINP.n129 4.5005
R45449 VINP.n392 VINP.n129 4.5005
R45450 VINP.n219 VINP.n129 4.5005
R45451 VINP.n394 VINP.n129 4.5005
R45452 VINP.n218 VINP.n129 4.5005
R45453 VINP.n396 VINP.n129 4.5005
R45454 VINP.n217 VINP.n129 4.5005
R45455 VINP.n398 VINP.n129 4.5005
R45456 VINP.n216 VINP.n129 4.5005
R45457 VINP.n400 VINP.n129 4.5005
R45458 VINP.n215 VINP.n129 4.5005
R45459 VINP.n654 VINP.n129 4.5005
R45460 VINP.n656 VINP.n129 4.5005
R45461 VINP.n129 VINP.n0 4.5005
R45462 VINP.n278 VINP.n172 4.5005
R45463 VINP.n276 VINP.n172 4.5005
R45464 VINP.n280 VINP.n172 4.5005
R45465 VINP.n275 VINP.n172 4.5005
R45466 VINP.n282 VINP.n172 4.5005
R45467 VINP.n274 VINP.n172 4.5005
R45468 VINP.n284 VINP.n172 4.5005
R45469 VINP.n273 VINP.n172 4.5005
R45470 VINP.n286 VINP.n172 4.5005
R45471 VINP.n272 VINP.n172 4.5005
R45472 VINP.n288 VINP.n172 4.5005
R45473 VINP.n271 VINP.n172 4.5005
R45474 VINP.n290 VINP.n172 4.5005
R45475 VINP.n270 VINP.n172 4.5005
R45476 VINP.n292 VINP.n172 4.5005
R45477 VINP.n269 VINP.n172 4.5005
R45478 VINP.n294 VINP.n172 4.5005
R45479 VINP.n268 VINP.n172 4.5005
R45480 VINP.n296 VINP.n172 4.5005
R45481 VINP.n267 VINP.n172 4.5005
R45482 VINP.n298 VINP.n172 4.5005
R45483 VINP.n266 VINP.n172 4.5005
R45484 VINP.n300 VINP.n172 4.5005
R45485 VINP.n265 VINP.n172 4.5005
R45486 VINP.n302 VINP.n172 4.5005
R45487 VINP.n264 VINP.n172 4.5005
R45488 VINP.n304 VINP.n172 4.5005
R45489 VINP.n263 VINP.n172 4.5005
R45490 VINP.n306 VINP.n172 4.5005
R45491 VINP.n262 VINP.n172 4.5005
R45492 VINP.n308 VINP.n172 4.5005
R45493 VINP.n261 VINP.n172 4.5005
R45494 VINP.n310 VINP.n172 4.5005
R45495 VINP.n260 VINP.n172 4.5005
R45496 VINP.n312 VINP.n172 4.5005
R45497 VINP.n259 VINP.n172 4.5005
R45498 VINP.n314 VINP.n172 4.5005
R45499 VINP.n258 VINP.n172 4.5005
R45500 VINP.n316 VINP.n172 4.5005
R45501 VINP.n257 VINP.n172 4.5005
R45502 VINP.n318 VINP.n172 4.5005
R45503 VINP.n256 VINP.n172 4.5005
R45504 VINP.n320 VINP.n172 4.5005
R45505 VINP.n255 VINP.n172 4.5005
R45506 VINP.n322 VINP.n172 4.5005
R45507 VINP.n254 VINP.n172 4.5005
R45508 VINP.n324 VINP.n172 4.5005
R45509 VINP.n253 VINP.n172 4.5005
R45510 VINP.n326 VINP.n172 4.5005
R45511 VINP.n252 VINP.n172 4.5005
R45512 VINP.n328 VINP.n172 4.5005
R45513 VINP.n251 VINP.n172 4.5005
R45514 VINP.n330 VINP.n172 4.5005
R45515 VINP.n250 VINP.n172 4.5005
R45516 VINP.n332 VINP.n172 4.5005
R45517 VINP.n249 VINP.n172 4.5005
R45518 VINP.n334 VINP.n172 4.5005
R45519 VINP.n248 VINP.n172 4.5005
R45520 VINP.n336 VINP.n172 4.5005
R45521 VINP.n247 VINP.n172 4.5005
R45522 VINP.n338 VINP.n172 4.5005
R45523 VINP.n246 VINP.n172 4.5005
R45524 VINP.n340 VINP.n172 4.5005
R45525 VINP.n245 VINP.n172 4.5005
R45526 VINP.n342 VINP.n172 4.5005
R45527 VINP.n244 VINP.n172 4.5005
R45528 VINP.n344 VINP.n172 4.5005
R45529 VINP.n243 VINP.n172 4.5005
R45530 VINP.n346 VINP.n172 4.5005
R45531 VINP.n242 VINP.n172 4.5005
R45532 VINP.n348 VINP.n172 4.5005
R45533 VINP.n241 VINP.n172 4.5005
R45534 VINP.n350 VINP.n172 4.5005
R45535 VINP.n240 VINP.n172 4.5005
R45536 VINP.n352 VINP.n172 4.5005
R45537 VINP.n239 VINP.n172 4.5005
R45538 VINP.n354 VINP.n172 4.5005
R45539 VINP.n238 VINP.n172 4.5005
R45540 VINP.n356 VINP.n172 4.5005
R45541 VINP.n237 VINP.n172 4.5005
R45542 VINP.n358 VINP.n172 4.5005
R45543 VINP.n236 VINP.n172 4.5005
R45544 VINP.n360 VINP.n172 4.5005
R45545 VINP.n235 VINP.n172 4.5005
R45546 VINP.n362 VINP.n172 4.5005
R45547 VINP.n234 VINP.n172 4.5005
R45548 VINP.n364 VINP.n172 4.5005
R45549 VINP.n233 VINP.n172 4.5005
R45550 VINP.n366 VINP.n172 4.5005
R45551 VINP.n232 VINP.n172 4.5005
R45552 VINP.n368 VINP.n172 4.5005
R45553 VINP.n231 VINP.n172 4.5005
R45554 VINP.n370 VINP.n172 4.5005
R45555 VINP.n230 VINP.n172 4.5005
R45556 VINP.n372 VINP.n172 4.5005
R45557 VINP.n229 VINP.n172 4.5005
R45558 VINP.n374 VINP.n172 4.5005
R45559 VINP.n228 VINP.n172 4.5005
R45560 VINP.n376 VINP.n172 4.5005
R45561 VINP.n227 VINP.n172 4.5005
R45562 VINP.n378 VINP.n172 4.5005
R45563 VINP.n226 VINP.n172 4.5005
R45564 VINP.n380 VINP.n172 4.5005
R45565 VINP.n225 VINP.n172 4.5005
R45566 VINP.n382 VINP.n172 4.5005
R45567 VINP.n224 VINP.n172 4.5005
R45568 VINP.n384 VINP.n172 4.5005
R45569 VINP.n223 VINP.n172 4.5005
R45570 VINP.n386 VINP.n172 4.5005
R45571 VINP.n222 VINP.n172 4.5005
R45572 VINP.n388 VINP.n172 4.5005
R45573 VINP.n221 VINP.n172 4.5005
R45574 VINP.n390 VINP.n172 4.5005
R45575 VINP.n220 VINP.n172 4.5005
R45576 VINP.n392 VINP.n172 4.5005
R45577 VINP.n219 VINP.n172 4.5005
R45578 VINP.n394 VINP.n172 4.5005
R45579 VINP.n218 VINP.n172 4.5005
R45580 VINP.n396 VINP.n172 4.5005
R45581 VINP.n217 VINP.n172 4.5005
R45582 VINP.n398 VINP.n172 4.5005
R45583 VINP.n216 VINP.n172 4.5005
R45584 VINP.n400 VINP.n172 4.5005
R45585 VINP.n215 VINP.n172 4.5005
R45586 VINP.n654 VINP.n172 4.5005
R45587 VINP.n656 VINP.n172 4.5005
R45588 VINP.n172 VINP.n0 4.5005
R45589 VINP.n278 VINP.n128 4.5005
R45590 VINP.n276 VINP.n128 4.5005
R45591 VINP.n280 VINP.n128 4.5005
R45592 VINP.n275 VINP.n128 4.5005
R45593 VINP.n282 VINP.n128 4.5005
R45594 VINP.n274 VINP.n128 4.5005
R45595 VINP.n284 VINP.n128 4.5005
R45596 VINP.n273 VINP.n128 4.5005
R45597 VINP.n286 VINP.n128 4.5005
R45598 VINP.n272 VINP.n128 4.5005
R45599 VINP.n288 VINP.n128 4.5005
R45600 VINP.n271 VINP.n128 4.5005
R45601 VINP.n290 VINP.n128 4.5005
R45602 VINP.n270 VINP.n128 4.5005
R45603 VINP.n292 VINP.n128 4.5005
R45604 VINP.n269 VINP.n128 4.5005
R45605 VINP.n294 VINP.n128 4.5005
R45606 VINP.n268 VINP.n128 4.5005
R45607 VINP.n296 VINP.n128 4.5005
R45608 VINP.n267 VINP.n128 4.5005
R45609 VINP.n298 VINP.n128 4.5005
R45610 VINP.n266 VINP.n128 4.5005
R45611 VINP.n300 VINP.n128 4.5005
R45612 VINP.n265 VINP.n128 4.5005
R45613 VINP.n302 VINP.n128 4.5005
R45614 VINP.n264 VINP.n128 4.5005
R45615 VINP.n304 VINP.n128 4.5005
R45616 VINP.n263 VINP.n128 4.5005
R45617 VINP.n306 VINP.n128 4.5005
R45618 VINP.n262 VINP.n128 4.5005
R45619 VINP.n308 VINP.n128 4.5005
R45620 VINP.n261 VINP.n128 4.5005
R45621 VINP.n310 VINP.n128 4.5005
R45622 VINP.n260 VINP.n128 4.5005
R45623 VINP.n312 VINP.n128 4.5005
R45624 VINP.n259 VINP.n128 4.5005
R45625 VINP.n314 VINP.n128 4.5005
R45626 VINP.n258 VINP.n128 4.5005
R45627 VINP.n316 VINP.n128 4.5005
R45628 VINP.n257 VINP.n128 4.5005
R45629 VINP.n318 VINP.n128 4.5005
R45630 VINP.n256 VINP.n128 4.5005
R45631 VINP.n320 VINP.n128 4.5005
R45632 VINP.n255 VINP.n128 4.5005
R45633 VINP.n322 VINP.n128 4.5005
R45634 VINP.n254 VINP.n128 4.5005
R45635 VINP.n324 VINP.n128 4.5005
R45636 VINP.n253 VINP.n128 4.5005
R45637 VINP.n326 VINP.n128 4.5005
R45638 VINP.n252 VINP.n128 4.5005
R45639 VINP.n328 VINP.n128 4.5005
R45640 VINP.n251 VINP.n128 4.5005
R45641 VINP.n330 VINP.n128 4.5005
R45642 VINP.n250 VINP.n128 4.5005
R45643 VINP.n332 VINP.n128 4.5005
R45644 VINP.n249 VINP.n128 4.5005
R45645 VINP.n334 VINP.n128 4.5005
R45646 VINP.n248 VINP.n128 4.5005
R45647 VINP.n336 VINP.n128 4.5005
R45648 VINP.n247 VINP.n128 4.5005
R45649 VINP.n338 VINP.n128 4.5005
R45650 VINP.n246 VINP.n128 4.5005
R45651 VINP.n340 VINP.n128 4.5005
R45652 VINP.n245 VINP.n128 4.5005
R45653 VINP.n342 VINP.n128 4.5005
R45654 VINP.n244 VINP.n128 4.5005
R45655 VINP.n344 VINP.n128 4.5005
R45656 VINP.n243 VINP.n128 4.5005
R45657 VINP.n346 VINP.n128 4.5005
R45658 VINP.n242 VINP.n128 4.5005
R45659 VINP.n348 VINP.n128 4.5005
R45660 VINP.n241 VINP.n128 4.5005
R45661 VINP.n350 VINP.n128 4.5005
R45662 VINP.n240 VINP.n128 4.5005
R45663 VINP.n352 VINP.n128 4.5005
R45664 VINP.n239 VINP.n128 4.5005
R45665 VINP.n354 VINP.n128 4.5005
R45666 VINP.n238 VINP.n128 4.5005
R45667 VINP.n356 VINP.n128 4.5005
R45668 VINP.n237 VINP.n128 4.5005
R45669 VINP.n358 VINP.n128 4.5005
R45670 VINP.n236 VINP.n128 4.5005
R45671 VINP.n360 VINP.n128 4.5005
R45672 VINP.n235 VINP.n128 4.5005
R45673 VINP.n362 VINP.n128 4.5005
R45674 VINP.n234 VINP.n128 4.5005
R45675 VINP.n364 VINP.n128 4.5005
R45676 VINP.n233 VINP.n128 4.5005
R45677 VINP.n366 VINP.n128 4.5005
R45678 VINP.n232 VINP.n128 4.5005
R45679 VINP.n368 VINP.n128 4.5005
R45680 VINP.n231 VINP.n128 4.5005
R45681 VINP.n370 VINP.n128 4.5005
R45682 VINP.n230 VINP.n128 4.5005
R45683 VINP.n372 VINP.n128 4.5005
R45684 VINP.n229 VINP.n128 4.5005
R45685 VINP.n374 VINP.n128 4.5005
R45686 VINP.n228 VINP.n128 4.5005
R45687 VINP.n376 VINP.n128 4.5005
R45688 VINP.n227 VINP.n128 4.5005
R45689 VINP.n378 VINP.n128 4.5005
R45690 VINP.n226 VINP.n128 4.5005
R45691 VINP.n380 VINP.n128 4.5005
R45692 VINP.n225 VINP.n128 4.5005
R45693 VINP.n382 VINP.n128 4.5005
R45694 VINP.n224 VINP.n128 4.5005
R45695 VINP.n384 VINP.n128 4.5005
R45696 VINP.n223 VINP.n128 4.5005
R45697 VINP.n386 VINP.n128 4.5005
R45698 VINP.n222 VINP.n128 4.5005
R45699 VINP.n388 VINP.n128 4.5005
R45700 VINP.n221 VINP.n128 4.5005
R45701 VINP.n390 VINP.n128 4.5005
R45702 VINP.n220 VINP.n128 4.5005
R45703 VINP.n392 VINP.n128 4.5005
R45704 VINP.n219 VINP.n128 4.5005
R45705 VINP.n394 VINP.n128 4.5005
R45706 VINP.n218 VINP.n128 4.5005
R45707 VINP.n396 VINP.n128 4.5005
R45708 VINP.n217 VINP.n128 4.5005
R45709 VINP.n398 VINP.n128 4.5005
R45710 VINP.n216 VINP.n128 4.5005
R45711 VINP.n400 VINP.n128 4.5005
R45712 VINP.n215 VINP.n128 4.5005
R45713 VINP.n654 VINP.n128 4.5005
R45714 VINP.n656 VINP.n128 4.5005
R45715 VINP.n128 VINP.n0 4.5005
R45716 VINP.n278 VINP.n173 4.5005
R45717 VINP.n276 VINP.n173 4.5005
R45718 VINP.n280 VINP.n173 4.5005
R45719 VINP.n275 VINP.n173 4.5005
R45720 VINP.n282 VINP.n173 4.5005
R45721 VINP.n274 VINP.n173 4.5005
R45722 VINP.n284 VINP.n173 4.5005
R45723 VINP.n273 VINP.n173 4.5005
R45724 VINP.n286 VINP.n173 4.5005
R45725 VINP.n272 VINP.n173 4.5005
R45726 VINP.n288 VINP.n173 4.5005
R45727 VINP.n271 VINP.n173 4.5005
R45728 VINP.n290 VINP.n173 4.5005
R45729 VINP.n270 VINP.n173 4.5005
R45730 VINP.n292 VINP.n173 4.5005
R45731 VINP.n269 VINP.n173 4.5005
R45732 VINP.n294 VINP.n173 4.5005
R45733 VINP.n268 VINP.n173 4.5005
R45734 VINP.n296 VINP.n173 4.5005
R45735 VINP.n267 VINP.n173 4.5005
R45736 VINP.n298 VINP.n173 4.5005
R45737 VINP.n266 VINP.n173 4.5005
R45738 VINP.n300 VINP.n173 4.5005
R45739 VINP.n265 VINP.n173 4.5005
R45740 VINP.n302 VINP.n173 4.5005
R45741 VINP.n264 VINP.n173 4.5005
R45742 VINP.n304 VINP.n173 4.5005
R45743 VINP.n263 VINP.n173 4.5005
R45744 VINP.n306 VINP.n173 4.5005
R45745 VINP.n262 VINP.n173 4.5005
R45746 VINP.n308 VINP.n173 4.5005
R45747 VINP.n261 VINP.n173 4.5005
R45748 VINP.n310 VINP.n173 4.5005
R45749 VINP.n260 VINP.n173 4.5005
R45750 VINP.n312 VINP.n173 4.5005
R45751 VINP.n259 VINP.n173 4.5005
R45752 VINP.n314 VINP.n173 4.5005
R45753 VINP.n258 VINP.n173 4.5005
R45754 VINP.n316 VINP.n173 4.5005
R45755 VINP.n257 VINP.n173 4.5005
R45756 VINP.n318 VINP.n173 4.5005
R45757 VINP.n256 VINP.n173 4.5005
R45758 VINP.n320 VINP.n173 4.5005
R45759 VINP.n255 VINP.n173 4.5005
R45760 VINP.n322 VINP.n173 4.5005
R45761 VINP.n254 VINP.n173 4.5005
R45762 VINP.n324 VINP.n173 4.5005
R45763 VINP.n253 VINP.n173 4.5005
R45764 VINP.n326 VINP.n173 4.5005
R45765 VINP.n252 VINP.n173 4.5005
R45766 VINP.n328 VINP.n173 4.5005
R45767 VINP.n251 VINP.n173 4.5005
R45768 VINP.n330 VINP.n173 4.5005
R45769 VINP.n250 VINP.n173 4.5005
R45770 VINP.n332 VINP.n173 4.5005
R45771 VINP.n249 VINP.n173 4.5005
R45772 VINP.n334 VINP.n173 4.5005
R45773 VINP.n248 VINP.n173 4.5005
R45774 VINP.n336 VINP.n173 4.5005
R45775 VINP.n247 VINP.n173 4.5005
R45776 VINP.n338 VINP.n173 4.5005
R45777 VINP.n246 VINP.n173 4.5005
R45778 VINP.n340 VINP.n173 4.5005
R45779 VINP.n245 VINP.n173 4.5005
R45780 VINP.n342 VINP.n173 4.5005
R45781 VINP.n244 VINP.n173 4.5005
R45782 VINP.n344 VINP.n173 4.5005
R45783 VINP.n243 VINP.n173 4.5005
R45784 VINP.n346 VINP.n173 4.5005
R45785 VINP.n242 VINP.n173 4.5005
R45786 VINP.n348 VINP.n173 4.5005
R45787 VINP.n241 VINP.n173 4.5005
R45788 VINP.n350 VINP.n173 4.5005
R45789 VINP.n240 VINP.n173 4.5005
R45790 VINP.n352 VINP.n173 4.5005
R45791 VINP.n239 VINP.n173 4.5005
R45792 VINP.n354 VINP.n173 4.5005
R45793 VINP.n238 VINP.n173 4.5005
R45794 VINP.n356 VINP.n173 4.5005
R45795 VINP.n237 VINP.n173 4.5005
R45796 VINP.n358 VINP.n173 4.5005
R45797 VINP.n236 VINP.n173 4.5005
R45798 VINP.n360 VINP.n173 4.5005
R45799 VINP.n235 VINP.n173 4.5005
R45800 VINP.n362 VINP.n173 4.5005
R45801 VINP.n234 VINP.n173 4.5005
R45802 VINP.n364 VINP.n173 4.5005
R45803 VINP.n233 VINP.n173 4.5005
R45804 VINP.n366 VINP.n173 4.5005
R45805 VINP.n232 VINP.n173 4.5005
R45806 VINP.n368 VINP.n173 4.5005
R45807 VINP.n231 VINP.n173 4.5005
R45808 VINP.n370 VINP.n173 4.5005
R45809 VINP.n230 VINP.n173 4.5005
R45810 VINP.n372 VINP.n173 4.5005
R45811 VINP.n229 VINP.n173 4.5005
R45812 VINP.n374 VINP.n173 4.5005
R45813 VINP.n228 VINP.n173 4.5005
R45814 VINP.n376 VINP.n173 4.5005
R45815 VINP.n227 VINP.n173 4.5005
R45816 VINP.n378 VINP.n173 4.5005
R45817 VINP.n226 VINP.n173 4.5005
R45818 VINP.n380 VINP.n173 4.5005
R45819 VINP.n225 VINP.n173 4.5005
R45820 VINP.n382 VINP.n173 4.5005
R45821 VINP.n224 VINP.n173 4.5005
R45822 VINP.n384 VINP.n173 4.5005
R45823 VINP.n223 VINP.n173 4.5005
R45824 VINP.n386 VINP.n173 4.5005
R45825 VINP.n222 VINP.n173 4.5005
R45826 VINP.n388 VINP.n173 4.5005
R45827 VINP.n221 VINP.n173 4.5005
R45828 VINP.n390 VINP.n173 4.5005
R45829 VINP.n220 VINP.n173 4.5005
R45830 VINP.n392 VINP.n173 4.5005
R45831 VINP.n219 VINP.n173 4.5005
R45832 VINP.n394 VINP.n173 4.5005
R45833 VINP.n218 VINP.n173 4.5005
R45834 VINP.n396 VINP.n173 4.5005
R45835 VINP.n217 VINP.n173 4.5005
R45836 VINP.n398 VINP.n173 4.5005
R45837 VINP.n216 VINP.n173 4.5005
R45838 VINP.n400 VINP.n173 4.5005
R45839 VINP.n215 VINP.n173 4.5005
R45840 VINP.n654 VINP.n173 4.5005
R45841 VINP.n656 VINP.n173 4.5005
R45842 VINP.n173 VINP.n0 4.5005
R45843 VINP.n278 VINP.n127 4.5005
R45844 VINP.n276 VINP.n127 4.5005
R45845 VINP.n280 VINP.n127 4.5005
R45846 VINP.n275 VINP.n127 4.5005
R45847 VINP.n282 VINP.n127 4.5005
R45848 VINP.n274 VINP.n127 4.5005
R45849 VINP.n284 VINP.n127 4.5005
R45850 VINP.n273 VINP.n127 4.5005
R45851 VINP.n286 VINP.n127 4.5005
R45852 VINP.n272 VINP.n127 4.5005
R45853 VINP.n288 VINP.n127 4.5005
R45854 VINP.n271 VINP.n127 4.5005
R45855 VINP.n290 VINP.n127 4.5005
R45856 VINP.n270 VINP.n127 4.5005
R45857 VINP.n292 VINP.n127 4.5005
R45858 VINP.n269 VINP.n127 4.5005
R45859 VINP.n294 VINP.n127 4.5005
R45860 VINP.n268 VINP.n127 4.5005
R45861 VINP.n296 VINP.n127 4.5005
R45862 VINP.n267 VINP.n127 4.5005
R45863 VINP.n298 VINP.n127 4.5005
R45864 VINP.n266 VINP.n127 4.5005
R45865 VINP.n300 VINP.n127 4.5005
R45866 VINP.n265 VINP.n127 4.5005
R45867 VINP.n302 VINP.n127 4.5005
R45868 VINP.n264 VINP.n127 4.5005
R45869 VINP.n304 VINP.n127 4.5005
R45870 VINP.n263 VINP.n127 4.5005
R45871 VINP.n306 VINP.n127 4.5005
R45872 VINP.n262 VINP.n127 4.5005
R45873 VINP.n308 VINP.n127 4.5005
R45874 VINP.n261 VINP.n127 4.5005
R45875 VINP.n310 VINP.n127 4.5005
R45876 VINP.n260 VINP.n127 4.5005
R45877 VINP.n312 VINP.n127 4.5005
R45878 VINP.n259 VINP.n127 4.5005
R45879 VINP.n314 VINP.n127 4.5005
R45880 VINP.n258 VINP.n127 4.5005
R45881 VINP.n316 VINP.n127 4.5005
R45882 VINP.n257 VINP.n127 4.5005
R45883 VINP.n318 VINP.n127 4.5005
R45884 VINP.n256 VINP.n127 4.5005
R45885 VINP.n320 VINP.n127 4.5005
R45886 VINP.n255 VINP.n127 4.5005
R45887 VINP.n322 VINP.n127 4.5005
R45888 VINP.n254 VINP.n127 4.5005
R45889 VINP.n324 VINP.n127 4.5005
R45890 VINP.n253 VINP.n127 4.5005
R45891 VINP.n326 VINP.n127 4.5005
R45892 VINP.n252 VINP.n127 4.5005
R45893 VINP.n328 VINP.n127 4.5005
R45894 VINP.n251 VINP.n127 4.5005
R45895 VINP.n330 VINP.n127 4.5005
R45896 VINP.n250 VINP.n127 4.5005
R45897 VINP.n332 VINP.n127 4.5005
R45898 VINP.n249 VINP.n127 4.5005
R45899 VINP.n334 VINP.n127 4.5005
R45900 VINP.n248 VINP.n127 4.5005
R45901 VINP.n336 VINP.n127 4.5005
R45902 VINP.n247 VINP.n127 4.5005
R45903 VINP.n338 VINP.n127 4.5005
R45904 VINP.n246 VINP.n127 4.5005
R45905 VINP.n340 VINP.n127 4.5005
R45906 VINP.n245 VINP.n127 4.5005
R45907 VINP.n342 VINP.n127 4.5005
R45908 VINP.n244 VINP.n127 4.5005
R45909 VINP.n344 VINP.n127 4.5005
R45910 VINP.n243 VINP.n127 4.5005
R45911 VINP.n346 VINP.n127 4.5005
R45912 VINP.n242 VINP.n127 4.5005
R45913 VINP.n348 VINP.n127 4.5005
R45914 VINP.n241 VINP.n127 4.5005
R45915 VINP.n350 VINP.n127 4.5005
R45916 VINP.n240 VINP.n127 4.5005
R45917 VINP.n352 VINP.n127 4.5005
R45918 VINP.n239 VINP.n127 4.5005
R45919 VINP.n354 VINP.n127 4.5005
R45920 VINP.n238 VINP.n127 4.5005
R45921 VINP.n356 VINP.n127 4.5005
R45922 VINP.n237 VINP.n127 4.5005
R45923 VINP.n358 VINP.n127 4.5005
R45924 VINP.n236 VINP.n127 4.5005
R45925 VINP.n360 VINP.n127 4.5005
R45926 VINP.n235 VINP.n127 4.5005
R45927 VINP.n362 VINP.n127 4.5005
R45928 VINP.n234 VINP.n127 4.5005
R45929 VINP.n364 VINP.n127 4.5005
R45930 VINP.n233 VINP.n127 4.5005
R45931 VINP.n366 VINP.n127 4.5005
R45932 VINP.n232 VINP.n127 4.5005
R45933 VINP.n368 VINP.n127 4.5005
R45934 VINP.n231 VINP.n127 4.5005
R45935 VINP.n370 VINP.n127 4.5005
R45936 VINP.n230 VINP.n127 4.5005
R45937 VINP.n372 VINP.n127 4.5005
R45938 VINP.n229 VINP.n127 4.5005
R45939 VINP.n374 VINP.n127 4.5005
R45940 VINP.n228 VINP.n127 4.5005
R45941 VINP.n376 VINP.n127 4.5005
R45942 VINP.n227 VINP.n127 4.5005
R45943 VINP.n378 VINP.n127 4.5005
R45944 VINP.n226 VINP.n127 4.5005
R45945 VINP.n380 VINP.n127 4.5005
R45946 VINP.n225 VINP.n127 4.5005
R45947 VINP.n382 VINP.n127 4.5005
R45948 VINP.n224 VINP.n127 4.5005
R45949 VINP.n384 VINP.n127 4.5005
R45950 VINP.n223 VINP.n127 4.5005
R45951 VINP.n386 VINP.n127 4.5005
R45952 VINP.n222 VINP.n127 4.5005
R45953 VINP.n388 VINP.n127 4.5005
R45954 VINP.n221 VINP.n127 4.5005
R45955 VINP.n390 VINP.n127 4.5005
R45956 VINP.n220 VINP.n127 4.5005
R45957 VINP.n392 VINP.n127 4.5005
R45958 VINP.n219 VINP.n127 4.5005
R45959 VINP.n394 VINP.n127 4.5005
R45960 VINP.n218 VINP.n127 4.5005
R45961 VINP.n396 VINP.n127 4.5005
R45962 VINP.n217 VINP.n127 4.5005
R45963 VINP.n398 VINP.n127 4.5005
R45964 VINP.n216 VINP.n127 4.5005
R45965 VINP.n400 VINP.n127 4.5005
R45966 VINP.n215 VINP.n127 4.5005
R45967 VINP.n654 VINP.n127 4.5005
R45968 VINP.n656 VINP.n127 4.5005
R45969 VINP.n127 VINP.n0 4.5005
R45970 VINP.n278 VINP.n174 4.5005
R45971 VINP.n276 VINP.n174 4.5005
R45972 VINP.n280 VINP.n174 4.5005
R45973 VINP.n275 VINP.n174 4.5005
R45974 VINP.n282 VINP.n174 4.5005
R45975 VINP.n274 VINP.n174 4.5005
R45976 VINP.n284 VINP.n174 4.5005
R45977 VINP.n273 VINP.n174 4.5005
R45978 VINP.n286 VINP.n174 4.5005
R45979 VINP.n272 VINP.n174 4.5005
R45980 VINP.n288 VINP.n174 4.5005
R45981 VINP.n271 VINP.n174 4.5005
R45982 VINP.n290 VINP.n174 4.5005
R45983 VINP.n270 VINP.n174 4.5005
R45984 VINP.n292 VINP.n174 4.5005
R45985 VINP.n269 VINP.n174 4.5005
R45986 VINP.n294 VINP.n174 4.5005
R45987 VINP.n268 VINP.n174 4.5005
R45988 VINP.n296 VINP.n174 4.5005
R45989 VINP.n267 VINP.n174 4.5005
R45990 VINP.n298 VINP.n174 4.5005
R45991 VINP.n266 VINP.n174 4.5005
R45992 VINP.n300 VINP.n174 4.5005
R45993 VINP.n265 VINP.n174 4.5005
R45994 VINP.n302 VINP.n174 4.5005
R45995 VINP.n264 VINP.n174 4.5005
R45996 VINP.n304 VINP.n174 4.5005
R45997 VINP.n263 VINP.n174 4.5005
R45998 VINP.n306 VINP.n174 4.5005
R45999 VINP.n262 VINP.n174 4.5005
R46000 VINP.n308 VINP.n174 4.5005
R46001 VINP.n261 VINP.n174 4.5005
R46002 VINP.n310 VINP.n174 4.5005
R46003 VINP.n260 VINP.n174 4.5005
R46004 VINP.n312 VINP.n174 4.5005
R46005 VINP.n259 VINP.n174 4.5005
R46006 VINP.n314 VINP.n174 4.5005
R46007 VINP.n258 VINP.n174 4.5005
R46008 VINP.n316 VINP.n174 4.5005
R46009 VINP.n257 VINP.n174 4.5005
R46010 VINP.n318 VINP.n174 4.5005
R46011 VINP.n256 VINP.n174 4.5005
R46012 VINP.n320 VINP.n174 4.5005
R46013 VINP.n255 VINP.n174 4.5005
R46014 VINP.n322 VINP.n174 4.5005
R46015 VINP.n254 VINP.n174 4.5005
R46016 VINP.n324 VINP.n174 4.5005
R46017 VINP.n253 VINP.n174 4.5005
R46018 VINP.n326 VINP.n174 4.5005
R46019 VINP.n252 VINP.n174 4.5005
R46020 VINP.n328 VINP.n174 4.5005
R46021 VINP.n251 VINP.n174 4.5005
R46022 VINP.n330 VINP.n174 4.5005
R46023 VINP.n250 VINP.n174 4.5005
R46024 VINP.n332 VINP.n174 4.5005
R46025 VINP.n249 VINP.n174 4.5005
R46026 VINP.n334 VINP.n174 4.5005
R46027 VINP.n248 VINP.n174 4.5005
R46028 VINP.n336 VINP.n174 4.5005
R46029 VINP.n247 VINP.n174 4.5005
R46030 VINP.n338 VINP.n174 4.5005
R46031 VINP.n246 VINP.n174 4.5005
R46032 VINP.n340 VINP.n174 4.5005
R46033 VINP.n245 VINP.n174 4.5005
R46034 VINP.n342 VINP.n174 4.5005
R46035 VINP.n244 VINP.n174 4.5005
R46036 VINP.n344 VINP.n174 4.5005
R46037 VINP.n243 VINP.n174 4.5005
R46038 VINP.n346 VINP.n174 4.5005
R46039 VINP.n242 VINP.n174 4.5005
R46040 VINP.n348 VINP.n174 4.5005
R46041 VINP.n241 VINP.n174 4.5005
R46042 VINP.n350 VINP.n174 4.5005
R46043 VINP.n240 VINP.n174 4.5005
R46044 VINP.n352 VINP.n174 4.5005
R46045 VINP.n239 VINP.n174 4.5005
R46046 VINP.n354 VINP.n174 4.5005
R46047 VINP.n238 VINP.n174 4.5005
R46048 VINP.n356 VINP.n174 4.5005
R46049 VINP.n237 VINP.n174 4.5005
R46050 VINP.n358 VINP.n174 4.5005
R46051 VINP.n236 VINP.n174 4.5005
R46052 VINP.n360 VINP.n174 4.5005
R46053 VINP.n235 VINP.n174 4.5005
R46054 VINP.n362 VINP.n174 4.5005
R46055 VINP.n234 VINP.n174 4.5005
R46056 VINP.n364 VINP.n174 4.5005
R46057 VINP.n233 VINP.n174 4.5005
R46058 VINP.n366 VINP.n174 4.5005
R46059 VINP.n232 VINP.n174 4.5005
R46060 VINP.n368 VINP.n174 4.5005
R46061 VINP.n231 VINP.n174 4.5005
R46062 VINP.n370 VINP.n174 4.5005
R46063 VINP.n230 VINP.n174 4.5005
R46064 VINP.n372 VINP.n174 4.5005
R46065 VINP.n229 VINP.n174 4.5005
R46066 VINP.n374 VINP.n174 4.5005
R46067 VINP.n228 VINP.n174 4.5005
R46068 VINP.n376 VINP.n174 4.5005
R46069 VINP.n227 VINP.n174 4.5005
R46070 VINP.n378 VINP.n174 4.5005
R46071 VINP.n226 VINP.n174 4.5005
R46072 VINP.n380 VINP.n174 4.5005
R46073 VINP.n225 VINP.n174 4.5005
R46074 VINP.n382 VINP.n174 4.5005
R46075 VINP.n224 VINP.n174 4.5005
R46076 VINP.n384 VINP.n174 4.5005
R46077 VINP.n223 VINP.n174 4.5005
R46078 VINP.n386 VINP.n174 4.5005
R46079 VINP.n222 VINP.n174 4.5005
R46080 VINP.n388 VINP.n174 4.5005
R46081 VINP.n221 VINP.n174 4.5005
R46082 VINP.n390 VINP.n174 4.5005
R46083 VINP.n220 VINP.n174 4.5005
R46084 VINP.n392 VINP.n174 4.5005
R46085 VINP.n219 VINP.n174 4.5005
R46086 VINP.n394 VINP.n174 4.5005
R46087 VINP.n218 VINP.n174 4.5005
R46088 VINP.n396 VINP.n174 4.5005
R46089 VINP.n217 VINP.n174 4.5005
R46090 VINP.n398 VINP.n174 4.5005
R46091 VINP.n216 VINP.n174 4.5005
R46092 VINP.n400 VINP.n174 4.5005
R46093 VINP.n215 VINP.n174 4.5005
R46094 VINP.n654 VINP.n174 4.5005
R46095 VINP.n656 VINP.n174 4.5005
R46096 VINP.n174 VINP.n0 4.5005
R46097 VINP.n278 VINP.n126 4.5005
R46098 VINP.n276 VINP.n126 4.5005
R46099 VINP.n280 VINP.n126 4.5005
R46100 VINP.n275 VINP.n126 4.5005
R46101 VINP.n282 VINP.n126 4.5005
R46102 VINP.n274 VINP.n126 4.5005
R46103 VINP.n284 VINP.n126 4.5005
R46104 VINP.n273 VINP.n126 4.5005
R46105 VINP.n286 VINP.n126 4.5005
R46106 VINP.n272 VINP.n126 4.5005
R46107 VINP.n288 VINP.n126 4.5005
R46108 VINP.n271 VINP.n126 4.5005
R46109 VINP.n290 VINP.n126 4.5005
R46110 VINP.n270 VINP.n126 4.5005
R46111 VINP.n292 VINP.n126 4.5005
R46112 VINP.n269 VINP.n126 4.5005
R46113 VINP.n294 VINP.n126 4.5005
R46114 VINP.n268 VINP.n126 4.5005
R46115 VINP.n296 VINP.n126 4.5005
R46116 VINP.n267 VINP.n126 4.5005
R46117 VINP.n298 VINP.n126 4.5005
R46118 VINP.n266 VINP.n126 4.5005
R46119 VINP.n300 VINP.n126 4.5005
R46120 VINP.n265 VINP.n126 4.5005
R46121 VINP.n302 VINP.n126 4.5005
R46122 VINP.n264 VINP.n126 4.5005
R46123 VINP.n304 VINP.n126 4.5005
R46124 VINP.n263 VINP.n126 4.5005
R46125 VINP.n306 VINP.n126 4.5005
R46126 VINP.n262 VINP.n126 4.5005
R46127 VINP.n308 VINP.n126 4.5005
R46128 VINP.n261 VINP.n126 4.5005
R46129 VINP.n310 VINP.n126 4.5005
R46130 VINP.n260 VINP.n126 4.5005
R46131 VINP.n312 VINP.n126 4.5005
R46132 VINP.n259 VINP.n126 4.5005
R46133 VINP.n314 VINP.n126 4.5005
R46134 VINP.n258 VINP.n126 4.5005
R46135 VINP.n316 VINP.n126 4.5005
R46136 VINP.n257 VINP.n126 4.5005
R46137 VINP.n318 VINP.n126 4.5005
R46138 VINP.n256 VINP.n126 4.5005
R46139 VINP.n320 VINP.n126 4.5005
R46140 VINP.n255 VINP.n126 4.5005
R46141 VINP.n322 VINP.n126 4.5005
R46142 VINP.n254 VINP.n126 4.5005
R46143 VINP.n324 VINP.n126 4.5005
R46144 VINP.n253 VINP.n126 4.5005
R46145 VINP.n326 VINP.n126 4.5005
R46146 VINP.n252 VINP.n126 4.5005
R46147 VINP.n328 VINP.n126 4.5005
R46148 VINP.n251 VINP.n126 4.5005
R46149 VINP.n330 VINP.n126 4.5005
R46150 VINP.n250 VINP.n126 4.5005
R46151 VINP.n332 VINP.n126 4.5005
R46152 VINP.n249 VINP.n126 4.5005
R46153 VINP.n334 VINP.n126 4.5005
R46154 VINP.n248 VINP.n126 4.5005
R46155 VINP.n336 VINP.n126 4.5005
R46156 VINP.n247 VINP.n126 4.5005
R46157 VINP.n338 VINP.n126 4.5005
R46158 VINP.n246 VINP.n126 4.5005
R46159 VINP.n340 VINP.n126 4.5005
R46160 VINP.n245 VINP.n126 4.5005
R46161 VINP.n342 VINP.n126 4.5005
R46162 VINP.n244 VINP.n126 4.5005
R46163 VINP.n344 VINP.n126 4.5005
R46164 VINP.n243 VINP.n126 4.5005
R46165 VINP.n346 VINP.n126 4.5005
R46166 VINP.n242 VINP.n126 4.5005
R46167 VINP.n348 VINP.n126 4.5005
R46168 VINP.n241 VINP.n126 4.5005
R46169 VINP.n350 VINP.n126 4.5005
R46170 VINP.n240 VINP.n126 4.5005
R46171 VINP.n352 VINP.n126 4.5005
R46172 VINP.n239 VINP.n126 4.5005
R46173 VINP.n354 VINP.n126 4.5005
R46174 VINP.n238 VINP.n126 4.5005
R46175 VINP.n356 VINP.n126 4.5005
R46176 VINP.n237 VINP.n126 4.5005
R46177 VINP.n358 VINP.n126 4.5005
R46178 VINP.n236 VINP.n126 4.5005
R46179 VINP.n360 VINP.n126 4.5005
R46180 VINP.n235 VINP.n126 4.5005
R46181 VINP.n362 VINP.n126 4.5005
R46182 VINP.n234 VINP.n126 4.5005
R46183 VINP.n364 VINP.n126 4.5005
R46184 VINP.n233 VINP.n126 4.5005
R46185 VINP.n366 VINP.n126 4.5005
R46186 VINP.n232 VINP.n126 4.5005
R46187 VINP.n368 VINP.n126 4.5005
R46188 VINP.n231 VINP.n126 4.5005
R46189 VINP.n370 VINP.n126 4.5005
R46190 VINP.n230 VINP.n126 4.5005
R46191 VINP.n372 VINP.n126 4.5005
R46192 VINP.n229 VINP.n126 4.5005
R46193 VINP.n374 VINP.n126 4.5005
R46194 VINP.n228 VINP.n126 4.5005
R46195 VINP.n376 VINP.n126 4.5005
R46196 VINP.n227 VINP.n126 4.5005
R46197 VINP.n378 VINP.n126 4.5005
R46198 VINP.n226 VINP.n126 4.5005
R46199 VINP.n380 VINP.n126 4.5005
R46200 VINP.n225 VINP.n126 4.5005
R46201 VINP.n382 VINP.n126 4.5005
R46202 VINP.n224 VINP.n126 4.5005
R46203 VINP.n384 VINP.n126 4.5005
R46204 VINP.n223 VINP.n126 4.5005
R46205 VINP.n386 VINP.n126 4.5005
R46206 VINP.n222 VINP.n126 4.5005
R46207 VINP.n388 VINP.n126 4.5005
R46208 VINP.n221 VINP.n126 4.5005
R46209 VINP.n390 VINP.n126 4.5005
R46210 VINP.n220 VINP.n126 4.5005
R46211 VINP.n392 VINP.n126 4.5005
R46212 VINP.n219 VINP.n126 4.5005
R46213 VINP.n394 VINP.n126 4.5005
R46214 VINP.n218 VINP.n126 4.5005
R46215 VINP.n396 VINP.n126 4.5005
R46216 VINP.n217 VINP.n126 4.5005
R46217 VINP.n398 VINP.n126 4.5005
R46218 VINP.n216 VINP.n126 4.5005
R46219 VINP.n400 VINP.n126 4.5005
R46220 VINP.n215 VINP.n126 4.5005
R46221 VINP.n654 VINP.n126 4.5005
R46222 VINP.n656 VINP.n126 4.5005
R46223 VINP.n126 VINP.n0 4.5005
R46224 VINP.n278 VINP.n175 4.5005
R46225 VINP.n276 VINP.n175 4.5005
R46226 VINP.n280 VINP.n175 4.5005
R46227 VINP.n275 VINP.n175 4.5005
R46228 VINP.n282 VINP.n175 4.5005
R46229 VINP.n274 VINP.n175 4.5005
R46230 VINP.n284 VINP.n175 4.5005
R46231 VINP.n273 VINP.n175 4.5005
R46232 VINP.n286 VINP.n175 4.5005
R46233 VINP.n272 VINP.n175 4.5005
R46234 VINP.n288 VINP.n175 4.5005
R46235 VINP.n271 VINP.n175 4.5005
R46236 VINP.n290 VINP.n175 4.5005
R46237 VINP.n270 VINP.n175 4.5005
R46238 VINP.n292 VINP.n175 4.5005
R46239 VINP.n269 VINP.n175 4.5005
R46240 VINP.n294 VINP.n175 4.5005
R46241 VINP.n268 VINP.n175 4.5005
R46242 VINP.n296 VINP.n175 4.5005
R46243 VINP.n267 VINP.n175 4.5005
R46244 VINP.n298 VINP.n175 4.5005
R46245 VINP.n266 VINP.n175 4.5005
R46246 VINP.n300 VINP.n175 4.5005
R46247 VINP.n265 VINP.n175 4.5005
R46248 VINP.n302 VINP.n175 4.5005
R46249 VINP.n264 VINP.n175 4.5005
R46250 VINP.n304 VINP.n175 4.5005
R46251 VINP.n263 VINP.n175 4.5005
R46252 VINP.n306 VINP.n175 4.5005
R46253 VINP.n262 VINP.n175 4.5005
R46254 VINP.n308 VINP.n175 4.5005
R46255 VINP.n261 VINP.n175 4.5005
R46256 VINP.n310 VINP.n175 4.5005
R46257 VINP.n260 VINP.n175 4.5005
R46258 VINP.n312 VINP.n175 4.5005
R46259 VINP.n259 VINP.n175 4.5005
R46260 VINP.n314 VINP.n175 4.5005
R46261 VINP.n258 VINP.n175 4.5005
R46262 VINP.n316 VINP.n175 4.5005
R46263 VINP.n257 VINP.n175 4.5005
R46264 VINP.n318 VINP.n175 4.5005
R46265 VINP.n256 VINP.n175 4.5005
R46266 VINP.n320 VINP.n175 4.5005
R46267 VINP.n255 VINP.n175 4.5005
R46268 VINP.n322 VINP.n175 4.5005
R46269 VINP.n254 VINP.n175 4.5005
R46270 VINP.n324 VINP.n175 4.5005
R46271 VINP.n253 VINP.n175 4.5005
R46272 VINP.n326 VINP.n175 4.5005
R46273 VINP.n252 VINP.n175 4.5005
R46274 VINP.n328 VINP.n175 4.5005
R46275 VINP.n251 VINP.n175 4.5005
R46276 VINP.n330 VINP.n175 4.5005
R46277 VINP.n250 VINP.n175 4.5005
R46278 VINP.n332 VINP.n175 4.5005
R46279 VINP.n249 VINP.n175 4.5005
R46280 VINP.n334 VINP.n175 4.5005
R46281 VINP.n248 VINP.n175 4.5005
R46282 VINP.n336 VINP.n175 4.5005
R46283 VINP.n247 VINP.n175 4.5005
R46284 VINP.n338 VINP.n175 4.5005
R46285 VINP.n246 VINP.n175 4.5005
R46286 VINP.n340 VINP.n175 4.5005
R46287 VINP.n245 VINP.n175 4.5005
R46288 VINP.n342 VINP.n175 4.5005
R46289 VINP.n244 VINP.n175 4.5005
R46290 VINP.n344 VINP.n175 4.5005
R46291 VINP.n243 VINP.n175 4.5005
R46292 VINP.n346 VINP.n175 4.5005
R46293 VINP.n242 VINP.n175 4.5005
R46294 VINP.n348 VINP.n175 4.5005
R46295 VINP.n241 VINP.n175 4.5005
R46296 VINP.n350 VINP.n175 4.5005
R46297 VINP.n240 VINP.n175 4.5005
R46298 VINP.n352 VINP.n175 4.5005
R46299 VINP.n239 VINP.n175 4.5005
R46300 VINP.n354 VINP.n175 4.5005
R46301 VINP.n238 VINP.n175 4.5005
R46302 VINP.n356 VINP.n175 4.5005
R46303 VINP.n237 VINP.n175 4.5005
R46304 VINP.n358 VINP.n175 4.5005
R46305 VINP.n236 VINP.n175 4.5005
R46306 VINP.n360 VINP.n175 4.5005
R46307 VINP.n235 VINP.n175 4.5005
R46308 VINP.n362 VINP.n175 4.5005
R46309 VINP.n234 VINP.n175 4.5005
R46310 VINP.n364 VINP.n175 4.5005
R46311 VINP.n233 VINP.n175 4.5005
R46312 VINP.n366 VINP.n175 4.5005
R46313 VINP.n232 VINP.n175 4.5005
R46314 VINP.n368 VINP.n175 4.5005
R46315 VINP.n231 VINP.n175 4.5005
R46316 VINP.n370 VINP.n175 4.5005
R46317 VINP.n230 VINP.n175 4.5005
R46318 VINP.n372 VINP.n175 4.5005
R46319 VINP.n229 VINP.n175 4.5005
R46320 VINP.n374 VINP.n175 4.5005
R46321 VINP.n228 VINP.n175 4.5005
R46322 VINP.n376 VINP.n175 4.5005
R46323 VINP.n227 VINP.n175 4.5005
R46324 VINP.n378 VINP.n175 4.5005
R46325 VINP.n226 VINP.n175 4.5005
R46326 VINP.n380 VINP.n175 4.5005
R46327 VINP.n225 VINP.n175 4.5005
R46328 VINP.n382 VINP.n175 4.5005
R46329 VINP.n224 VINP.n175 4.5005
R46330 VINP.n384 VINP.n175 4.5005
R46331 VINP.n223 VINP.n175 4.5005
R46332 VINP.n386 VINP.n175 4.5005
R46333 VINP.n222 VINP.n175 4.5005
R46334 VINP.n388 VINP.n175 4.5005
R46335 VINP.n221 VINP.n175 4.5005
R46336 VINP.n390 VINP.n175 4.5005
R46337 VINP.n220 VINP.n175 4.5005
R46338 VINP.n392 VINP.n175 4.5005
R46339 VINP.n219 VINP.n175 4.5005
R46340 VINP.n394 VINP.n175 4.5005
R46341 VINP.n218 VINP.n175 4.5005
R46342 VINP.n396 VINP.n175 4.5005
R46343 VINP.n217 VINP.n175 4.5005
R46344 VINP.n398 VINP.n175 4.5005
R46345 VINP.n216 VINP.n175 4.5005
R46346 VINP.n400 VINP.n175 4.5005
R46347 VINP.n215 VINP.n175 4.5005
R46348 VINP.n654 VINP.n175 4.5005
R46349 VINP.n656 VINP.n175 4.5005
R46350 VINP.n175 VINP.n0 4.5005
R46351 VINP.n278 VINP.n125 4.5005
R46352 VINP.n276 VINP.n125 4.5005
R46353 VINP.n280 VINP.n125 4.5005
R46354 VINP.n275 VINP.n125 4.5005
R46355 VINP.n282 VINP.n125 4.5005
R46356 VINP.n274 VINP.n125 4.5005
R46357 VINP.n284 VINP.n125 4.5005
R46358 VINP.n273 VINP.n125 4.5005
R46359 VINP.n286 VINP.n125 4.5005
R46360 VINP.n272 VINP.n125 4.5005
R46361 VINP.n288 VINP.n125 4.5005
R46362 VINP.n271 VINP.n125 4.5005
R46363 VINP.n290 VINP.n125 4.5005
R46364 VINP.n270 VINP.n125 4.5005
R46365 VINP.n292 VINP.n125 4.5005
R46366 VINP.n269 VINP.n125 4.5005
R46367 VINP.n294 VINP.n125 4.5005
R46368 VINP.n268 VINP.n125 4.5005
R46369 VINP.n296 VINP.n125 4.5005
R46370 VINP.n267 VINP.n125 4.5005
R46371 VINP.n298 VINP.n125 4.5005
R46372 VINP.n266 VINP.n125 4.5005
R46373 VINP.n300 VINP.n125 4.5005
R46374 VINP.n265 VINP.n125 4.5005
R46375 VINP.n302 VINP.n125 4.5005
R46376 VINP.n264 VINP.n125 4.5005
R46377 VINP.n304 VINP.n125 4.5005
R46378 VINP.n263 VINP.n125 4.5005
R46379 VINP.n306 VINP.n125 4.5005
R46380 VINP.n262 VINP.n125 4.5005
R46381 VINP.n308 VINP.n125 4.5005
R46382 VINP.n261 VINP.n125 4.5005
R46383 VINP.n310 VINP.n125 4.5005
R46384 VINP.n260 VINP.n125 4.5005
R46385 VINP.n312 VINP.n125 4.5005
R46386 VINP.n259 VINP.n125 4.5005
R46387 VINP.n314 VINP.n125 4.5005
R46388 VINP.n258 VINP.n125 4.5005
R46389 VINP.n316 VINP.n125 4.5005
R46390 VINP.n257 VINP.n125 4.5005
R46391 VINP.n318 VINP.n125 4.5005
R46392 VINP.n256 VINP.n125 4.5005
R46393 VINP.n320 VINP.n125 4.5005
R46394 VINP.n255 VINP.n125 4.5005
R46395 VINP.n322 VINP.n125 4.5005
R46396 VINP.n254 VINP.n125 4.5005
R46397 VINP.n324 VINP.n125 4.5005
R46398 VINP.n253 VINP.n125 4.5005
R46399 VINP.n326 VINP.n125 4.5005
R46400 VINP.n252 VINP.n125 4.5005
R46401 VINP.n328 VINP.n125 4.5005
R46402 VINP.n251 VINP.n125 4.5005
R46403 VINP.n330 VINP.n125 4.5005
R46404 VINP.n250 VINP.n125 4.5005
R46405 VINP.n332 VINP.n125 4.5005
R46406 VINP.n249 VINP.n125 4.5005
R46407 VINP.n334 VINP.n125 4.5005
R46408 VINP.n248 VINP.n125 4.5005
R46409 VINP.n336 VINP.n125 4.5005
R46410 VINP.n247 VINP.n125 4.5005
R46411 VINP.n338 VINP.n125 4.5005
R46412 VINP.n246 VINP.n125 4.5005
R46413 VINP.n340 VINP.n125 4.5005
R46414 VINP.n245 VINP.n125 4.5005
R46415 VINP.n342 VINP.n125 4.5005
R46416 VINP.n244 VINP.n125 4.5005
R46417 VINP.n344 VINP.n125 4.5005
R46418 VINP.n243 VINP.n125 4.5005
R46419 VINP.n346 VINP.n125 4.5005
R46420 VINP.n242 VINP.n125 4.5005
R46421 VINP.n348 VINP.n125 4.5005
R46422 VINP.n241 VINP.n125 4.5005
R46423 VINP.n350 VINP.n125 4.5005
R46424 VINP.n240 VINP.n125 4.5005
R46425 VINP.n352 VINP.n125 4.5005
R46426 VINP.n239 VINP.n125 4.5005
R46427 VINP.n354 VINP.n125 4.5005
R46428 VINP.n238 VINP.n125 4.5005
R46429 VINP.n356 VINP.n125 4.5005
R46430 VINP.n237 VINP.n125 4.5005
R46431 VINP.n358 VINP.n125 4.5005
R46432 VINP.n236 VINP.n125 4.5005
R46433 VINP.n360 VINP.n125 4.5005
R46434 VINP.n235 VINP.n125 4.5005
R46435 VINP.n362 VINP.n125 4.5005
R46436 VINP.n234 VINP.n125 4.5005
R46437 VINP.n364 VINP.n125 4.5005
R46438 VINP.n233 VINP.n125 4.5005
R46439 VINP.n366 VINP.n125 4.5005
R46440 VINP.n232 VINP.n125 4.5005
R46441 VINP.n368 VINP.n125 4.5005
R46442 VINP.n231 VINP.n125 4.5005
R46443 VINP.n370 VINP.n125 4.5005
R46444 VINP.n230 VINP.n125 4.5005
R46445 VINP.n372 VINP.n125 4.5005
R46446 VINP.n229 VINP.n125 4.5005
R46447 VINP.n374 VINP.n125 4.5005
R46448 VINP.n228 VINP.n125 4.5005
R46449 VINP.n376 VINP.n125 4.5005
R46450 VINP.n227 VINP.n125 4.5005
R46451 VINP.n378 VINP.n125 4.5005
R46452 VINP.n226 VINP.n125 4.5005
R46453 VINP.n380 VINP.n125 4.5005
R46454 VINP.n225 VINP.n125 4.5005
R46455 VINP.n382 VINP.n125 4.5005
R46456 VINP.n224 VINP.n125 4.5005
R46457 VINP.n384 VINP.n125 4.5005
R46458 VINP.n223 VINP.n125 4.5005
R46459 VINP.n386 VINP.n125 4.5005
R46460 VINP.n222 VINP.n125 4.5005
R46461 VINP.n388 VINP.n125 4.5005
R46462 VINP.n221 VINP.n125 4.5005
R46463 VINP.n390 VINP.n125 4.5005
R46464 VINP.n220 VINP.n125 4.5005
R46465 VINP.n392 VINP.n125 4.5005
R46466 VINP.n219 VINP.n125 4.5005
R46467 VINP.n394 VINP.n125 4.5005
R46468 VINP.n218 VINP.n125 4.5005
R46469 VINP.n396 VINP.n125 4.5005
R46470 VINP.n217 VINP.n125 4.5005
R46471 VINP.n398 VINP.n125 4.5005
R46472 VINP.n216 VINP.n125 4.5005
R46473 VINP.n400 VINP.n125 4.5005
R46474 VINP.n215 VINP.n125 4.5005
R46475 VINP.n654 VINP.n125 4.5005
R46476 VINP.n656 VINP.n125 4.5005
R46477 VINP.n125 VINP.n0 4.5005
R46478 VINP.n278 VINP.n176 4.5005
R46479 VINP.n276 VINP.n176 4.5005
R46480 VINP.n280 VINP.n176 4.5005
R46481 VINP.n275 VINP.n176 4.5005
R46482 VINP.n282 VINP.n176 4.5005
R46483 VINP.n274 VINP.n176 4.5005
R46484 VINP.n284 VINP.n176 4.5005
R46485 VINP.n273 VINP.n176 4.5005
R46486 VINP.n286 VINP.n176 4.5005
R46487 VINP.n272 VINP.n176 4.5005
R46488 VINP.n288 VINP.n176 4.5005
R46489 VINP.n271 VINP.n176 4.5005
R46490 VINP.n290 VINP.n176 4.5005
R46491 VINP.n270 VINP.n176 4.5005
R46492 VINP.n292 VINP.n176 4.5005
R46493 VINP.n269 VINP.n176 4.5005
R46494 VINP.n294 VINP.n176 4.5005
R46495 VINP.n268 VINP.n176 4.5005
R46496 VINP.n296 VINP.n176 4.5005
R46497 VINP.n267 VINP.n176 4.5005
R46498 VINP.n298 VINP.n176 4.5005
R46499 VINP.n266 VINP.n176 4.5005
R46500 VINP.n300 VINP.n176 4.5005
R46501 VINP.n265 VINP.n176 4.5005
R46502 VINP.n302 VINP.n176 4.5005
R46503 VINP.n264 VINP.n176 4.5005
R46504 VINP.n304 VINP.n176 4.5005
R46505 VINP.n263 VINP.n176 4.5005
R46506 VINP.n306 VINP.n176 4.5005
R46507 VINP.n262 VINP.n176 4.5005
R46508 VINP.n308 VINP.n176 4.5005
R46509 VINP.n261 VINP.n176 4.5005
R46510 VINP.n310 VINP.n176 4.5005
R46511 VINP.n260 VINP.n176 4.5005
R46512 VINP.n312 VINP.n176 4.5005
R46513 VINP.n259 VINP.n176 4.5005
R46514 VINP.n314 VINP.n176 4.5005
R46515 VINP.n258 VINP.n176 4.5005
R46516 VINP.n316 VINP.n176 4.5005
R46517 VINP.n257 VINP.n176 4.5005
R46518 VINP.n318 VINP.n176 4.5005
R46519 VINP.n256 VINP.n176 4.5005
R46520 VINP.n320 VINP.n176 4.5005
R46521 VINP.n255 VINP.n176 4.5005
R46522 VINP.n322 VINP.n176 4.5005
R46523 VINP.n254 VINP.n176 4.5005
R46524 VINP.n324 VINP.n176 4.5005
R46525 VINP.n253 VINP.n176 4.5005
R46526 VINP.n326 VINP.n176 4.5005
R46527 VINP.n252 VINP.n176 4.5005
R46528 VINP.n328 VINP.n176 4.5005
R46529 VINP.n251 VINP.n176 4.5005
R46530 VINP.n330 VINP.n176 4.5005
R46531 VINP.n250 VINP.n176 4.5005
R46532 VINP.n332 VINP.n176 4.5005
R46533 VINP.n249 VINP.n176 4.5005
R46534 VINP.n334 VINP.n176 4.5005
R46535 VINP.n248 VINP.n176 4.5005
R46536 VINP.n336 VINP.n176 4.5005
R46537 VINP.n247 VINP.n176 4.5005
R46538 VINP.n338 VINP.n176 4.5005
R46539 VINP.n246 VINP.n176 4.5005
R46540 VINP.n340 VINP.n176 4.5005
R46541 VINP.n245 VINP.n176 4.5005
R46542 VINP.n342 VINP.n176 4.5005
R46543 VINP.n244 VINP.n176 4.5005
R46544 VINP.n344 VINP.n176 4.5005
R46545 VINP.n243 VINP.n176 4.5005
R46546 VINP.n346 VINP.n176 4.5005
R46547 VINP.n242 VINP.n176 4.5005
R46548 VINP.n348 VINP.n176 4.5005
R46549 VINP.n241 VINP.n176 4.5005
R46550 VINP.n350 VINP.n176 4.5005
R46551 VINP.n240 VINP.n176 4.5005
R46552 VINP.n352 VINP.n176 4.5005
R46553 VINP.n239 VINP.n176 4.5005
R46554 VINP.n354 VINP.n176 4.5005
R46555 VINP.n238 VINP.n176 4.5005
R46556 VINP.n356 VINP.n176 4.5005
R46557 VINP.n237 VINP.n176 4.5005
R46558 VINP.n358 VINP.n176 4.5005
R46559 VINP.n236 VINP.n176 4.5005
R46560 VINP.n360 VINP.n176 4.5005
R46561 VINP.n235 VINP.n176 4.5005
R46562 VINP.n362 VINP.n176 4.5005
R46563 VINP.n234 VINP.n176 4.5005
R46564 VINP.n364 VINP.n176 4.5005
R46565 VINP.n233 VINP.n176 4.5005
R46566 VINP.n366 VINP.n176 4.5005
R46567 VINP.n232 VINP.n176 4.5005
R46568 VINP.n368 VINP.n176 4.5005
R46569 VINP.n231 VINP.n176 4.5005
R46570 VINP.n370 VINP.n176 4.5005
R46571 VINP.n230 VINP.n176 4.5005
R46572 VINP.n372 VINP.n176 4.5005
R46573 VINP.n229 VINP.n176 4.5005
R46574 VINP.n374 VINP.n176 4.5005
R46575 VINP.n228 VINP.n176 4.5005
R46576 VINP.n376 VINP.n176 4.5005
R46577 VINP.n227 VINP.n176 4.5005
R46578 VINP.n378 VINP.n176 4.5005
R46579 VINP.n226 VINP.n176 4.5005
R46580 VINP.n380 VINP.n176 4.5005
R46581 VINP.n225 VINP.n176 4.5005
R46582 VINP.n382 VINP.n176 4.5005
R46583 VINP.n224 VINP.n176 4.5005
R46584 VINP.n384 VINP.n176 4.5005
R46585 VINP.n223 VINP.n176 4.5005
R46586 VINP.n386 VINP.n176 4.5005
R46587 VINP.n222 VINP.n176 4.5005
R46588 VINP.n388 VINP.n176 4.5005
R46589 VINP.n221 VINP.n176 4.5005
R46590 VINP.n390 VINP.n176 4.5005
R46591 VINP.n220 VINP.n176 4.5005
R46592 VINP.n392 VINP.n176 4.5005
R46593 VINP.n219 VINP.n176 4.5005
R46594 VINP.n394 VINP.n176 4.5005
R46595 VINP.n218 VINP.n176 4.5005
R46596 VINP.n396 VINP.n176 4.5005
R46597 VINP.n217 VINP.n176 4.5005
R46598 VINP.n398 VINP.n176 4.5005
R46599 VINP.n216 VINP.n176 4.5005
R46600 VINP.n400 VINP.n176 4.5005
R46601 VINP.n215 VINP.n176 4.5005
R46602 VINP.n654 VINP.n176 4.5005
R46603 VINP.n656 VINP.n176 4.5005
R46604 VINP.n176 VINP.n0 4.5005
R46605 VINP.n278 VINP.n124 4.5005
R46606 VINP.n276 VINP.n124 4.5005
R46607 VINP.n280 VINP.n124 4.5005
R46608 VINP.n275 VINP.n124 4.5005
R46609 VINP.n282 VINP.n124 4.5005
R46610 VINP.n274 VINP.n124 4.5005
R46611 VINP.n284 VINP.n124 4.5005
R46612 VINP.n273 VINP.n124 4.5005
R46613 VINP.n286 VINP.n124 4.5005
R46614 VINP.n272 VINP.n124 4.5005
R46615 VINP.n288 VINP.n124 4.5005
R46616 VINP.n271 VINP.n124 4.5005
R46617 VINP.n290 VINP.n124 4.5005
R46618 VINP.n270 VINP.n124 4.5005
R46619 VINP.n292 VINP.n124 4.5005
R46620 VINP.n269 VINP.n124 4.5005
R46621 VINP.n294 VINP.n124 4.5005
R46622 VINP.n268 VINP.n124 4.5005
R46623 VINP.n296 VINP.n124 4.5005
R46624 VINP.n267 VINP.n124 4.5005
R46625 VINP.n298 VINP.n124 4.5005
R46626 VINP.n266 VINP.n124 4.5005
R46627 VINP.n300 VINP.n124 4.5005
R46628 VINP.n265 VINP.n124 4.5005
R46629 VINP.n302 VINP.n124 4.5005
R46630 VINP.n264 VINP.n124 4.5005
R46631 VINP.n304 VINP.n124 4.5005
R46632 VINP.n263 VINP.n124 4.5005
R46633 VINP.n306 VINP.n124 4.5005
R46634 VINP.n262 VINP.n124 4.5005
R46635 VINP.n308 VINP.n124 4.5005
R46636 VINP.n261 VINP.n124 4.5005
R46637 VINP.n310 VINP.n124 4.5005
R46638 VINP.n260 VINP.n124 4.5005
R46639 VINP.n312 VINP.n124 4.5005
R46640 VINP.n259 VINP.n124 4.5005
R46641 VINP.n314 VINP.n124 4.5005
R46642 VINP.n258 VINP.n124 4.5005
R46643 VINP.n316 VINP.n124 4.5005
R46644 VINP.n257 VINP.n124 4.5005
R46645 VINP.n318 VINP.n124 4.5005
R46646 VINP.n256 VINP.n124 4.5005
R46647 VINP.n320 VINP.n124 4.5005
R46648 VINP.n255 VINP.n124 4.5005
R46649 VINP.n322 VINP.n124 4.5005
R46650 VINP.n254 VINP.n124 4.5005
R46651 VINP.n324 VINP.n124 4.5005
R46652 VINP.n253 VINP.n124 4.5005
R46653 VINP.n326 VINP.n124 4.5005
R46654 VINP.n252 VINP.n124 4.5005
R46655 VINP.n328 VINP.n124 4.5005
R46656 VINP.n251 VINP.n124 4.5005
R46657 VINP.n330 VINP.n124 4.5005
R46658 VINP.n250 VINP.n124 4.5005
R46659 VINP.n332 VINP.n124 4.5005
R46660 VINP.n249 VINP.n124 4.5005
R46661 VINP.n334 VINP.n124 4.5005
R46662 VINP.n248 VINP.n124 4.5005
R46663 VINP.n336 VINP.n124 4.5005
R46664 VINP.n247 VINP.n124 4.5005
R46665 VINP.n338 VINP.n124 4.5005
R46666 VINP.n246 VINP.n124 4.5005
R46667 VINP.n340 VINP.n124 4.5005
R46668 VINP.n245 VINP.n124 4.5005
R46669 VINP.n342 VINP.n124 4.5005
R46670 VINP.n244 VINP.n124 4.5005
R46671 VINP.n344 VINP.n124 4.5005
R46672 VINP.n243 VINP.n124 4.5005
R46673 VINP.n346 VINP.n124 4.5005
R46674 VINP.n242 VINP.n124 4.5005
R46675 VINP.n348 VINP.n124 4.5005
R46676 VINP.n241 VINP.n124 4.5005
R46677 VINP.n350 VINP.n124 4.5005
R46678 VINP.n240 VINP.n124 4.5005
R46679 VINP.n352 VINP.n124 4.5005
R46680 VINP.n239 VINP.n124 4.5005
R46681 VINP.n354 VINP.n124 4.5005
R46682 VINP.n238 VINP.n124 4.5005
R46683 VINP.n356 VINP.n124 4.5005
R46684 VINP.n237 VINP.n124 4.5005
R46685 VINP.n358 VINP.n124 4.5005
R46686 VINP.n236 VINP.n124 4.5005
R46687 VINP.n360 VINP.n124 4.5005
R46688 VINP.n235 VINP.n124 4.5005
R46689 VINP.n362 VINP.n124 4.5005
R46690 VINP.n234 VINP.n124 4.5005
R46691 VINP.n364 VINP.n124 4.5005
R46692 VINP.n233 VINP.n124 4.5005
R46693 VINP.n366 VINP.n124 4.5005
R46694 VINP.n232 VINP.n124 4.5005
R46695 VINP.n368 VINP.n124 4.5005
R46696 VINP.n231 VINP.n124 4.5005
R46697 VINP.n370 VINP.n124 4.5005
R46698 VINP.n230 VINP.n124 4.5005
R46699 VINP.n372 VINP.n124 4.5005
R46700 VINP.n229 VINP.n124 4.5005
R46701 VINP.n374 VINP.n124 4.5005
R46702 VINP.n228 VINP.n124 4.5005
R46703 VINP.n376 VINP.n124 4.5005
R46704 VINP.n227 VINP.n124 4.5005
R46705 VINP.n378 VINP.n124 4.5005
R46706 VINP.n226 VINP.n124 4.5005
R46707 VINP.n380 VINP.n124 4.5005
R46708 VINP.n225 VINP.n124 4.5005
R46709 VINP.n382 VINP.n124 4.5005
R46710 VINP.n224 VINP.n124 4.5005
R46711 VINP.n384 VINP.n124 4.5005
R46712 VINP.n223 VINP.n124 4.5005
R46713 VINP.n386 VINP.n124 4.5005
R46714 VINP.n222 VINP.n124 4.5005
R46715 VINP.n388 VINP.n124 4.5005
R46716 VINP.n221 VINP.n124 4.5005
R46717 VINP.n390 VINP.n124 4.5005
R46718 VINP.n220 VINP.n124 4.5005
R46719 VINP.n392 VINP.n124 4.5005
R46720 VINP.n219 VINP.n124 4.5005
R46721 VINP.n394 VINP.n124 4.5005
R46722 VINP.n218 VINP.n124 4.5005
R46723 VINP.n396 VINP.n124 4.5005
R46724 VINP.n217 VINP.n124 4.5005
R46725 VINP.n398 VINP.n124 4.5005
R46726 VINP.n216 VINP.n124 4.5005
R46727 VINP.n400 VINP.n124 4.5005
R46728 VINP.n215 VINP.n124 4.5005
R46729 VINP.n654 VINP.n124 4.5005
R46730 VINP.n656 VINP.n124 4.5005
R46731 VINP.n124 VINP.n0 4.5005
R46732 VINP.n278 VINP.n177 4.5005
R46733 VINP.n276 VINP.n177 4.5005
R46734 VINP.n280 VINP.n177 4.5005
R46735 VINP.n275 VINP.n177 4.5005
R46736 VINP.n282 VINP.n177 4.5005
R46737 VINP.n274 VINP.n177 4.5005
R46738 VINP.n284 VINP.n177 4.5005
R46739 VINP.n273 VINP.n177 4.5005
R46740 VINP.n286 VINP.n177 4.5005
R46741 VINP.n272 VINP.n177 4.5005
R46742 VINP.n288 VINP.n177 4.5005
R46743 VINP.n271 VINP.n177 4.5005
R46744 VINP.n290 VINP.n177 4.5005
R46745 VINP.n270 VINP.n177 4.5005
R46746 VINP.n292 VINP.n177 4.5005
R46747 VINP.n269 VINP.n177 4.5005
R46748 VINP.n294 VINP.n177 4.5005
R46749 VINP.n268 VINP.n177 4.5005
R46750 VINP.n296 VINP.n177 4.5005
R46751 VINP.n267 VINP.n177 4.5005
R46752 VINP.n298 VINP.n177 4.5005
R46753 VINP.n266 VINP.n177 4.5005
R46754 VINP.n300 VINP.n177 4.5005
R46755 VINP.n265 VINP.n177 4.5005
R46756 VINP.n302 VINP.n177 4.5005
R46757 VINP.n264 VINP.n177 4.5005
R46758 VINP.n304 VINP.n177 4.5005
R46759 VINP.n263 VINP.n177 4.5005
R46760 VINP.n306 VINP.n177 4.5005
R46761 VINP.n262 VINP.n177 4.5005
R46762 VINP.n308 VINP.n177 4.5005
R46763 VINP.n261 VINP.n177 4.5005
R46764 VINP.n310 VINP.n177 4.5005
R46765 VINP.n260 VINP.n177 4.5005
R46766 VINP.n312 VINP.n177 4.5005
R46767 VINP.n259 VINP.n177 4.5005
R46768 VINP.n314 VINP.n177 4.5005
R46769 VINP.n258 VINP.n177 4.5005
R46770 VINP.n316 VINP.n177 4.5005
R46771 VINP.n257 VINP.n177 4.5005
R46772 VINP.n318 VINP.n177 4.5005
R46773 VINP.n256 VINP.n177 4.5005
R46774 VINP.n320 VINP.n177 4.5005
R46775 VINP.n255 VINP.n177 4.5005
R46776 VINP.n322 VINP.n177 4.5005
R46777 VINP.n254 VINP.n177 4.5005
R46778 VINP.n324 VINP.n177 4.5005
R46779 VINP.n253 VINP.n177 4.5005
R46780 VINP.n326 VINP.n177 4.5005
R46781 VINP.n252 VINP.n177 4.5005
R46782 VINP.n328 VINP.n177 4.5005
R46783 VINP.n251 VINP.n177 4.5005
R46784 VINP.n330 VINP.n177 4.5005
R46785 VINP.n250 VINP.n177 4.5005
R46786 VINP.n332 VINP.n177 4.5005
R46787 VINP.n249 VINP.n177 4.5005
R46788 VINP.n334 VINP.n177 4.5005
R46789 VINP.n248 VINP.n177 4.5005
R46790 VINP.n336 VINP.n177 4.5005
R46791 VINP.n247 VINP.n177 4.5005
R46792 VINP.n338 VINP.n177 4.5005
R46793 VINP.n246 VINP.n177 4.5005
R46794 VINP.n340 VINP.n177 4.5005
R46795 VINP.n245 VINP.n177 4.5005
R46796 VINP.n342 VINP.n177 4.5005
R46797 VINP.n244 VINP.n177 4.5005
R46798 VINP.n344 VINP.n177 4.5005
R46799 VINP.n243 VINP.n177 4.5005
R46800 VINP.n346 VINP.n177 4.5005
R46801 VINP.n242 VINP.n177 4.5005
R46802 VINP.n348 VINP.n177 4.5005
R46803 VINP.n241 VINP.n177 4.5005
R46804 VINP.n350 VINP.n177 4.5005
R46805 VINP.n240 VINP.n177 4.5005
R46806 VINP.n352 VINP.n177 4.5005
R46807 VINP.n239 VINP.n177 4.5005
R46808 VINP.n354 VINP.n177 4.5005
R46809 VINP.n238 VINP.n177 4.5005
R46810 VINP.n356 VINP.n177 4.5005
R46811 VINP.n237 VINP.n177 4.5005
R46812 VINP.n358 VINP.n177 4.5005
R46813 VINP.n236 VINP.n177 4.5005
R46814 VINP.n360 VINP.n177 4.5005
R46815 VINP.n235 VINP.n177 4.5005
R46816 VINP.n362 VINP.n177 4.5005
R46817 VINP.n234 VINP.n177 4.5005
R46818 VINP.n364 VINP.n177 4.5005
R46819 VINP.n233 VINP.n177 4.5005
R46820 VINP.n366 VINP.n177 4.5005
R46821 VINP.n232 VINP.n177 4.5005
R46822 VINP.n368 VINP.n177 4.5005
R46823 VINP.n231 VINP.n177 4.5005
R46824 VINP.n370 VINP.n177 4.5005
R46825 VINP.n230 VINP.n177 4.5005
R46826 VINP.n372 VINP.n177 4.5005
R46827 VINP.n229 VINP.n177 4.5005
R46828 VINP.n374 VINP.n177 4.5005
R46829 VINP.n228 VINP.n177 4.5005
R46830 VINP.n376 VINP.n177 4.5005
R46831 VINP.n227 VINP.n177 4.5005
R46832 VINP.n378 VINP.n177 4.5005
R46833 VINP.n226 VINP.n177 4.5005
R46834 VINP.n380 VINP.n177 4.5005
R46835 VINP.n225 VINP.n177 4.5005
R46836 VINP.n382 VINP.n177 4.5005
R46837 VINP.n224 VINP.n177 4.5005
R46838 VINP.n384 VINP.n177 4.5005
R46839 VINP.n223 VINP.n177 4.5005
R46840 VINP.n386 VINP.n177 4.5005
R46841 VINP.n222 VINP.n177 4.5005
R46842 VINP.n388 VINP.n177 4.5005
R46843 VINP.n221 VINP.n177 4.5005
R46844 VINP.n390 VINP.n177 4.5005
R46845 VINP.n220 VINP.n177 4.5005
R46846 VINP.n392 VINP.n177 4.5005
R46847 VINP.n219 VINP.n177 4.5005
R46848 VINP.n394 VINP.n177 4.5005
R46849 VINP.n218 VINP.n177 4.5005
R46850 VINP.n396 VINP.n177 4.5005
R46851 VINP.n217 VINP.n177 4.5005
R46852 VINP.n398 VINP.n177 4.5005
R46853 VINP.n216 VINP.n177 4.5005
R46854 VINP.n400 VINP.n177 4.5005
R46855 VINP.n215 VINP.n177 4.5005
R46856 VINP.n654 VINP.n177 4.5005
R46857 VINP.n656 VINP.n177 4.5005
R46858 VINP.n177 VINP.n0 4.5005
R46859 VINP.n278 VINP.n123 4.5005
R46860 VINP.n276 VINP.n123 4.5005
R46861 VINP.n280 VINP.n123 4.5005
R46862 VINP.n275 VINP.n123 4.5005
R46863 VINP.n282 VINP.n123 4.5005
R46864 VINP.n274 VINP.n123 4.5005
R46865 VINP.n284 VINP.n123 4.5005
R46866 VINP.n273 VINP.n123 4.5005
R46867 VINP.n286 VINP.n123 4.5005
R46868 VINP.n272 VINP.n123 4.5005
R46869 VINP.n288 VINP.n123 4.5005
R46870 VINP.n271 VINP.n123 4.5005
R46871 VINP.n290 VINP.n123 4.5005
R46872 VINP.n270 VINP.n123 4.5005
R46873 VINP.n292 VINP.n123 4.5005
R46874 VINP.n269 VINP.n123 4.5005
R46875 VINP.n294 VINP.n123 4.5005
R46876 VINP.n268 VINP.n123 4.5005
R46877 VINP.n296 VINP.n123 4.5005
R46878 VINP.n267 VINP.n123 4.5005
R46879 VINP.n298 VINP.n123 4.5005
R46880 VINP.n266 VINP.n123 4.5005
R46881 VINP.n300 VINP.n123 4.5005
R46882 VINP.n265 VINP.n123 4.5005
R46883 VINP.n302 VINP.n123 4.5005
R46884 VINP.n264 VINP.n123 4.5005
R46885 VINP.n304 VINP.n123 4.5005
R46886 VINP.n263 VINP.n123 4.5005
R46887 VINP.n306 VINP.n123 4.5005
R46888 VINP.n262 VINP.n123 4.5005
R46889 VINP.n308 VINP.n123 4.5005
R46890 VINP.n261 VINP.n123 4.5005
R46891 VINP.n310 VINP.n123 4.5005
R46892 VINP.n260 VINP.n123 4.5005
R46893 VINP.n312 VINP.n123 4.5005
R46894 VINP.n259 VINP.n123 4.5005
R46895 VINP.n314 VINP.n123 4.5005
R46896 VINP.n258 VINP.n123 4.5005
R46897 VINP.n316 VINP.n123 4.5005
R46898 VINP.n257 VINP.n123 4.5005
R46899 VINP.n318 VINP.n123 4.5005
R46900 VINP.n256 VINP.n123 4.5005
R46901 VINP.n320 VINP.n123 4.5005
R46902 VINP.n255 VINP.n123 4.5005
R46903 VINP.n322 VINP.n123 4.5005
R46904 VINP.n254 VINP.n123 4.5005
R46905 VINP.n324 VINP.n123 4.5005
R46906 VINP.n253 VINP.n123 4.5005
R46907 VINP.n326 VINP.n123 4.5005
R46908 VINP.n252 VINP.n123 4.5005
R46909 VINP.n328 VINP.n123 4.5005
R46910 VINP.n251 VINP.n123 4.5005
R46911 VINP.n330 VINP.n123 4.5005
R46912 VINP.n250 VINP.n123 4.5005
R46913 VINP.n332 VINP.n123 4.5005
R46914 VINP.n249 VINP.n123 4.5005
R46915 VINP.n334 VINP.n123 4.5005
R46916 VINP.n248 VINP.n123 4.5005
R46917 VINP.n336 VINP.n123 4.5005
R46918 VINP.n247 VINP.n123 4.5005
R46919 VINP.n338 VINP.n123 4.5005
R46920 VINP.n246 VINP.n123 4.5005
R46921 VINP.n340 VINP.n123 4.5005
R46922 VINP.n245 VINP.n123 4.5005
R46923 VINP.n342 VINP.n123 4.5005
R46924 VINP.n244 VINP.n123 4.5005
R46925 VINP.n344 VINP.n123 4.5005
R46926 VINP.n243 VINP.n123 4.5005
R46927 VINP.n346 VINP.n123 4.5005
R46928 VINP.n242 VINP.n123 4.5005
R46929 VINP.n348 VINP.n123 4.5005
R46930 VINP.n241 VINP.n123 4.5005
R46931 VINP.n350 VINP.n123 4.5005
R46932 VINP.n240 VINP.n123 4.5005
R46933 VINP.n352 VINP.n123 4.5005
R46934 VINP.n239 VINP.n123 4.5005
R46935 VINP.n354 VINP.n123 4.5005
R46936 VINP.n238 VINP.n123 4.5005
R46937 VINP.n356 VINP.n123 4.5005
R46938 VINP.n237 VINP.n123 4.5005
R46939 VINP.n358 VINP.n123 4.5005
R46940 VINP.n236 VINP.n123 4.5005
R46941 VINP.n360 VINP.n123 4.5005
R46942 VINP.n235 VINP.n123 4.5005
R46943 VINP.n362 VINP.n123 4.5005
R46944 VINP.n234 VINP.n123 4.5005
R46945 VINP.n364 VINP.n123 4.5005
R46946 VINP.n233 VINP.n123 4.5005
R46947 VINP.n366 VINP.n123 4.5005
R46948 VINP.n232 VINP.n123 4.5005
R46949 VINP.n368 VINP.n123 4.5005
R46950 VINP.n231 VINP.n123 4.5005
R46951 VINP.n370 VINP.n123 4.5005
R46952 VINP.n230 VINP.n123 4.5005
R46953 VINP.n372 VINP.n123 4.5005
R46954 VINP.n229 VINP.n123 4.5005
R46955 VINP.n374 VINP.n123 4.5005
R46956 VINP.n228 VINP.n123 4.5005
R46957 VINP.n376 VINP.n123 4.5005
R46958 VINP.n227 VINP.n123 4.5005
R46959 VINP.n378 VINP.n123 4.5005
R46960 VINP.n226 VINP.n123 4.5005
R46961 VINP.n380 VINP.n123 4.5005
R46962 VINP.n225 VINP.n123 4.5005
R46963 VINP.n382 VINP.n123 4.5005
R46964 VINP.n224 VINP.n123 4.5005
R46965 VINP.n384 VINP.n123 4.5005
R46966 VINP.n223 VINP.n123 4.5005
R46967 VINP.n386 VINP.n123 4.5005
R46968 VINP.n222 VINP.n123 4.5005
R46969 VINP.n388 VINP.n123 4.5005
R46970 VINP.n221 VINP.n123 4.5005
R46971 VINP.n390 VINP.n123 4.5005
R46972 VINP.n220 VINP.n123 4.5005
R46973 VINP.n392 VINP.n123 4.5005
R46974 VINP.n219 VINP.n123 4.5005
R46975 VINP.n394 VINP.n123 4.5005
R46976 VINP.n218 VINP.n123 4.5005
R46977 VINP.n396 VINP.n123 4.5005
R46978 VINP.n217 VINP.n123 4.5005
R46979 VINP.n398 VINP.n123 4.5005
R46980 VINP.n216 VINP.n123 4.5005
R46981 VINP.n400 VINP.n123 4.5005
R46982 VINP.n215 VINP.n123 4.5005
R46983 VINP.n654 VINP.n123 4.5005
R46984 VINP.n656 VINP.n123 4.5005
R46985 VINP.n123 VINP.n0 4.5005
R46986 VINP.n278 VINP.n178 4.5005
R46987 VINP.n276 VINP.n178 4.5005
R46988 VINP.n280 VINP.n178 4.5005
R46989 VINP.n275 VINP.n178 4.5005
R46990 VINP.n282 VINP.n178 4.5005
R46991 VINP.n274 VINP.n178 4.5005
R46992 VINP.n284 VINP.n178 4.5005
R46993 VINP.n273 VINP.n178 4.5005
R46994 VINP.n286 VINP.n178 4.5005
R46995 VINP.n272 VINP.n178 4.5005
R46996 VINP.n288 VINP.n178 4.5005
R46997 VINP.n271 VINP.n178 4.5005
R46998 VINP.n290 VINP.n178 4.5005
R46999 VINP.n270 VINP.n178 4.5005
R47000 VINP.n292 VINP.n178 4.5005
R47001 VINP.n269 VINP.n178 4.5005
R47002 VINP.n294 VINP.n178 4.5005
R47003 VINP.n268 VINP.n178 4.5005
R47004 VINP.n296 VINP.n178 4.5005
R47005 VINP.n267 VINP.n178 4.5005
R47006 VINP.n298 VINP.n178 4.5005
R47007 VINP.n266 VINP.n178 4.5005
R47008 VINP.n300 VINP.n178 4.5005
R47009 VINP.n265 VINP.n178 4.5005
R47010 VINP.n302 VINP.n178 4.5005
R47011 VINP.n264 VINP.n178 4.5005
R47012 VINP.n304 VINP.n178 4.5005
R47013 VINP.n263 VINP.n178 4.5005
R47014 VINP.n306 VINP.n178 4.5005
R47015 VINP.n262 VINP.n178 4.5005
R47016 VINP.n308 VINP.n178 4.5005
R47017 VINP.n261 VINP.n178 4.5005
R47018 VINP.n310 VINP.n178 4.5005
R47019 VINP.n260 VINP.n178 4.5005
R47020 VINP.n312 VINP.n178 4.5005
R47021 VINP.n259 VINP.n178 4.5005
R47022 VINP.n314 VINP.n178 4.5005
R47023 VINP.n258 VINP.n178 4.5005
R47024 VINP.n316 VINP.n178 4.5005
R47025 VINP.n257 VINP.n178 4.5005
R47026 VINP.n318 VINP.n178 4.5005
R47027 VINP.n256 VINP.n178 4.5005
R47028 VINP.n320 VINP.n178 4.5005
R47029 VINP.n255 VINP.n178 4.5005
R47030 VINP.n322 VINP.n178 4.5005
R47031 VINP.n254 VINP.n178 4.5005
R47032 VINP.n324 VINP.n178 4.5005
R47033 VINP.n253 VINP.n178 4.5005
R47034 VINP.n326 VINP.n178 4.5005
R47035 VINP.n252 VINP.n178 4.5005
R47036 VINP.n328 VINP.n178 4.5005
R47037 VINP.n251 VINP.n178 4.5005
R47038 VINP.n330 VINP.n178 4.5005
R47039 VINP.n250 VINP.n178 4.5005
R47040 VINP.n332 VINP.n178 4.5005
R47041 VINP.n249 VINP.n178 4.5005
R47042 VINP.n334 VINP.n178 4.5005
R47043 VINP.n248 VINP.n178 4.5005
R47044 VINP.n336 VINP.n178 4.5005
R47045 VINP.n247 VINP.n178 4.5005
R47046 VINP.n338 VINP.n178 4.5005
R47047 VINP.n246 VINP.n178 4.5005
R47048 VINP.n340 VINP.n178 4.5005
R47049 VINP.n245 VINP.n178 4.5005
R47050 VINP.n342 VINP.n178 4.5005
R47051 VINP.n244 VINP.n178 4.5005
R47052 VINP.n344 VINP.n178 4.5005
R47053 VINP.n243 VINP.n178 4.5005
R47054 VINP.n346 VINP.n178 4.5005
R47055 VINP.n242 VINP.n178 4.5005
R47056 VINP.n348 VINP.n178 4.5005
R47057 VINP.n241 VINP.n178 4.5005
R47058 VINP.n350 VINP.n178 4.5005
R47059 VINP.n240 VINP.n178 4.5005
R47060 VINP.n352 VINP.n178 4.5005
R47061 VINP.n239 VINP.n178 4.5005
R47062 VINP.n354 VINP.n178 4.5005
R47063 VINP.n238 VINP.n178 4.5005
R47064 VINP.n356 VINP.n178 4.5005
R47065 VINP.n237 VINP.n178 4.5005
R47066 VINP.n358 VINP.n178 4.5005
R47067 VINP.n236 VINP.n178 4.5005
R47068 VINP.n360 VINP.n178 4.5005
R47069 VINP.n235 VINP.n178 4.5005
R47070 VINP.n362 VINP.n178 4.5005
R47071 VINP.n234 VINP.n178 4.5005
R47072 VINP.n364 VINP.n178 4.5005
R47073 VINP.n233 VINP.n178 4.5005
R47074 VINP.n366 VINP.n178 4.5005
R47075 VINP.n232 VINP.n178 4.5005
R47076 VINP.n368 VINP.n178 4.5005
R47077 VINP.n231 VINP.n178 4.5005
R47078 VINP.n370 VINP.n178 4.5005
R47079 VINP.n230 VINP.n178 4.5005
R47080 VINP.n372 VINP.n178 4.5005
R47081 VINP.n229 VINP.n178 4.5005
R47082 VINP.n374 VINP.n178 4.5005
R47083 VINP.n228 VINP.n178 4.5005
R47084 VINP.n376 VINP.n178 4.5005
R47085 VINP.n227 VINP.n178 4.5005
R47086 VINP.n378 VINP.n178 4.5005
R47087 VINP.n226 VINP.n178 4.5005
R47088 VINP.n380 VINP.n178 4.5005
R47089 VINP.n225 VINP.n178 4.5005
R47090 VINP.n382 VINP.n178 4.5005
R47091 VINP.n224 VINP.n178 4.5005
R47092 VINP.n384 VINP.n178 4.5005
R47093 VINP.n223 VINP.n178 4.5005
R47094 VINP.n386 VINP.n178 4.5005
R47095 VINP.n222 VINP.n178 4.5005
R47096 VINP.n388 VINP.n178 4.5005
R47097 VINP.n221 VINP.n178 4.5005
R47098 VINP.n390 VINP.n178 4.5005
R47099 VINP.n220 VINP.n178 4.5005
R47100 VINP.n392 VINP.n178 4.5005
R47101 VINP.n219 VINP.n178 4.5005
R47102 VINP.n394 VINP.n178 4.5005
R47103 VINP.n218 VINP.n178 4.5005
R47104 VINP.n396 VINP.n178 4.5005
R47105 VINP.n217 VINP.n178 4.5005
R47106 VINP.n398 VINP.n178 4.5005
R47107 VINP.n216 VINP.n178 4.5005
R47108 VINP.n400 VINP.n178 4.5005
R47109 VINP.n215 VINP.n178 4.5005
R47110 VINP.n654 VINP.n178 4.5005
R47111 VINP.n656 VINP.n178 4.5005
R47112 VINP.n178 VINP.n0 4.5005
R47113 VINP.n278 VINP.n122 4.5005
R47114 VINP.n276 VINP.n122 4.5005
R47115 VINP.n280 VINP.n122 4.5005
R47116 VINP.n275 VINP.n122 4.5005
R47117 VINP.n282 VINP.n122 4.5005
R47118 VINP.n274 VINP.n122 4.5005
R47119 VINP.n284 VINP.n122 4.5005
R47120 VINP.n273 VINP.n122 4.5005
R47121 VINP.n286 VINP.n122 4.5005
R47122 VINP.n272 VINP.n122 4.5005
R47123 VINP.n288 VINP.n122 4.5005
R47124 VINP.n271 VINP.n122 4.5005
R47125 VINP.n290 VINP.n122 4.5005
R47126 VINP.n270 VINP.n122 4.5005
R47127 VINP.n292 VINP.n122 4.5005
R47128 VINP.n269 VINP.n122 4.5005
R47129 VINP.n294 VINP.n122 4.5005
R47130 VINP.n268 VINP.n122 4.5005
R47131 VINP.n296 VINP.n122 4.5005
R47132 VINP.n267 VINP.n122 4.5005
R47133 VINP.n298 VINP.n122 4.5005
R47134 VINP.n266 VINP.n122 4.5005
R47135 VINP.n300 VINP.n122 4.5005
R47136 VINP.n265 VINP.n122 4.5005
R47137 VINP.n302 VINP.n122 4.5005
R47138 VINP.n264 VINP.n122 4.5005
R47139 VINP.n304 VINP.n122 4.5005
R47140 VINP.n263 VINP.n122 4.5005
R47141 VINP.n306 VINP.n122 4.5005
R47142 VINP.n262 VINP.n122 4.5005
R47143 VINP.n308 VINP.n122 4.5005
R47144 VINP.n261 VINP.n122 4.5005
R47145 VINP.n310 VINP.n122 4.5005
R47146 VINP.n260 VINP.n122 4.5005
R47147 VINP.n312 VINP.n122 4.5005
R47148 VINP.n259 VINP.n122 4.5005
R47149 VINP.n314 VINP.n122 4.5005
R47150 VINP.n258 VINP.n122 4.5005
R47151 VINP.n316 VINP.n122 4.5005
R47152 VINP.n257 VINP.n122 4.5005
R47153 VINP.n318 VINP.n122 4.5005
R47154 VINP.n256 VINP.n122 4.5005
R47155 VINP.n320 VINP.n122 4.5005
R47156 VINP.n255 VINP.n122 4.5005
R47157 VINP.n322 VINP.n122 4.5005
R47158 VINP.n254 VINP.n122 4.5005
R47159 VINP.n324 VINP.n122 4.5005
R47160 VINP.n253 VINP.n122 4.5005
R47161 VINP.n326 VINP.n122 4.5005
R47162 VINP.n252 VINP.n122 4.5005
R47163 VINP.n328 VINP.n122 4.5005
R47164 VINP.n251 VINP.n122 4.5005
R47165 VINP.n330 VINP.n122 4.5005
R47166 VINP.n250 VINP.n122 4.5005
R47167 VINP.n332 VINP.n122 4.5005
R47168 VINP.n249 VINP.n122 4.5005
R47169 VINP.n334 VINP.n122 4.5005
R47170 VINP.n248 VINP.n122 4.5005
R47171 VINP.n336 VINP.n122 4.5005
R47172 VINP.n247 VINP.n122 4.5005
R47173 VINP.n338 VINP.n122 4.5005
R47174 VINP.n246 VINP.n122 4.5005
R47175 VINP.n340 VINP.n122 4.5005
R47176 VINP.n245 VINP.n122 4.5005
R47177 VINP.n342 VINP.n122 4.5005
R47178 VINP.n244 VINP.n122 4.5005
R47179 VINP.n344 VINP.n122 4.5005
R47180 VINP.n243 VINP.n122 4.5005
R47181 VINP.n346 VINP.n122 4.5005
R47182 VINP.n242 VINP.n122 4.5005
R47183 VINP.n348 VINP.n122 4.5005
R47184 VINP.n241 VINP.n122 4.5005
R47185 VINP.n350 VINP.n122 4.5005
R47186 VINP.n240 VINP.n122 4.5005
R47187 VINP.n352 VINP.n122 4.5005
R47188 VINP.n239 VINP.n122 4.5005
R47189 VINP.n354 VINP.n122 4.5005
R47190 VINP.n238 VINP.n122 4.5005
R47191 VINP.n356 VINP.n122 4.5005
R47192 VINP.n237 VINP.n122 4.5005
R47193 VINP.n358 VINP.n122 4.5005
R47194 VINP.n236 VINP.n122 4.5005
R47195 VINP.n360 VINP.n122 4.5005
R47196 VINP.n235 VINP.n122 4.5005
R47197 VINP.n362 VINP.n122 4.5005
R47198 VINP.n234 VINP.n122 4.5005
R47199 VINP.n364 VINP.n122 4.5005
R47200 VINP.n233 VINP.n122 4.5005
R47201 VINP.n366 VINP.n122 4.5005
R47202 VINP.n232 VINP.n122 4.5005
R47203 VINP.n368 VINP.n122 4.5005
R47204 VINP.n231 VINP.n122 4.5005
R47205 VINP.n370 VINP.n122 4.5005
R47206 VINP.n230 VINP.n122 4.5005
R47207 VINP.n372 VINP.n122 4.5005
R47208 VINP.n229 VINP.n122 4.5005
R47209 VINP.n374 VINP.n122 4.5005
R47210 VINP.n228 VINP.n122 4.5005
R47211 VINP.n376 VINP.n122 4.5005
R47212 VINP.n227 VINP.n122 4.5005
R47213 VINP.n378 VINP.n122 4.5005
R47214 VINP.n226 VINP.n122 4.5005
R47215 VINP.n380 VINP.n122 4.5005
R47216 VINP.n225 VINP.n122 4.5005
R47217 VINP.n382 VINP.n122 4.5005
R47218 VINP.n224 VINP.n122 4.5005
R47219 VINP.n384 VINP.n122 4.5005
R47220 VINP.n223 VINP.n122 4.5005
R47221 VINP.n386 VINP.n122 4.5005
R47222 VINP.n222 VINP.n122 4.5005
R47223 VINP.n388 VINP.n122 4.5005
R47224 VINP.n221 VINP.n122 4.5005
R47225 VINP.n390 VINP.n122 4.5005
R47226 VINP.n220 VINP.n122 4.5005
R47227 VINP.n392 VINP.n122 4.5005
R47228 VINP.n219 VINP.n122 4.5005
R47229 VINP.n394 VINP.n122 4.5005
R47230 VINP.n218 VINP.n122 4.5005
R47231 VINP.n396 VINP.n122 4.5005
R47232 VINP.n217 VINP.n122 4.5005
R47233 VINP.n398 VINP.n122 4.5005
R47234 VINP.n216 VINP.n122 4.5005
R47235 VINP.n400 VINP.n122 4.5005
R47236 VINP.n215 VINP.n122 4.5005
R47237 VINP.n654 VINP.n122 4.5005
R47238 VINP.n656 VINP.n122 4.5005
R47239 VINP.n122 VINP.n0 4.5005
R47240 VINP.n278 VINP.n179 4.5005
R47241 VINP.n276 VINP.n179 4.5005
R47242 VINP.n280 VINP.n179 4.5005
R47243 VINP.n275 VINP.n179 4.5005
R47244 VINP.n282 VINP.n179 4.5005
R47245 VINP.n274 VINP.n179 4.5005
R47246 VINP.n284 VINP.n179 4.5005
R47247 VINP.n273 VINP.n179 4.5005
R47248 VINP.n286 VINP.n179 4.5005
R47249 VINP.n272 VINP.n179 4.5005
R47250 VINP.n288 VINP.n179 4.5005
R47251 VINP.n271 VINP.n179 4.5005
R47252 VINP.n290 VINP.n179 4.5005
R47253 VINP.n270 VINP.n179 4.5005
R47254 VINP.n292 VINP.n179 4.5005
R47255 VINP.n269 VINP.n179 4.5005
R47256 VINP.n294 VINP.n179 4.5005
R47257 VINP.n268 VINP.n179 4.5005
R47258 VINP.n296 VINP.n179 4.5005
R47259 VINP.n267 VINP.n179 4.5005
R47260 VINP.n298 VINP.n179 4.5005
R47261 VINP.n266 VINP.n179 4.5005
R47262 VINP.n300 VINP.n179 4.5005
R47263 VINP.n265 VINP.n179 4.5005
R47264 VINP.n302 VINP.n179 4.5005
R47265 VINP.n264 VINP.n179 4.5005
R47266 VINP.n304 VINP.n179 4.5005
R47267 VINP.n263 VINP.n179 4.5005
R47268 VINP.n306 VINP.n179 4.5005
R47269 VINP.n262 VINP.n179 4.5005
R47270 VINP.n308 VINP.n179 4.5005
R47271 VINP.n261 VINP.n179 4.5005
R47272 VINP.n310 VINP.n179 4.5005
R47273 VINP.n260 VINP.n179 4.5005
R47274 VINP.n312 VINP.n179 4.5005
R47275 VINP.n259 VINP.n179 4.5005
R47276 VINP.n314 VINP.n179 4.5005
R47277 VINP.n258 VINP.n179 4.5005
R47278 VINP.n316 VINP.n179 4.5005
R47279 VINP.n257 VINP.n179 4.5005
R47280 VINP.n318 VINP.n179 4.5005
R47281 VINP.n256 VINP.n179 4.5005
R47282 VINP.n320 VINP.n179 4.5005
R47283 VINP.n255 VINP.n179 4.5005
R47284 VINP.n322 VINP.n179 4.5005
R47285 VINP.n254 VINP.n179 4.5005
R47286 VINP.n324 VINP.n179 4.5005
R47287 VINP.n253 VINP.n179 4.5005
R47288 VINP.n326 VINP.n179 4.5005
R47289 VINP.n252 VINP.n179 4.5005
R47290 VINP.n328 VINP.n179 4.5005
R47291 VINP.n251 VINP.n179 4.5005
R47292 VINP.n330 VINP.n179 4.5005
R47293 VINP.n250 VINP.n179 4.5005
R47294 VINP.n332 VINP.n179 4.5005
R47295 VINP.n249 VINP.n179 4.5005
R47296 VINP.n334 VINP.n179 4.5005
R47297 VINP.n248 VINP.n179 4.5005
R47298 VINP.n336 VINP.n179 4.5005
R47299 VINP.n247 VINP.n179 4.5005
R47300 VINP.n338 VINP.n179 4.5005
R47301 VINP.n246 VINP.n179 4.5005
R47302 VINP.n340 VINP.n179 4.5005
R47303 VINP.n245 VINP.n179 4.5005
R47304 VINP.n342 VINP.n179 4.5005
R47305 VINP.n244 VINP.n179 4.5005
R47306 VINP.n344 VINP.n179 4.5005
R47307 VINP.n243 VINP.n179 4.5005
R47308 VINP.n346 VINP.n179 4.5005
R47309 VINP.n242 VINP.n179 4.5005
R47310 VINP.n348 VINP.n179 4.5005
R47311 VINP.n241 VINP.n179 4.5005
R47312 VINP.n350 VINP.n179 4.5005
R47313 VINP.n240 VINP.n179 4.5005
R47314 VINP.n352 VINP.n179 4.5005
R47315 VINP.n239 VINP.n179 4.5005
R47316 VINP.n354 VINP.n179 4.5005
R47317 VINP.n238 VINP.n179 4.5005
R47318 VINP.n356 VINP.n179 4.5005
R47319 VINP.n237 VINP.n179 4.5005
R47320 VINP.n358 VINP.n179 4.5005
R47321 VINP.n236 VINP.n179 4.5005
R47322 VINP.n360 VINP.n179 4.5005
R47323 VINP.n235 VINP.n179 4.5005
R47324 VINP.n362 VINP.n179 4.5005
R47325 VINP.n234 VINP.n179 4.5005
R47326 VINP.n364 VINP.n179 4.5005
R47327 VINP.n233 VINP.n179 4.5005
R47328 VINP.n366 VINP.n179 4.5005
R47329 VINP.n232 VINP.n179 4.5005
R47330 VINP.n368 VINP.n179 4.5005
R47331 VINP.n231 VINP.n179 4.5005
R47332 VINP.n370 VINP.n179 4.5005
R47333 VINP.n230 VINP.n179 4.5005
R47334 VINP.n372 VINP.n179 4.5005
R47335 VINP.n229 VINP.n179 4.5005
R47336 VINP.n374 VINP.n179 4.5005
R47337 VINP.n228 VINP.n179 4.5005
R47338 VINP.n376 VINP.n179 4.5005
R47339 VINP.n227 VINP.n179 4.5005
R47340 VINP.n378 VINP.n179 4.5005
R47341 VINP.n226 VINP.n179 4.5005
R47342 VINP.n380 VINP.n179 4.5005
R47343 VINP.n225 VINP.n179 4.5005
R47344 VINP.n382 VINP.n179 4.5005
R47345 VINP.n224 VINP.n179 4.5005
R47346 VINP.n384 VINP.n179 4.5005
R47347 VINP.n223 VINP.n179 4.5005
R47348 VINP.n386 VINP.n179 4.5005
R47349 VINP.n222 VINP.n179 4.5005
R47350 VINP.n388 VINP.n179 4.5005
R47351 VINP.n221 VINP.n179 4.5005
R47352 VINP.n390 VINP.n179 4.5005
R47353 VINP.n220 VINP.n179 4.5005
R47354 VINP.n392 VINP.n179 4.5005
R47355 VINP.n219 VINP.n179 4.5005
R47356 VINP.n394 VINP.n179 4.5005
R47357 VINP.n218 VINP.n179 4.5005
R47358 VINP.n396 VINP.n179 4.5005
R47359 VINP.n217 VINP.n179 4.5005
R47360 VINP.n398 VINP.n179 4.5005
R47361 VINP.n216 VINP.n179 4.5005
R47362 VINP.n400 VINP.n179 4.5005
R47363 VINP.n215 VINP.n179 4.5005
R47364 VINP.n654 VINP.n179 4.5005
R47365 VINP.n656 VINP.n179 4.5005
R47366 VINP.n179 VINP.n0 4.5005
R47367 VINP.n278 VINP.n121 4.5005
R47368 VINP.n276 VINP.n121 4.5005
R47369 VINP.n280 VINP.n121 4.5005
R47370 VINP.n275 VINP.n121 4.5005
R47371 VINP.n282 VINP.n121 4.5005
R47372 VINP.n274 VINP.n121 4.5005
R47373 VINP.n284 VINP.n121 4.5005
R47374 VINP.n273 VINP.n121 4.5005
R47375 VINP.n286 VINP.n121 4.5005
R47376 VINP.n272 VINP.n121 4.5005
R47377 VINP.n288 VINP.n121 4.5005
R47378 VINP.n271 VINP.n121 4.5005
R47379 VINP.n290 VINP.n121 4.5005
R47380 VINP.n270 VINP.n121 4.5005
R47381 VINP.n292 VINP.n121 4.5005
R47382 VINP.n269 VINP.n121 4.5005
R47383 VINP.n294 VINP.n121 4.5005
R47384 VINP.n268 VINP.n121 4.5005
R47385 VINP.n296 VINP.n121 4.5005
R47386 VINP.n267 VINP.n121 4.5005
R47387 VINP.n298 VINP.n121 4.5005
R47388 VINP.n266 VINP.n121 4.5005
R47389 VINP.n300 VINP.n121 4.5005
R47390 VINP.n265 VINP.n121 4.5005
R47391 VINP.n302 VINP.n121 4.5005
R47392 VINP.n264 VINP.n121 4.5005
R47393 VINP.n304 VINP.n121 4.5005
R47394 VINP.n263 VINP.n121 4.5005
R47395 VINP.n306 VINP.n121 4.5005
R47396 VINP.n262 VINP.n121 4.5005
R47397 VINP.n308 VINP.n121 4.5005
R47398 VINP.n261 VINP.n121 4.5005
R47399 VINP.n310 VINP.n121 4.5005
R47400 VINP.n260 VINP.n121 4.5005
R47401 VINP.n312 VINP.n121 4.5005
R47402 VINP.n259 VINP.n121 4.5005
R47403 VINP.n314 VINP.n121 4.5005
R47404 VINP.n258 VINP.n121 4.5005
R47405 VINP.n316 VINP.n121 4.5005
R47406 VINP.n257 VINP.n121 4.5005
R47407 VINP.n318 VINP.n121 4.5005
R47408 VINP.n256 VINP.n121 4.5005
R47409 VINP.n320 VINP.n121 4.5005
R47410 VINP.n255 VINP.n121 4.5005
R47411 VINP.n322 VINP.n121 4.5005
R47412 VINP.n254 VINP.n121 4.5005
R47413 VINP.n324 VINP.n121 4.5005
R47414 VINP.n253 VINP.n121 4.5005
R47415 VINP.n326 VINP.n121 4.5005
R47416 VINP.n252 VINP.n121 4.5005
R47417 VINP.n328 VINP.n121 4.5005
R47418 VINP.n251 VINP.n121 4.5005
R47419 VINP.n330 VINP.n121 4.5005
R47420 VINP.n250 VINP.n121 4.5005
R47421 VINP.n332 VINP.n121 4.5005
R47422 VINP.n249 VINP.n121 4.5005
R47423 VINP.n334 VINP.n121 4.5005
R47424 VINP.n248 VINP.n121 4.5005
R47425 VINP.n336 VINP.n121 4.5005
R47426 VINP.n247 VINP.n121 4.5005
R47427 VINP.n338 VINP.n121 4.5005
R47428 VINP.n246 VINP.n121 4.5005
R47429 VINP.n340 VINP.n121 4.5005
R47430 VINP.n245 VINP.n121 4.5005
R47431 VINP.n342 VINP.n121 4.5005
R47432 VINP.n244 VINP.n121 4.5005
R47433 VINP.n344 VINP.n121 4.5005
R47434 VINP.n243 VINP.n121 4.5005
R47435 VINP.n346 VINP.n121 4.5005
R47436 VINP.n242 VINP.n121 4.5005
R47437 VINP.n348 VINP.n121 4.5005
R47438 VINP.n241 VINP.n121 4.5005
R47439 VINP.n350 VINP.n121 4.5005
R47440 VINP.n240 VINP.n121 4.5005
R47441 VINP.n352 VINP.n121 4.5005
R47442 VINP.n239 VINP.n121 4.5005
R47443 VINP.n354 VINP.n121 4.5005
R47444 VINP.n238 VINP.n121 4.5005
R47445 VINP.n356 VINP.n121 4.5005
R47446 VINP.n237 VINP.n121 4.5005
R47447 VINP.n358 VINP.n121 4.5005
R47448 VINP.n236 VINP.n121 4.5005
R47449 VINP.n360 VINP.n121 4.5005
R47450 VINP.n235 VINP.n121 4.5005
R47451 VINP.n362 VINP.n121 4.5005
R47452 VINP.n234 VINP.n121 4.5005
R47453 VINP.n364 VINP.n121 4.5005
R47454 VINP.n233 VINP.n121 4.5005
R47455 VINP.n366 VINP.n121 4.5005
R47456 VINP.n232 VINP.n121 4.5005
R47457 VINP.n368 VINP.n121 4.5005
R47458 VINP.n231 VINP.n121 4.5005
R47459 VINP.n370 VINP.n121 4.5005
R47460 VINP.n230 VINP.n121 4.5005
R47461 VINP.n372 VINP.n121 4.5005
R47462 VINP.n229 VINP.n121 4.5005
R47463 VINP.n374 VINP.n121 4.5005
R47464 VINP.n228 VINP.n121 4.5005
R47465 VINP.n376 VINP.n121 4.5005
R47466 VINP.n227 VINP.n121 4.5005
R47467 VINP.n378 VINP.n121 4.5005
R47468 VINP.n226 VINP.n121 4.5005
R47469 VINP.n380 VINP.n121 4.5005
R47470 VINP.n225 VINP.n121 4.5005
R47471 VINP.n382 VINP.n121 4.5005
R47472 VINP.n224 VINP.n121 4.5005
R47473 VINP.n384 VINP.n121 4.5005
R47474 VINP.n223 VINP.n121 4.5005
R47475 VINP.n386 VINP.n121 4.5005
R47476 VINP.n222 VINP.n121 4.5005
R47477 VINP.n388 VINP.n121 4.5005
R47478 VINP.n221 VINP.n121 4.5005
R47479 VINP.n390 VINP.n121 4.5005
R47480 VINP.n220 VINP.n121 4.5005
R47481 VINP.n392 VINP.n121 4.5005
R47482 VINP.n219 VINP.n121 4.5005
R47483 VINP.n394 VINP.n121 4.5005
R47484 VINP.n218 VINP.n121 4.5005
R47485 VINP.n396 VINP.n121 4.5005
R47486 VINP.n217 VINP.n121 4.5005
R47487 VINP.n398 VINP.n121 4.5005
R47488 VINP.n216 VINP.n121 4.5005
R47489 VINP.n400 VINP.n121 4.5005
R47490 VINP.n215 VINP.n121 4.5005
R47491 VINP.n654 VINP.n121 4.5005
R47492 VINP.n656 VINP.n121 4.5005
R47493 VINP.n121 VINP.n0 4.5005
R47494 VINP.n278 VINP.n180 4.5005
R47495 VINP.n276 VINP.n180 4.5005
R47496 VINP.n280 VINP.n180 4.5005
R47497 VINP.n275 VINP.n180 4.5005
R47498 VINP.n282 VINP.n180 4.5005
R47499 VINP.n274 VINP.n180 4.5005
R47500 VINP.n284 VINP.n180 4.5005
R47501 VINP.n273 VINP.n180 4.5005
R47502 VINP.n286 VINP.n180 4.5005
R47503 VINP.n272 VINP.n180 4.5005
R47504 VINP.n288 VINP.n180 4.5005
R47505 VINP.n271 VINP.n180 4.5005
R47506 VINP.n290 VINP.n180 4.5005
R47507 VINP.n270 VINP.n180 4.5005
R47508 VINP.n292 VINP.n180 4.5005
R47509 VINP.n269 VINP.n180 4.5005
R47510 VINP.n294 VINP.n180 4.5005
R47511 VINP.n268 VINP.n180 4.5005
R47512 VINP.n296 VINP.n180 4.5005
R47513 VINP.n267 VINP.n180 4.5005
R47514 VINP.n298 VINP.n180 4.5005
R47515 VINP.n266 VINP.n180 4.5005
R47516 VINP.n300 VINP.n180 4.5005
R47517 VINP.n265 VINP.n180 4.5005
R47518 VINP.n302 VINP.n180 4.5005
R47519 VINP.n264 VINP.n180 4.5005
R47520 VINP.n304 VINP.n180 4.5005
R47521 VINP.n263 VINP.n180 4.5005
R47522 VINP.n306 VINP.n180 4.5005
R47523 VINP.n262 VINP.n180 4.5005
R47524 VINP.n308 VINP.n180 4.5005
R47525 VINP.n261 VINP.n180 4.5005
R47526 VINP.n310 VINP.n180 4.5005
R47527 VINP.n260 VINP.n180 4.5005
R47528 VINP.n312 VINP.n180 4.5005
R47529 VINP.n259 VINP.n180 4.5005
R47530 VINP.n314 VINP.n180 4.5005
R47531 VINP.n258 VINP.n180 4.5005
R47532 VINP.n316 VINP.n180 4.5005
R47533 VINP.n257 VINP.n180 4.5005
R47534 VINP.n318 VINP.n180 4.5005
R47535 VINP.n256 VINP.n180 4.5005
R47536 VINP.n320 VINP.n180 4.5005
R47537 VINP.n255 VINP.n180 4.5005
R47538 VINP.n322 VINP.n180 4.5005
R47539 VINP.n254 VINP.n180 4.5005
R47540 VINP.n324 VINP.n180 4.5005
R47541 VINP.n253 VINP.n180 4.5005
R47542 VINP.n326 VINP.n180 4.5005
R47543 VINP.n252 VINP.n180 4.5005
R47544 VINP.n328 VINP.n180 4.5005
R47545 VINP.n251 VINP.n180 4.5005
R47546 VINP.n330 VINP.n180 4.5005
R47547 VINP.n250 VINP.n180 4.5005
R47548 VINP.n332 VINP.n180 4.5005
R47549 VINP.n249 VINP.n180 4.5005
R47550 VINP.n334 VINP.n180 4.5005
R47551 VINP.n248 VINP.n180 4.5005
R47552 VINP.n336 VINP.n180 4.5005
R47553 VINP.n247 VINP.n180 4.5005
R47554 VINP.n338 VINP.n180 4.5005
R47555 VINP.n246 VINP.n180 4.5005
R47556 VINP.n340 VINP.n180 4.5005
R47557 VINP.n245 VINP.n180 4.5005
R47558 VINP.n342 VINP.n180 4.5005
R47559 VINP.n244 VINP.n180 4.5005
R47560 VINP.n344 VINP.n180 4.5005
R47561 VINP.n243 VINP.n180 4.5005
R47562 VINP.n346 VINP.n180 4.5005
R47563 VINP.n242 VINP.n180 4.5005
R47564 VINP.n348 VINP.n180 4.5005
R47565 VINP.n241 VINP.n180 4.5005
R47566 VINP.n350 VINP.n180 4.5005
R47567 VINP.n240 VINP.n180 4.5005
R47568 VINP.n352 VINP.n180 4.5005
R47569 VINP.n239 VINP.n180 4.5005
R47570 VINP.n354 VINP.n180 4.5005
R47571 VINP.n238 VINP.n180 4.5005
R47572 VINP.n356 VINP.n180 4.5005
R47573 VINP.n237 VINP.n180 4.5005
R47574 VINP.n358 VINP.n180 4.5005
R47575 VINP.n236 VINP.n180 4.5005
R47576 VINP.n360 VINP.n180 4.5005
R47577 VINP.n235 VINP.n180 4.5005
R47578 VINP.n362 VINP.n180 4.5005
R47579 VINP.n234 VINP.n180 4.5005
R47580 VINP.n364 VINP.n180 4.5005
R47581 VINP.n233 VINP.n180 4.5005
R47582 VINP.n366 VINP.n180 4.5005
R47583 VINP.n232 VINP.n180 4.5005
R47584 VINP.n368 VINP.n180 4.5005
R47585 VINP.n231 VINP.n180 4.5005
R47586 VINP.n370 VINP.n180 4.5005
R47587 VINP.n230 VINP.n180 4.5005
R47588 VINP.n372 VINP.n180 4.5005
R47589 VINP.n229 VINP.n180 4.5005
R47590 VINP.n374 VINP.n180 4.5005
R47591 VINP.n228 VINP.n180 4.5005
R47592 VINP.n376 VINP.n180 4.5005
R47593 VINP.n227 VINP.n180 4.5005
R47594 VINP.n378 VINP.n180 4.5005
R47595 VINP.n226 VINP.n180 4.5005
R47596 VINP.n380 VINP.n180 4.5005
R47597 VINP.n225 VINP.n180 4.5005
R47598 VINP.n382 VINP.n180 4.5005
R47599 VINP.n224 VINP.n180 4.5005
R47600 VINP.n384 VINP.n180 4.5005
R47601 VINP.n223 VINP.n180 4.5005
R47602 VINP.n386 VINP.n180 4.5005
R47603 VINP.n222 VINP.n180 4.5005
R47604 VINP.n388 VINP.n180 4.5005
R47605 VINP.n221 VINP.n180 4.5005
R47606 VINP.n390 VINP.n180 4.5005
R47607 VINP.n220 VINP.n180 4.5005
R47608 VINP.n392 VINP.n180 4.5005
R47609 VINP.n219 VINP.n180 4.5005
R47610 VINP.n394 VINP.n180 4.5005
R47611 VINP.n218 VINP.n180 4.5005
R47612 VINP.n396 VINP.n180 4.5005
R47613 VINP.n217 VINP.n180 4.5005
R47614 VINP.n398 VINP.n180 4.5005
R47615 VINP.n216 VINP.n180 4.5005
R47616 VINP.n400 VINP.n180 4.5005
R47617 VINP.n215 VINP.n180 4.5005
R47618 VINP.n654 VINP.n180 4.5005
R47619 VINP.n656 VINP.n180 4.5005
R47620 VINP.n180 VINP.n0 4.5005
R47621 VINP.n278 VINP.n120 4.5005
R47622 VINP.n276 VINP.n120 4.5005
R47623 VINP.n280 VINP.n120 4.5005
R47624 VINP.n275 VINP.n120 4.5005
R47625 VINP.n282 VINP.n120 4.5005
R47626 VINP.n274 VINP.n120 4.5005
R47627 VINP.n284 VINP.n120 4.5005
R47628 VINP.n273 VINP.n120 4.5005
R47629 VINP.n286 VINP.n120 4.5005
R47630 VINP.n272 VINP.n120 4.5005
R47631 VINP.n288 VINP.n120 4.5005
R47632 VINP.n271 VINP.n120 4.5005
R47633 VINP.n290 VINP.n120 4.5005
R47634 VINP.n270 VINP.n120 4.5005
R47635 VINP.n292 VINP.n120 4.5005
R47636 VINP.n269 VINP.n120 4.5005
R47637 VINP.n294 VINP.n120 4.5005
R47638 VINP.n268 VINP.n120 4.5005
R47639 VINP.n296 VINP.n120 4.5005
R47640 VINP.n267 VINP.n120 4.5005
R47641 VINP.n298 VINP.n120 4.5005
R47642 VINP.n266 VINP.n120 4.5005
R47643 VINP.n300 VINP.n120 4.5005
R47644 VINP.n265 VINP.n120 4.5005
R47645 VINP.n302 VINP.n120 4.5005
R47646 VINP.n264 VINP.n120 4.5005
R47647 VINP.n304 VINP.n120 4.5005
R47648 VINP.n263 VINP.n120 4.5005
R47649 VINP.n306 VINP.n120 4.5005
R47650 VINP.n262 VINP.n120 4.5005
R47651 VINP.n308 VINP.n120 4.5005
R47652 VINP.n261 VINP.n120 4.5005
R47653 VINP.n310 VINP.n120 4.5005
R47654 VINP.n260 VINP.n120 4.5005
R47655 VINP.n312 VINP.n120 4.5005
R47656 VINP.n259 VINP.n120 4.5005
R47657 VINP.n314 VINP.n120 4.5005
R47658 VINP.n258 VINP.n120 4.5005
R47659 VINP.n316 VINP.n120 4.5005
R47660 VINP.n257 VINP.n120 4.5005
R47661 VINP.n318 VINP.n120 4.5005
R47662 VINP.n256 VINP.n120 4.5005
R47663 VINP.n320 VINP.n120 4.5005
R47664 VINP.n255 VINP.n120 4.5005
R47665 VINP.n322 VINP.n120 4.5005
R47666 VINP.n254 VINP.n120 4.5005
R47667 VINP.n324 VINP.n120 4.5005
R47668 VINP.n253 VINP.n120 4.5005
R47669 VINP.n326 VINP.n120 4.5005
R47670 VINP.n252 VINP.n120 4.5005
R47671 VINP.n328 VINP.n120 4.5005
R47672 VINP.n251 VINP.n120 4.5005
R47673 VINP.n330 VINP.n120 4.5005
R47674 VINP.n250 VINP.n120 4.5005
R47675 VINP.n332 VINP.n120 4.5005
R47676 VINP.n249 VINP.n120 4.5005
R47677 VINP.n334 VINP.n120 4.5005
R47678 VINP.n248 VINP.n120 4.5005
R47679 VINP.n336 VINP.n120 4.5005
R47680 VINP.n247 VINP.n120 4.5005
R47681 VINP.n338 VINP.n120 4.5005
R47682 VINP.n246 VINP.n120 4.5005
R47683 VINP.n340 VINP.n120 4.5005
R47684 VINP.n245 VINP.n120 4.5005
R47685 VINP.n342 VINP.n120 4.5005
R47686 VINP.n244 VINP.n120 4.5005
R47687 VINP.n344 VINP.n120 4.5005
R47688 VINP.n243 VINP.n120 4.5005
R47689 VINP.n346 VINP.n120 4.5005
R47690 VINP.n242 VINP.n120 4.5005
R47691 VINP.n348 VINP.n120 4.5005
R47692 VINP.n241 VINP.n120 4.5005
R47693 VINP.n350 VINP.n120 4.5005
R47694 VINP.n240 VINP.n120 4.5005
R47695 VINP.n352 VINP.n120 4.5005
R47696 VINP.n239 VINP.n120 4.5005
R47697 VINP.n354 VINP.n120 4.5005
R47698 VINP.n238 VINP.n120 4.5005
R47699 VINP.n356 VINP.n120 4.5005
R47700 VINP.n237 VINP.n120 4.5005
R47701 VINP.n358 VINP.n120 4.5005
R47702 VINP.n236 VINP.n120 4.5005
R47703 VINP.n360 VINP.n120 4.5005
R47704 VINP.n235 VINP.n120 4.5005
R47705 VINP.n362 VINP.n120 4.5005
R47706 VINP.n234 VINP.n120 4.5005
R47707 VINP.n364 VINP.n120 4.5005
R47708 VINP.n233 VINP.n120 4.5005
R47709 VINP.n366 VINP.n120 4.5005
R47710 VINP.n232 VINP.n120 4.5005
R47711 VINP.n368 VINP.n120 4.5005
R47712 VINP.n231 VINP.n120 4.5005
R47713 VINP.n370 VINP.n120 4.5005
R47714 VINP.n230 VINP.n120 4.5005
R47715 VINP.n372 VINP.n120 4.5005
R47716 VINP.n229 VINP.n120 4.5005
R47717 VINP.n374 VINP.n120 4.5005
R47718 VINP.n228 VINP.n120 4.5005
R47719 VINP.n376 VINP.n120 4.5005
R47720 VINP.n227 VINP.n120 4.5005
R47721 VINP.n378 VINP.n120 4.5005
R47722 VINP.n226 VINP.n120 4.5005
R47723 VINP.n380 VINP.n120 4.5005
R47724 VINP.n225 VINP.n120 4.5005
R47725 VINP.n382 VINP.n120 4.5005
R47726 VINP.n224 VINP.n120 4.5005
R47727 VINP.n384 VINP.n120 4.5005
R47728 VINP.n223 VINP.n120 4.5005
R47729 VINP.n386 VINP.n120 4.5005
R47730 VINP.n222 VINP.n120 4.5005
R47731 VINP.n388 VINP.n120 4.5005
R47732 VINP.n221 VINP.n120 4.5005
R47733 VINP.n390 VINP.n120 4.5005
R47734 VINP.n220 VINP.n120 4.5005
R47735 VINP.n392 VINP.n120 4.5005
R47736 VINP.n219 VINP.n120 4.5005
R47737 VINP.n394 VINP.n120 4.5005
R47738 VINP.n218 VINP.n120 4.5005
R47739 VINP.n396 VINP.n120 4.5005
R47740 VINP.n217 VINP.n120 4.5005
R47741 VINP.n398 VINP.n120 4.5005
R47742 VINP.n216 VINP.n120 4.5005
R47743 VINP.n400 VINP.n120 4.5005
R47744 VINP.n215 VINP.n120 4.5005
R47745 VINP.n654 VINP.n120 4.5005
R47746 VINP.n656 VINP.n120 4.5005
R47747 VINP.n120 VINP.n0 4.5005
R47748 VINP.n278 VINP.n181 4.5005
R47749 VINP.n276 VINP.n181 4.5005
R47750 VINP.n280 VINP.n181 4.5005
R47751 VINP.n275 VINP.n181 4.5005
R47752 VINP.n282 VINP.n181 4.5005
R47753 VINP.n274 VINP.n181 4.5005
R47754 VINP.n284 VINP.n181 4.5005
R47755 VINP.n273 VINP.n181 4.5005
R47756 VINP.n286 VINP.n181 4.5005
R47757 VINP.n272 VINP.n181 4.5005
R47758 VINP.n288 VINP.n181 4.5005
R47759 VINP.n271 VINP.n181 4.5005
R47760 VINP.n290 VINP.n181 4.5005
R47761 VINP.n270 VINP.n181 4.5005
R47762 VINP.n292 VINP.n181 4.5005
R47763 VINP.n269 VINP.n181 4.5005
R47764 VINP.n294 VINP.n181 4.5005
R47765 VINP.n268 VINP.n181 4.5005
R47766 VINP.n296 VINP.n181 4.5005
R47767 VINP.n267 VINP.n181 4.5005
R47768 VINP.n298 VINP.n181 4.5005
R47769 VINP.n266 VINP.n181 4.5005
R47770 VINP.n300 VINP.n181 4.5005
R47771 VINP.n265 VINP.n181 4.5005
R47772 VINP.n302 VINP.n181 4.5005
R47773 VINP.n264 VINP.n181 4.5005
R47774 VINP.n304 VINP.n181 4.5005
R47775 VINP.n263 VINP.n181 4.5005
R47776 VINP.n306 VINP.n181 4.5005
R47777 VINP.n262 VINP.n181 4.5005
R47778 VINP.n308 VINP.n181 4.5005
R47779 VINP.n261 VINP.n181 4.5005
R47780 VINP.n310 VINP.n181 4.5005
R47781 VINP.n260 VINP.n181 4.5005
R47782 VINP.n312 VINP.n181 4.5005
R47783 VINP.n259 VINP.n181 4.5005
R47784 VINP.n314 VINP.n181 4.5005
R47785 VINP.n258 VINP.n181 4.5005
R47786 VINP.n316 VINP.n181 4.5005
R47787 VINP.n257 VINP.n181 4.5005
R47788 VINP.n318 VINP.n181 4.5005
R47789 VINP.n256 VINP.n181 4.5005
R47790 VINP.n320 VINP.n181 4.5005
R47791 VINP.n255 VINP.n181 4.5005
R47792 VINP.n322 VINP.n181 4.5005
R47793 VINP.n254 VINP.n181 4.5005
R47794 VINP.n324 VINP.n181 4.5005
R47795 VINP.n253 VINP.n181 4.5005
R47796 VINP.n326 VINP.n181 4.5005
R47797 VINP.n252 VINP.n181 4.5005
R47798 VINP.n328 VINP.n181 4.5005
R47799 VINP.n251 VINP.n181 4.5005
R47800 VINP.n330 VINP.n181 4.5005
R47801 VINP.n250 VINP.n181 4.5005
R47802 VINP.n332 VINP.n181 4.5005
R47803 VINP.n249 VINP.n181 4.5005
R47804 VINP.n334 VINP.n181 4.5005
R47805 VINP.n248 VINP.n181 4.5005
R47806 VINP.n336 VINP.n181 4.5005
R47807 VINP.n247 VINP.n181 4.5005
R47808 VINP.n338 VINP.n181 4.5005
R47809 VINP.n246 VINP.n181 4.5005
R47810 VINP.n340 VINP.n181 4.5005
R47811 VINP.n245 VINP.n181 4.5005
R47812 VINP.n342 VINP.n181 4.5005
R47813 VINP.n244 VINP.n181 4.5005
R47814 VINP.n344 VINP.n181 4.5005
R47815 VINP.n243 VINP.n181 4.5005
R47816 VINP.n346 VINP.n181 4.5005
R47817 VINP.n242 VINP.n181 4.5005
R47818 VINP.n348 VINP.n181 4.5005
R47819 VINP.n241 VINP.n181 4.5005
R47820 VINP.n350 VINP.n181 4.5005
R47821 VINP.n240 VINP.n181 4.5005
R47822 VINP.n352 VINP.n181 4.5005
R47823 VINP.n239 VINP.n181 4.5005
R47824 VINP.n354 VINP.n181 4.5005
R47825 VINP.n238 VINP.n181 4.5005
R47826 VINP.n356 VINP.n181 4.5005
R47827 VINP.n237 VINP.n181 4.5005
R47828 VINP.n358 VINP.n181 4.5005
R47829 VINP.n236 VINP.n181 4.5005
R47830 VINP.n360 VINP.n181 4.5005
R47831 VINP.n235 VINP.n181 4.5005
R47832 VINP.n362 VINP.n181 4.5005
R47833 VINP.n234 VINP.n181 4.5005
R47834 VINP.n364 VINP.n181 4.5005
R47835 VINP.n233 VINP.n181 4.5005
R47836 VINP.n366 VINP.n181 4.5005
R47837 VINP.n232 VINP.n181 4.5005
R47838 VINP.n368 VINP.n181 4.5005
R47839 VINP.n231 VINP.n181 4.5005
R47840 VINP.n370 VINP.n181 4.5005
R47841 VINP.n230 VINP.n181 4.5005
R47842 VINP.n372 VINP.n181 4.5005
R47843 VINP.n229 VINP.n181 4.5005
R47844 VINP.n374 VINP.n181 4.5005
R47845 VINP.n228 VINP.n181 4.5005
R47846 VINP.n376 VINP.n181 4.5005
R47847 VINP.n227 VINP.n181 4.5005
R47848 VINP.n378 VINP.n181 4.5005
R47849 VINP.n226 VINP.n181 4.5005
R47850 VINP.n380 VINP.n181 4.5005
R47851 VINP.n225 VINP.n181 4.5005
R47852 VINP.n382 VINP.n181 4.5005
R47853 VINP.n224 VINP.n181 4.5005
R47854 VINP.n384 VINP.n181 4.5005
R47855 VINP.n223 VINP.n181 4.5005
R47856 VINP.n386 VINP.n181 4.5005
R47857 VINP.n222 VINP.n181 4.5005
R47858 VINP.n388 VINP.n181 4.5005
R47859 VINP.n221 VINP.n181 4.5005
R47860 VINP.n390 VINP.n181 4.5005
R47861 VINP.n220 VINP.n181 4.5005
R47862 VINP.n392 VINP.n181 4.5005
R47863 VINP.n219 VINP.n181 4.5005
R47864 VINP.n394 VINP.n181 4.5005
R47865 VINP.n218 VINP.n181 4.5005
R47866 VINP.n396 VINP.n181 4.5005
R47867 VINP.n217 VINP.n181 4.5005
R47868 VINP.n398 VINP.n181 4.5005
R47869 VINP.n216 VINP.n181 4.5005
R47870 VINP.n400 VINP.n181 4.5005
R47871 VINP.n215 VINP.n181 4.5005
R47872 VINP.n654 VINP.n181 4.5005
R47873 VINP.n656 VINP.n181 4.5005
R47874 VINP.n181 VINP.n0 4.5005
R47875 VINP.n278 VINP.n119 4.5005
R47876 VINP.n276 VINP.n119 4.5005
R47877 VINP.n280 VINP.n119 4.5005
R47878 VINP.n275 VINP.n119 4.5005
R47879 VINP.n282 VINP.n119 4.5005
R47880 VINP.n274 VINP.n119 4.5005
R47881 VINP.n284 VINP.n119 4.5005
R47882 VINP.n273 VINP.n119 4.5005
R47883 VINP.n286 VINP.n119 4.5005
R47884 VINP.n272 VINP.n119 4.5005
R47885 VINP.n288 VINP.n119 4.5005
R47886 VINP.n271 VINP.n119 4.5005
R47887 VINP.n290 VINP.n119 4.5005
R47888 VINP.n270 VINP.n119 4.5005
R47889 VINP.n292 VINP.n119 4.5005
R47890 VINP.n269 VINP.n119 4.5005
R47891 VINP.n294 VINP.n119 4.5005
R47892 VINP.n268 VINP.n119 4.5005
R47893 VINP.n296 VINP.n119 4.5005
R47894 VINP.n267 VINP.n119 4.5005
R47895 VINP.n298 VINP.n119 4.5005
R47896 VINP.n266 VINP.n119 4.5005
R47897 VINP.n300 VINP.n119 4.5005
R47898 VINP.n265 VINP.n119 4.5005
R47899 VINP.n302 VINP.n119 4.5005
R47900 VINP.n264 VINP.n119 4.5005
R47901 VINP.n304 VINP.n119 4.5005
R47902 VINP.n263 VINP.n119 4.5005
R47903 VINP.n306 VINP.n119 4.5005
R47904 VINP.n262 VINP.n119 4.5005
R47905 VINP.n308 VINP.n119 4.5005
R47906 VINP.n261 VINP.n119 4.5005
R47907 VINP.n310 VINP.n119 4.5005
R47908 VINP.n260 VINP.n119 4.5005
R47909 VINP.n312 VINP.n119 4.5005
R47910 VINP.n259 VINP.n119 4.5005
R47911 VINP.n314 VINP.n119 4.5005
R47912 VINP.n258 VINP.n119 4.5005
R47913 VINP.n316 VINP.n119 4.5005
R47914 VINP.n257 VINP.n119 4.5005
R47915 VINP.n318 VINP.n119 4.5005
R47916 VINP.n256 VINP.n119 4.5005
R47917 VINP.n320 VINP.n119 4.5005
R47918 VINP.n255 VINP.n119 4.5005
R47919 VINP.n322 VINP.n119 4.5005
R47920 VINP.n254 VINP.n119 4.5005
R47921 VINP.n324 VINP.n119 4.5005
R47922 VINP.n253 VINP.n119 4.5005
R47923 VINP.n326 VINP.n119 4.5005
R47924 VINP.n252 VINP.n119 4.5005
R47925 VINP.n328 VINP.n119 4.5005
R47926 VINP.n251 VINP.n119 4.5005
R47927 VINP.n330 VINP.n119 4.5005
R47928 VINP.n250 VINP.n119 4.5005
R47929 VINP.n332 VINP.n119 4.5005
R47930 VINP.n249 VINP.n119 4.5005
R47931 VINP.n334 VINP.n119 4.5005
R47932 VINP.n248 VINP.n119 4.5005
R47933 VINP.n336 VINP.n119 4.5005
R47934 VINP.n247 VINP.n119 4.5005
R47935 VINP.n338 VINP.n119 4.5005
R47936 VINP.n246 VINP.n119 4.5005
R47937 VINP.n340 VINP.n119 4.5005
R47938 VINP.n245 VINP.n119 4.5005
R47939 VINP.n342 VINP.n119 4.5005
R47940 VINP.n244 VINP.n119 4.5005
R47941 VINP.n344 VINP.n119 4.5005
R47942 VINP.n243 VINP.n119 4.5005
R47943 VINP.n346 VINP.n119 4.5005
R47944 VINP.n242 VINP.n119 4.5005
R47945 VINP.n348 VINP.n119 4.5005
R47946 VINP.n241 VINP.n119 4.5005
R47947 VINP.n350 VINP.n119 4.5005
R47948 VINP.n240 VINP.n119 4.5005
R47949 VINP.n352 VINP.n119 4.5005
R47950 VINP.n239 VINP.n119 4.5005
R47951 VINP.n354 VINP.n119 4.5005
R47952 VINP.n238 VINP.n119 4.5005
R47953 VINP.n356 VINP.n119 4.5005
R47954 VINP.n237 VINP.n119 4.5005
R47955 VINP.n358 VINP.n119 4.5005
R47956 VINP.n236 VINP.n119 4.5005
R47957 VINP.n360 VINP.n119 4.5005
R47958 VINP.n235 VINP.n119 4.5005
R47959 VINP.n362 VINP.n119 4.5005
R47960 VINP.n234 VINP.n119 4.5005
R47961 VINP.n364 VINP.n119 4.5005
R47962 VINP.n233 VINP.n119 4.5005
R47963 VINP.n366 VINP.n119 4.5005
R47964 VINP.n232 VINP.n119 4.5005
R47965 VINP.n368 VINP.n119 4.5005
R47966 VINP.n231 VINP.n119 4.5005
R47967 VINP.n370 VINP.n119 4.5005
R47968 VINP.n230 VINP.n119 4.5005
R47969 VINP.n372 VINP.n119 4.5005
R47970 VINP.n229 VINP.n119 4.5005
R47971 VINP.n374 VINP.n119 4.5005
R47972 VINP.n228 VINP.n119 4.5005
R47973 VINP.n376 VINP.n119 4.5005
R47974 VINP.n227 VINP.n119 4.5005
R47975 VINP.n378 VINP.n119 4.5005
R47976 VINP.n226 VINP.n119 4.5005
R47977 VINP.n380 VINP.n119 4.5005
R47978 VINP.n225 VINP.n119 4.5005
R47979 VINP.n382 VINP.n119 4.5005
R47980 VINP.n224 VINP.n119 4.5005
R47981 VINP.n384 VINP.n119 4.5005
R47982 VINP.n223 VINP.n119 4.5005
R47983 VINP.n386 VINP.n119 4.5005
R47984 VINP.n222 VINP.n119 4.5005
R47985 VINP.n388 VINP.n119 4.5005
R47986 VINP.n221 VINP.n119 4.5005
R47987 VINP.n390 VINP.n119 4.5005
R47988 VINP.n220 VINP.n119 4.5005
R47989 VINP.n392 VINP.n119 4.5005
R47990 VINP.n219 VINP.n119 4.5005
R47991 VINP.n394 VINP.n119 4.5005
R47992 VINP.n218 VINP.n119 4.5005
R47993 VINP.n396 VINP.n119 4.5005
R47994 VINP.n217 VINP.n119 4.5005
R47995 VINP.n398 VINP.n119 4.5005
R47996 VINP.n216 VINP.n119 4.5005
R47997 VINP.n400 VINP.n119 4.5005
R47998 VINP.n215 VINP.n119 4.5005
R47999 VINP.n654 VINP.n119 4.5005
R48000 VINP.n656 VINP.n119 4.5005
R48001 VINP.n119 VINP.n0 4.5005
R48002 VINP.n278 VINP.n182 4.5005
R48003 VINP.n276 VINP.n182 4.5005
R48004 VINP.n280 VINP.n182 4.5005
R48005 VINP.n275 VINP.n182 4.5005
R48006 VINP.n282 VINP.n182 4.5005
R48007 VINP.n274 VINP.n182 4.5005
R48008 VINP.n284 VINP.n182 4.5005
R48009 VINP.n273 VINP.n182 4.5005
R48010 VINP.n286 VINP.n182 4.5005
R48011 VINP.n272 VINP.n182 4.5005
R48012 VINP.n288 VINP.n182 4.5005
R48013 VINP.n271 VINP.n182 4.5005
R48014 VINP.n290 VINP.n182 4.5005
R48015 VINP.n270 VINP.n182 4.5005
R48016 VINP.n292 VINP.n182 4.5005
R48017 VINP.n269 VINP.n182 4.5005
R48018 VINP.n294 VINP.n182 4.5005
R48019 VINP.n268 VINP.n182 4.5005
R48020 VINP.n296 VINP.n182 4.5005
R48021 VINP.n267 VINP.n182 4.5005
R48022 VINP.n298 VINP.n182 4.5005
R48023 VINP.n266 VINP.n182 4.5005
R48024 VINP.n300 VINP.n182 4.5005
R48025 VINP.n265 VINP.n182 4.5005
R48026 VINP.n302 VINP.n182 4.5005
R48027 VINP.n264 VINP.n182 4.5005
R48028 VINP.n304 VINP.n182 4.5005
R48029 VINP.n263 VINP.n182 4.5005
R48030 VINP.n306 VINP.n182 4.5005
R48031 VINP.n262 VINP.n182 4.5005
R48032 VINP.n308 VINP.n182 4.5005
R48033 VINP.n261 VINP.n182 4.5005
R48034 VINP.n310 VINP.n182 4.5005
R48035 VINP.n260 VINP.n182 4.5005
R48036 VINP.n312 VINP.n182 4.5005
R48037 VINP.n259 VINP.n182 4.5005
R48038 VINP.n314 VINP.n182 4.5005
R48039 VINP.n258 VINP.n182 4.5005
R48040 VINP.n316 VINP.n182 4.5005
R48041 VINP.n257 VINP.n182 4.5005
R48042 VINP.n318 VINP.n182 4.5005
R48043 VINP.n256 VINP.n182 4.5005
R48044 VINP.n320 VINP.n182 4.5005
R48045 VINP.n255 VINP.n182 4.5005
R48046 VINP.n322 VINP.n182 4.5005
R48047 VINP.n254 VINP.n182 4.5005
R48048 VINP.n324 VINP.n182 4.5005
R48049 VINP.n253 VINP.n182 4.5005
R48050 VINP.n326 VINP.n182 4.5005
R48051 VINP.n252 VINP.n182 4.5005
R48052 VINP.n328 VINP.n182 4.5005
R48053 VINP.n251 VINP.n182 4.5005
R48054 VINP.n330 VINP.n182 4.5005
R48055 VINP.n250 VINP.n182 4.5005
R48056 VINP.n332 VINP.n182 4.5005
R48057 VINP.n249 VINP.n182 4.5005
R48058 VINP.n334 VINP.n182 4.5005
R48059 VINP.n248 VINP.n182 4.5005
R48060 VINP.n336 VINP.n182 4.5005
R48061 VINP.n247 VINP.n182 4.5005
R48062 VINP.n338 VINP.n182 4.5005
R48063 VINP.n246 VINP.n182 4.5005
R48064 VINP.n340 VINP.n182 4.5005
R48065 VINP.n245 VINP.n182 4.5005
R48066 VINP.n342 VINP.n182 4.5005
R48067 VINP.n244 VINP.n182 4.5005
R48068 VINP.n344 VINP.n182 4.5005
R48069 VINP.n243 VINP.n182 4.5005
R48070 VINP.n346 VINP.n182 4.5005
R48071 VINP.n242 VINP.n182 4.5005
R48072 VINP.n348 VINP.n182 4.5005
R48073 VINP.n241 VINP.n182 4.5005
R48074 VINP.n350 VINP.n182 4.5005
R48075 VINP.n240 VINP.n182 4.5005
R48076 VINP.n352 VINP.n182 4.5005
R48077 VINP.n239 VINP.n182 4.5005
R48078 VINP.n354 VINP.n182 4.5005
R48079 VINP.n238 VINP.n182 4.5005
R48080 VINP.n356 VINP.n182 4.5005
R48081 VINP.n237 VINP.n182 4.5005
R48082 VINP.n358 VINP.n182 4.5005
R48083 VINP.n236 VINP.n182 4.5005
R48084 VINP.n360 VINP.n182 4.5005
R48085 VINP.n235 VINP.n182 4.5005
R48086 VINP.n362 VINP.n182 4.5005
R48087 VINP.n234 VINP.n182 4.5005
R48088 VINP.n364 VINP.n182 4.5005
R48089 VINP.n233 VINP.n182 4.5005
R48090 VINP.n366 VINP.n182 4.5005
R48091 VINP.n232 VINP.n182 4.5005
R48092 VINP.n368 VINP.n182 4.5005
R48093 VINP.n231 VINP.n182 4.5005
R48094 VINP.n370 VINP.n182 4.5005
R48095 VINP.n230 VINP.n182 4.5005
R48096 VINP.n372 VINP.n182 4.5005
R48097 VINP.n229 VINP.n182 4.5005
R48098 VINP.n374 VINP.n182 4.5005
R48099 VINP.n228 VINP.n182 4.5005
R48100 VINP.n376 VINP.n182 4.5005
R48101 VINP.n227 VINP.n182 4.5005
R48102 VINP.n378 VINP.n182 4.5005
R48103 VINP.n226 VINP.n182 4.5005
R48104 VINP.n380 VINP.n182 4.5005
R48105 VINP.n225 VINP.n182 4.5005
R48106 VINP.n382 VINP.n182 4.5005
R48107 VINP.n224 VINP.n182 4.5005
R48108 VINP.n384 VINP.n182 4.5005
R48109 VINP.n223 VINP.n182 4.5005
R48110 VINP.n386 VINP.n182 4.5005
R48111 VINP.n222 VINP.n182 4.5005
R48112 VINP.n388 VINP.n182 4.5005
R48113 VINP.n221 VINP.n182 4.5005
R48114 VINP.n390 VINP.n182 4.5005
R48115 VINP.n220 VINP.n182 4.5005
R48116 VINP.n392 VINP.n182 4.5005
R48117 VINP.n219 VINP.n182 4.5005
R48118 VINP.n394 VINP.n182 4.5005
R48119 VINP.n218 VINP.n182 4.5005
R48120 VINP.n396 VINP.n182 4.5005
R48121 VINP.n217 VINP.n182 4.5005
R48122 VINP.n398 VINP.n182 4.5005
R48123 VINP.n216 VINP.n182 4.5005
R48124 VINP.n400 VINP.n182 4.5005
R48125 VINP.n215 VINP.n182 4.5005
R48126 VINP.n654 VINP.n182 4.5005
R48127 VINP.n656 VINP.n182 4.5005
R48128 VINP.n182 VINP.n0 4.5005
R48129 VINP.n278 VINP.n118 4.5005
R48130 VINP.n276 VINP.n118 4.5005
R48131 VINP.n280 VINP.n118 4.5005
R48132 VINP.n275 VINP.n118 4.5005
R48133 VINP.n282 VINP.n118 4.5005
R48134 VINP.n274 VINP.n118 4.5005
R48135 VINP.n284 VINP.n118 4.5005
R48136 VINP.n273 VINP.n118 4.5005
R48137 VINP.n286 VINP.n118 4.5005
R48138 VINP.n272 VINP.n118 4.5005
R48139 VINP.n288 VINP.n118 4.5005
R48140 VINP.n271 VINP.n118 4.5005
R48141 VINP.n290 VINP.n118 4.5005
R48142 VINP.n270 VINP.n118 4.5005
R48143 VINP.n292 VINP.n118 4.5005
R48144 VINP.n269 VINP.n118 4.5005
R48145 VINP.n294 VINP.n118 4.5005
R48146 VINP.n268 VINP.n118 4.5005
R48147 VINP.n296 VINP.n118 4.5005
R48148 VINP.n267 VINP.n118 4.5005
R48149 VINP.n298 VINP.n118 4.5005
R48150 VINP.n266 VINP.n118 4.5005
R48151 VINP.n300 VINP.n118 4.5005
R48152 VINP.n265 VINP.n118 4.5005
R48153 VINP.n302 VINP.n118 4.5005
R48154 VINP.n264 VINP.n118 4.5005
R48155 VINP.n304 VINP.n118 4.5005
R48156 VINP.n263 VINP.n118 4.5005
R48157 VINP.n306 VINP.n118 4.5005
R48158 VINP.n262 VINP.n118 4.5005
R48159 VINP.n308 VINP.n118 4.5005
R48160 VINP.n261 VINP.n118 4.5005
R48161 VINP.n310 VINP.n118 4.5005
R48162 VINP.n260 VINP.n118 4.5005
R48163 VINP.n312 VINP.n118 4.5005
R48164 VINP.n259 VINP.n118 4.5005
R48165 VINP.n314 VINP.n118 4.5005
R48166 VINP.n258 VINP.n118 4.5005
R48167 VINP.n316 VINP.n118 4.5005
R48168 VINP.n257 VINP.n118 4.5005
R48169 VINP.n318 VINP.n118 4.5005
R48170 VINP.n256 VINP.n118 4.5005
R48171 VINP.n320 VINP.n118 4.5005
R48172 VINP.n255 VINP.n118 4.5005
R48173 VINP.n322 VINP.n118 4.5005
R48174 VINP.n254 VINP.n118 4.5005
R48175 VINP.n324 VINP.n118 4.5005
R48176 VINP.n253 VINP.n118 4.5005
R48177 VINP.n326 VINP.n118 4.5005
R48178 VINP.n252 VINP.n118 4.5005
R48179 VINP.n328 VINP.n118 4.5005
R48180 VINP.n251 VINP.n118 4.5005
R48181 VINP.n330 VINP.n118 4.5005
R48182 VINP.n250 VINP.n118 4.5005
R48183 VINP.n332 VINP.n118 4.5005
R48184 VINP.n249 VINP.n118 4.5005
R48185 VINP.n334 VINP.n118 4.5005
R48186 VINP.n248 VINP.n118 4.5005
R48187 VINP.n336 VINP.n118 4.5005
R48188 VINP.n247 VINP.n118 4.5005
R48189 VINP.n338 VINP.n118 4.5005
R48190 VINP.n246 VINP.n118 4.5005
R48191 VINP.n340 VINP.n118 4.5005
R48192 VINP.n245 VINP.n118 4.5005
R48193 VINP.n342 VINP.n118 4.5005
R48194 VINP.n244 VINP.n118 4.5005
R48195 VINP.n344 VINP.n118 4.5005
R48196 VINP.n243 VINP.n118 4.5005
R48197 VINP.n346 VINP.n118 4.5005
R48198 VINP.n242 VINP.n118 4.5005
R48199 VINP.n348 VINP.n118 4.5005
R48200 VINP.n241 VINP.n118 4.5005
R48201 VINP.n350 VINP.n118 4.5005
R48202 VINP.n240 VINP.n118 4.5005
R48203 VINP.n352 VINP.n118 4.5005
R48204 VINP.n239 VINP.n118 4.5005
R48205 VINP.n354 VINP.n118 4.5005
R48206 VINP.n238 VINP.n118 4.5005
R48207 VINP.n356 VINP.n118 4.5005
R48208 VINP.n237 VINP.n118 4.5005
R48209 VINP.n358 VINP.n118 4.5005
R48210 VINP.n236 VINP.n118 4.5005
R48211 VINP.n360 VINP.n118 4.5005
R48212 VINP.n235 VINP.n118 4.5005
R48213 VINP.n362 VINP.n118 4.5005
R48214 VINP.n234 VINP.n118 4.5005
R48215 VINP.n364 VINP.n118 4.5005
R48216 VINP.n233 VINP.n118 4.5005
R48217 VINP.n366 VINP.n118 4.5005
R48218 VINP.n232 VINP.n118 4.5005
R48219 VINP.n368 VINP.n118 4.5005
R48220 VINP.n231 VINP.n118 4.5005
R48221 VINP.n370 VINP.n118 4.5005
R48222 VINP.n230 VINP.n118 4.5005
R48223 VINP.n372 VINP.n118 4.5005
R48224 VINP.n229 VINP.n118 4.5005
R48225 VINP.n374 VINP.n118 4.5005
R48226 VINP.n228 VINP.n118 4.5005
R48227 VINP.n376 VINP.n118 4.5005
R48228 VINP.n227 VINP.n118 4.5005
R48229 VINP.n378 VINP.n118 4.5005
R48230 VINP.n226 VINP.n118 4.5005
R48231 VINP.n380 VINP.n118 4.5005
R48232 VINP.n225 VINP.n118 4.5005
R48233 VINP.n382 VINP.n118 4.5005
R48234 VINP.n224 VINP.n118 4.5005
R48235 VINP.n384 VINP.n118 4.5005
R48236 VINP.n223 VINP.n118 4.5005
R48237 VINP.n386 VINP.n118 4.5005
R48238 VINP.n222 VINP.n118 4.5005
R48239 VINP.n388 VINP.n118 4.5005
R48240 VINP.n221 VINP.n118 4.5005
R48241 VINP.n390 VINP.n118 4.5005
R48242 VINP.n220 VINP.n118 4.5005
R48243 VINP.n392 VINP.n118 4.5005
R48244 VINP.n219 VINP.n118 4.5005
R48245 VINP.n394 VINP.n118 4.5005
R48246 VINP.n218 VINP.n118 4.5005
R48247 VINP.n396 VINP.n118 4.5005
R48248 VINP.n217 VINP.n118 4.5005
R48249 VINP.n398 VINP.n118 4.5005
R48250 VINP.n216 VINP.n118 4.5005
R48251 VINP.n400 VINP.n118 4.5005
R48252 VINP.n215 VINP.n118 4.5005
R48253 VINP.n654 VINP.n118 4.5005
R48254 VINP.n656 VINP.n118 4.5005
R48255 VINP.n118 VINP.n0 4.5005
R48256 VINP.n278 VINP.n183 4.5005
R48257 VINP.n276 VINP.n183 4.5005
R48258 VINP.n280 VINP.n183 4.5005
R48259 VINP.n275 VINP.n183 4.5005
R48260 VINP.n282 VINP.n183 4.5005
R48261 VINP.n274 VINP.n183 4.5005
R48262 VINP.n284 VINP.n183 4.5005
R48263 VINP.n273 VINP.n183 4.5005
R48264 VINP.n286 VINP.n183 4.5005
R48265 VINP.n272 VINP.n183 4.5005
R48266 VINP.n288 VINP.n183 4.5005
R48267 VINP.n271 VINP.n183 4.5005
R48268 VINP.n290 VINP.n183 4.5005
R48269 VINP.n270 VINP.n183 4.5005
R48270 VINP.n292 VINP.n183 4.5005
R48271 VINP.n269 VINP.n183 4.5005
R48272 VINP.n294 VINP.n183 4.5005
R48273 VINP.n268 VINP.n183 4.5005
R48274 VINP.n296 VINP.n183 4.5005
R48275 VINP.n267 VINP.n183 4.5005
R48276 VINP.n298 VINP.n183 4.5005
R48277 VINP.n266 VINP.n183 4.5005
R48278 VINP.n300 VINP.n183 4.5005
R48279 VINP.n265 VINP.n183 4.5005
R48280 VINP.n302 VINP.n183 4.5005
R48281 VINP.n264 VINP.n183 4.5005
R48282 VINP.n304 VINP.n183 4.5005
R48283 VINP.n263 VINP.n183 4.5005
R48284 VINP.n306 VINP.n183 4.5005
R48285 VINP.n262 VINP.n183 4.5005
R48286 VINP.n308 VINP.n183 4.5005
R48287 VINP.n261 VINP.n183 4.5005
R48288 VINP.n310 VINP.n183 4.5005
R48289 VINP.n260 VINP.n183 4.5005
R48290 VINP.n312 VINP.n183 4.5005
R48291 VINP.n259 VINP.n183 4.5005
R48292 VINP.n314 VINP.n183 4.5005
R48293 VINP.n258 VINP.n183 4.5005
R48294 VINP.n316 VINP.n183 4.5005
R48295 VINP.n257 VINP.n183 4.5005
R48296 VINP.n318 VINP.n183 4.5005
R48297 VINP.n256 VINP.n183 4.5005
R48298 VINP.n320 VINP.n183 4.5005
R48299 VINP.n255 VINP.n183 4.5005
R48300 VINP.n322 VINP.n183 4.5005
R48301 VINP.n254 VINP.n183 4.5005
R48302 VINP.n324 VINP.n183 4.5005
R48303 VINP.n253 VINP.n183 4.5005
R48304 VINP.n326 VINP.n183 4.5005
R48305 VINP.n252 VINP.n183 4.5005
R48306 VINP.n328 VINP.n183 4.5005
R48307 VINP.n251 VINP.n183 4.5005
R48308 VINP.n330 VINP.n183 4.5005
R48309 VINP.n250 VINP.n183 4.5005
R48310 VINP.n332 VINP.n183 4.5005
R48311 VINP.n249 VINP.n183 4.5005
R48312 VINP.n334 VINP.n183 4.5005
R48313 VINP.n248 VINP.n183 4.5005
R48314 VINP.n336 VINP.n183 4.5005
R48315 VINP.n247 VINP.n183 4.5005
R48316 VINP.n338 VINP.n183 4.5005
R48317 VINP.n246 VINP.n183 4.5005
R48318 VINP.n340 VINP.n183 4.5005
R48319 VINP.n245 VINP.n183 4.5005
R48320 VINP.n342 VINP.n183 4.5005
R48321 VINP.n244 VINP.n183 4.5005
R48322 VINP.n344 VINP.n183 4.5005
R48323 VINP.n243 VINP.n183 4.5005
R48324 VINP.n346 VINP.n183 4.5005
R48325 VINP.n242 VINP.n183 4.5005
R48326 VINP.n348 VINP.n183 4.5005
R48327 VINP.n241 VINP.n183 4.5005
R48328 VINP.n350 VINP.n183 4.5005
R48329 VINP.n240 VINP.n183 4.5005
R48330 VINP.n352 VINP.n183 4.5005
R48331 VINP.n239 VINP.n183 4.5005
R48332 VINP.n354 VINP.n183 4.5005
R48333 VINP.n238 VINP.n183 4.5005
R48334 VINP.n356 VINP.n183 4.5005
R48335 VINP.n237 VINP.n183 4.5005
R48336 VINP.n358 VINP.n183 4.5005
R48337 VINP.n236 VINP.n183 4.5005
R48338 VINP.n360 VINP.n183 4.5005
R48339 VINP.n235 VINP.n183 4.5005
R48340 VINP.n362 VINP.n183 4.5005
R48341 VINP.n234 VINP.n183 4.5005
R48342 VINP.n364 VINP.n183 4.5005
R48343 VINP.n233 VINP.n183 4.5005
R48344 VINP.n366 VINP.n183 4.5005
R48345 VINP.n232 VINP.n183 4.5005
R48346 VINP.n368 VINP.n183 4.5005
R48347 VINP.n231 VINP.n183 4.5005
R48348 VINP.n370 VINP.n183 4.5005
R48349 VINP.n230 VINP.n183 4.5005
R48350 VINP.n372 VINP.n183 4.5005
R48351 VINP.n229 VINP.n183 4.5005
R48352 VINP.n374 VINP.n183 4.5005
R48353 VINP.n228 VINP.n183 4.5005
R48354 VINP.n376 VINP.n183 4.5005
R48355 VINP.n227 VINP.n183 4.5005
R48356 VINP.n378 VINP.n183 4.5005
R48357 VINP.n226 VINP.n183 4.5005
R48358 VINP.n380 VINP.n183 4.5005
R48359 VINP.n225 VINP.n183 4.5005
R48360 VINP.n382 VINP.n183 4.5005
R48361 VINP.n224 VINP.n183 4.5005
R48362 VINP.n384 VINP.n183 4.5005
R48363 VINP.n223 VINP.n183 4.5005
R48364 VINP.n386 VINP.n183 4.5005
R48365 VINP.n222 VINP.n183 4.5005
R48366 VINP.n388 VINP.n183 4.5005
R48367 VINP.n221 VINP.n183 4.5005
R48368 VINP.n390 VINP.n183 4.5005
R48369 VINP.n220 VINP.n183 4.5005
R48370 VINP.n392 VINP.n183 4.5005
R48371 VINP.n219 VINP.n183 4.5005
R48372 VINP.n394 VINP.n183 4.5005
R48373 VINP.n218 VINP.n183 4.5005
R48374 VINP.n396 VINP.n183 4.5005
R48375 VINP.n217 VINP.n183 4.5005
R48376 VINP.n398 VINP.n183 4.5005
R48377 VINP.n216 VINP.n183 4.5005
R48378 VINP.n400 VINP.n183 4.5005
R48379 VINP.n215 VINP.n183 4.5005
R48380 VINP.n654 VINP.n183 4.5005
R48381 VINP.n656 VINP.n183 4.5005
R48382 VINP.n183 VINP.n0 4.5005
R48383 VINP.n278 VINP.n117 4.5005
R48384 VINP.n276 VINP.n117 4.5005
R48385 VINP.n280 VINP.n117 4.5005
R48386 VINP.n275 VINP.n117 4.5005
R48387 VINP.n282 VINP.n117 4.5005
R48388 VINP.n274 VINP.n117 4.5005
R48389 VINP.n284 VINP.n117 4.5005
R48390 VINP.n273 VINP.n117 4.5005
R48391 VINP.n286 VINP.n117 4.5005
R48392 VINP.n272 VINP.n117 4.5005
R48393 VINP.n288 VINP.n117 4.5005
R48394 VINP.n271 VINP.n117 4.5005
R48395 VINP.n290 VINP.n117 4.5005
R48396 VINP.n270 VINP.n117 4.5005
R48397 VINP.n292 VINP.n117 4.5005
R48398 VINP.n269 VINP.n117 4.5005
R48399 VINP.n294 VINP.n117 4.5005
R48400 VINP.n268 VINP.n117 4.5005
R48401 VINP.n296 VINP.n117 4.5005
R48402 VINP.n267 VINP.n117 4.5005
R48403 VINP.n298 VINP.n117 4.5005
R48404 VINP.n266 VINP.n117 4.5005
R48405 VINP.n300 VINP.n117 4.5005
R48406 VINP.n265 VINP.n117 4.5005
R48407 VINP.n302 VINP.n117 4.5005
R48408 VINP.n264 VINP.n117 4.5005
R48409 VINP.n304 VINP.n117 4.5005
R48410 VINP.n263 VINP.n117 4.5005
R48411 VINP.n306 VINP.n117 4.5005
R48412 VINP.n262 VINP.n117 4.5005
R48413 VINP.n308 VINP.n117 4.5005
R48414 VINP.n261 VINP.n117 4.5005
R48415 VINP.n310 VINP.n117 4.5005
R48416 VINP.n260 VINP.n117 4.5005
R48417 VINP.n312 VINP.n117 4.5005
R48418 VINP.n259 VINP.n117 4.5005
R48419 VINP.n314 VINP.n117 4.5005
R48420 VINP.n258 VINP.n117 4.5005
R48421 VINP.n316 VINP.n117 4.5005
R48422 VINP.n257 VINP.n117 4.5005
R48423 VINP.n318 VINP.n117 4.5005
R48424 VINP.n256 VINP.n117 4.5005
R48425 VINP.n320 VINP.n117 4.5005
R48426 VINP.n255 VINP.n117 4.5005
R48427 VINP.n322 VINP.n117 4.5005
R48428 VINP.n254 VINP.n117 4.5005
R48429 VINP.n324 VINP.n117 4.5005
R48430 VINP.n253 VINP.n117 4.5005
R48431 VINP.n326 VINP.n117 4.5005
R48432 VINP.n252 VINP.n117 4.5005
R48433 VINP.n328 VINP.n117 4.5005
R48434 VINP.n251 VINP.n117 4.5005
R48435 VINP.n330 VINP.n117 4.5005
R48436 VINP.n250 VINP.n117 4.5005
R48437 VINP.n332 VINP.n117 4.5005
R48438 VINP.n249 VINP.n117 4.5005
R48439 VINP.n334 VINP.n117 4.5005
R48440 VINP.n248 VINP.n117 4.5005
R48441 VINP.n336 VINP.n117 4.5005
R48442 VINP.n247 VINP.n117 4.5005
R48443 VINP.n338 VINP.n117 4.5005
R48444 VINP.n246 VINP.n117 4.5005
R48445 VINP.n340 VINP.n117 4.5005
R48446 VINP.n245 VINP.n117 4.5005
R48447 VINP.n342 VINP.n117 4.5005
R48448 VINP.n244 VINP.n117 4.5005
R48449 VINP.n344 VINP.n117 4.5005
R48450 VINP.n243 VINP.n117 4.5005
R48451 VINP.n346 VINP.n117 4.5005
R48452 VINP.n242 VINP.n117 4.5005
R48453 VINP.n348 VINP.n117 4.5005
R48454 VINP.n241 VINP.n117 4.5005
R48455 VINP.n350 VINP.n117 4.5005
R48456 VINP.n240 VINP.n117 4.5005
R48457 VINP.n352 VINP.n117 4.5005
R48458 VINP.n239 VINP.n117 4.5005
R48459 VINP.n354 VINP.n117 4.5005
R48460 VINP.n238 VINP.n117 4.5005
R48461 VINP.n356 VINP.n117 4.5005
R48462 VINP.n237 VINP.n117 4.5005
R48463 VINP.n358 VINP.n117 4.5005
R48464 VINP.n236 VINP.n117 4.5005
R48465 VINP.n360 VINP.n117 4.5005
R48466 VINP.n235 VINP.n117 4.5005
R48467 VINP.n362 VINP.n117 4.5005
R48468 VINP.n234 VINP.n117 4.5005
R48469 VINP.n364 VINP.n117 4.5005
R48470 VINP.n233 VINP.n117 4.5005
R48471 VINP.n366 VINP.n117 4.5005
R48472 VINP.n232 VINP.n117 4.5005
R48473 VINP.n368 VINP.n117 4.5005
R48474 VINP.n231 VINP.n117 4.5005
R48475 VINP.n370 VINP.n117 4.5005
R48476 VINP.n230 VINP.n117 4.5005
R48477 VINP.n372 VINP.n117 4.5005
R48478 VINP.n229 VINP.n117 4.5005
R48479 VINP.n374 VINP.n117 4.5005
R48480 VINP.n228 VINP.n117 4.5005
R48481 VINP.n376 VINP.n117 4.5005
R48482 VINP.n227 VINP.n117 4.5005
R48483 VINP.n378 VINP.n117 4.5005
R48484 VINP.n226 VINP.n117 4.5005
R48485 VINP.n380 VINP.n117 4.5005
R48486 VINP.n225 VINP.n117 4.5005
R48487 VINP.n382 VINP.n117 4.5005
R48488 VINP.n224 VINP.n117 4.5005
R48489 VINP.n384 VINP.n117 4.5005
R48490 VINP.n223 VINP.n117 4.5005
R48491 VINP.n386 VINP.n117 4.5005
R48492 VINP.n222 VINP.n117 4.5005
R48493 VINP.n388 VINP.n117 4.5005
R48494 VINP.n221 VINP.n117 4.5005
R48495 VINP.n390 VINP.n117 4.5005
R48496 VINP.n220 VINP.n117 4.5005
R48497 VINP.n392 VINP.n117 4.5005
R48498 VINP.n219 VINP.n117 4.5005
R48499 VINP.n394 VINP.n117 4.5005
R48500 VINP.n218 VINP.n117 4.5005
R48501 VINP.n396 VINP.n117 4.5005
R48502 VINP.n217 VINP.n117 4.5005
R48503 VINP.n398 VINP.n117 4.5005
R48504 VINP.n216 VINP.n117 4.5005
R48505 VINP.n400 VINP.n117 4.5005
R48506 VINP.n215 VINP.n117 4.5005
R48507 VINP.n654 VINP.n117 4.5005
R48508 VINP.n656 VINP.n117 4.5005
R48509 VINP.n117 VINP.n0 4.5005
R48510 VINP.n278 VINP.n184 4.5005
R48511 VINP.n276 VINP.n184 4.5005
R48512 VINP.n280 VINP.n184 4.5005
R48513 VINP.n275 VINP.n184 4.5005
R48514 VINP.n282 VINP.n184 4.5005
R48515 VINP.n274 VINP.n184 4.5005
R48516 VINP.n284 VINP.n184 4.5005
R48517 VINP.n273 VINP.n184 4.5005
R48518 VINP.n286 VINP.n184 4.5005
R48519 VINP.n272 VINP.n184 4.5005
R48520 VINP.n288 VINP.n184 4.5005
R48521 VINP.n271 VINP.n184 4.5005
R48522 VINP.n290 VINP.n184 4.5005
R48523 VINP.n270 VINP.n184 4.5005
R48524 VINP.n292 VINP.n184 4.5005
R48525 VINP.n269 VINP.n184 4.5005
R48526 VINP.n294 VINP.n184 4.5005
R48527 VINP.n268 VINP.n184 4.5005
R48528 VINP.n296 VINP.n184 4.5005
R48529 VINP.n267 VINP.n184 4.5005
R48530 VINP.n298 VINP.n184 4.5005
R48531 VINP.n266 VINP.n184 4.5005
R48532 VINP.n300 VINP.n184 4.5005
R48533 VINP.n265 VINP.n184 4.5005
R48534 VINP.n302 VINP.n184 4.5005
R48535 VINP.n264 VINP.n184 4.5005
R48536 VINP.n304 VINP.n184 4.5005
R48537 VINP.n263 VINP.n184 4.5005
R48538 VINP.n306 VINP.n184 4.5005
R48539 VINP.n262 VINP.n184 4.5005
R48540 VINP.n308 VINP.n184 4.5005
R48541 VINP.n261 VINP.n184 4.5005
R48542 VINP.n310 VINP.n184 4.5005
R48543 VINP.n260 VINP.n184 4.5005
R48544 VINP.n312 VINP.n184 4.5005
R48545 VINP.n259 VINP.n184 4.5005
R48546 VINP.n314 VINP.n184 4.5005
R48547 VINP.n258 VINP.n184 4.5005
R48548 VINP.n316 VINP.n184 4.5005
R48549 VINP.n257 VINP.n184 4.5005
R48550 VINP.n318 VINP.n184 4.5005
R48551 VINP.n256 VINP.n184 4.5005
R48552 VINP.n320 VINP.n184 4.5005
R48553 VINP.n255 VINP.n184 4.5005
R48554 VINP.n322 VINP.n184 4.5005
R48555 VINP.n254 VINP.n184 4.5005
R48556 VINP.n324 VINP.n184 4.5005
R48557 VINP.n253 VINP.n184 4.5005
R48558 VINP.n326 VINP.n184 4.5005
R48559 VINP.n252 VINP.n184 4.5005
R48560 VINP.n328 VINP.n184 4.5005
R48561 VINP.n251 VINP.n184 4.5005
R48562 VINP.n330 VINP.n184 4.5005
R48563 VINP.n250 VINP.n184 4.5005
R48564 VINP.n332 VINP.n184 4.5005
R48565 VINP.n249 VINP.n184 4.5005
R48566 VINP.n334 VINP.n184 4.5005
R48567 VINP.n248 VINP.n184 4.5005
R48568 VINP.n336 VINP.n184 4.5005
R48569 VINP.n247 VINP.n184 4.5005
R48570 VINP.n338 VINP.n184 4.5005
R48571 VINP.n246 VINP.n184 4.5005
R48572 VINP.n340 VINP.n184 4.5005
R48573 VINP.n245 VINP.n184 4.5005
R48574 VINP.n342 VINP.n184 4.5005
R48575 VINP.n244 VINP.n184 4.5005
R48576 VINP.n344 VINP.n184 4.5005
R48577 VINP.n243 VINP.n184 4.5005
R48578 VINP.n346 VINP.n184 4.5005
R48579 VINP.n242 VINP.n184 4.5005
R48580 VINP.n348 VINP.n184 4.5005
R48581 VINP.n241 VINP.n184 4.5005
R48582 VINP.n350 VINP.n184 4.5005
R48583 VINP.n240 VINP.n184 4.5005
R48584 VINP.n352 VINP.n184 4.5005
R48585 VINP.n239 VINP.n184 4.5005
R48586 VINP.n354 VINP.n184 4.5005
R48587 VINP.n238 VINP.n184 4.5005
R48588 VINP.n356 VINP.n184 4.5005
R48589 VINP.n237 VINP.n184 4.5005
R48590 VINP.n358 VINP.n184 4.5005
R48591 VINP.n236 VINP.n184 4.5005
R48592 VINP.n360 VINP.n184 4.5005
R48593 VINP.n235 VINP.n184 4.5005
R48594 VINP.n362 VINP.n184 4.5005
R48595 VINP.n234 VINP.n184 4.5005
R48596 VINP.n364 VINP.n184 4.5005
R48597 VINP.n233 VINP.n184 4.5005
R48598 VINP.n366 VINP.n184 4.5005
R48599 VINP.n232 VINP.n184 4.5005
R48600 VINP.n368 VINP.n184 4.5005
R48601 VINP.n231 VINP.n184 4.5005
R48602 VINP.n370 VINP.n184 4.5005
R48603 VINP.n230 VINP.n184 4.5005
R48604 VINP.n372 VINP.n184 4.5005
R48605 VINP.n229 VINP.n184 4.5005
R48606 VINP.n374 VINP.n184 4.5005
R48607 VINP.n228 VINP.n184 4.5005
R48608 VINP.n376 VINP.n184 4.5005
R48609 VINP.n227 VINP.n184 4.5005
R48610 VINP.n378 VINP.n184 4.5005
R48611 VINP.n226 VINP.n184 4.5005
R48612 VINP.n380 VINP.n184 4.5005
R48613 VINP.n225 VINP.n184 4.5005
R48614 VINP.n382 VINP.n184 4.5005
R48615 VINP.n224 VINP.n184 4.5005
R48616 VINP.n384 VINP.n184 4.5005
R48617 VINP.n223 VINP.n184 4.5005
R48618 VINP.n386 VINP.n184 4.5005
R48619 VINP.n222 VINP.n184 4.5005
R48620 VINP.n388 VINP.n184 4.5005
R48621 VINP.n221 VINP.n184 4.5005
R48622 VINP.n390 VINP.n184 4.5005
R48623 VINP.n220 VINP.n184 4.5005
R48624 VINP.n392 VINP.n184 4.5005
R48625 VINP.n219 VINP.n184 4.5005
R48626 VINP.n394 VINP.n184 4.5005
R48627 VINP.n218 VINP.n184 4.5005
R48628 VINP.n396 VINP.n184 4.5005
R48629 VINP.n217 VINP.n184 4.5005
R48630 VINP.n398 VINP.n184 4.5005
R48631 VINP.n216 VINP.n184 4.5005
R48632 VINP.n400 VINP.n184 4.5005
R48633 VINP.n215 VINP.n184 4.5005
R48634 VINP.n654 VINP.n184 4.5005
R48635 VINP.n656 VINP.n184 4.5005
R48636 VINP.n184 VINP.n0 4.5005
R48637 VINP.n278 VINP.n116 4.5005
R48638 VINP.n276 VINP.n116 4.5005
R48639 VINP.n280 VINP.n116 4.5005
R48640 VINP.n275 VINP.n116 4.5005
R48641 VINP.n282 VINP.n116 4.5005
R48642 VINP.n274 VINP.n116 4.5005
R48643 VINP.n284 VINP.n116 4.5005
R48644 VINP.n273 VINP.n116 4.5005
R48645 VINP.n286 VINP.n116 4.5005
R48646 VINP.n272 VINP.n116 4.5005
R48647 VINP.n288 VINP.n116 4.5005
R48648 VINP.n271 VINP.n116 4.5005
R48649 VINP.n290 VINP.n116 4.5005
R48650 VINP.n270 VINP.n116 4.5005
R48651 VINP.n292 VINP.n116 4.5005
R48652 VINP.n269 VINP.n116 4.5005
R48653 VINP.n294 VINP.n116 4.5005
R48654 VINP.n268 VINP.n116 4.5005
R48655 VINP.n296 VINP.n116 4.5005
R48656 VINP.n267 VINP.n116 4.5005
R48657 VINP.n298 VINP.n116 4.5005
R48658 VINP.n266 VINP.n116 4.5005
R48659 VINP.n300 VINP.n116 4.5005
R48660 VINP.n265 VINP.n116 4.5005
R48661 VINP.n302 VINP.n116 4.5005
R48662 VINP.n264 VINP.n116 4.5005
R48663 VINP.n304 VINP.n116 4.5005
R48664 VINP.n263 VINP.n116 4.5005
R48665 VINP.n306 VINP.n116 4.5005
R48666 VINP.n262 VINP.n116 4.5005
R48667 VINP.n308 VINP.n116 4.5005
R48668 VINP.n261 VINP.n116 4.5005
R48669 VINP.n310 VINP.n116 4.5005
R48670 VINP.n260 VINP.n116 4.5005
R48671 VINP.n312 VINP.n116 4.5005
R48672 VINP.n259 VINP.n116 4.5005
R48673 VINP.n314 VINP.n116 4.5005
R48674 VINP.n258 VINP.n116 4.5005
R48675 VINP.n316 VINP.n116 4.5005
R48676 VINP.n257 VINP.n116 4.5005
R48677 VINP.n318 VINP.n116 4.5005
R48678 VINP.n256 VINP.n116 4.5005
R48679 VINP.n320 VINP.n116 4.5005
R48680 VINP.n255 VINP.n116 4.5005
R48681 VINP.n322 VINP.n116 4.5005
R48682 VINP.n254 VINP.n116 4.5005
R48683 VINP.n324 VINP.n116 4.5005
R48684 VINP.n253 VINP.n116 4.5005
R48685 VINP.n326 VINP.n116 4.5005
R48686 VINP.n252 VINP.n116 4.5005
R48687 VINP.n328 VINP.n116 4.5005
R48688 VINP.n251 VINP.n116 4.5005
R48689 VINP.n330 VINP.n116 4.5005
R48690 VINP.n250 VINP.n116 4.5005
R48691 VINP.n332 VINP.n116 4.5005
R48692 VINP.n249 VINP.n116 4.5005
R48693 VINP.n334 VINP.n116 4.5005
R48694 VINP.n248 VINP.n116 4.5005
R48695 VINP.n336 VINP.n116 4.5005
R48696 VINP.n247 VINP.n116 4.5005
R48697 VINP.n338 VINP.n116 4.5005
R48698 VINP.n246 VINP.n116 4.5005
R48699 VINP.n340 VINP.n116 4.5005
R48700 VINP.n245 VINP.n116 4.5005
R48701 VINP.n342 VINP.n116 4.5005
R48702 VINP.n244 VINP.n116 4.5005
R48703 VINP.n344 VINP.n116 4.5005
R48704 VINP.n243 VINP.n116 4.5005
R48705 VINP.n346 VINP.n116 4.5005
R48706 VINP.n242 VINP.n116 4.5005
R48707 VINP.n348 VINP.n116 4.5005
R48708 VINP.n241 VINP.n116 4.5005
R48709 VINP.n350 VINP.n116 4.5005
R48710 VINP.n240 VINP.n116 4.5005
R48711 VINP.n352 VINP.n116 4.5005
R48712 VINP.n239 VINP.n116 4.5005
R48713 VINP.n354 VINP.n116 4.5005
R48714 VINP.n238 VINP.n116 4.5005
R48715 VINP.n356 VINP.n116 4.5005
R48716 VINP.n237 VINP.n116 4.5005
R48717 VINP.n358 VINP.n116 4.5005
R48718 VINP.n236 VINP.n116 4.5005
R48719 VINP.n360 VINP.n116 4.5005
R48720 VINP.n235 VINP.n116 4.5005
R48721 VINP.n362 VINP.n116 4.5005
R48722 VINP.n234 VINP.n116 4.5005
R48723 VINP.n364 VINP.n116 4.5005
R48724 VINP.n233 VINP.n116 4.5005
R48725 VINP.n366 VINP.n116 4.5005
R48726 VINP.n232 VINP.n116 4.5005
R48727 VINP.n368 VINP.n116 4.5005
R48728 VINP.n231 VINP.n116 4.5005
R48729 VINP.n370 VINP.n116 4.5005
R48730 VINP.n230 VINP.n116 4.5005
R48731 VINP.n372 VINP.n116 4.5005
R48732 VINP.n229 VINP.n116 4.5005
R48733 VINP.n374 VINP.n116 4.5005
R48734 VINP.n228 VINP.n116 4.5005
R48735 VINP.n376 VINP.n116 4.5005
R48736 VINP.n227 VINP.n116 4.5005
R48737 VINP.n378 VINP.n116 4.5005
R48738 VINP.n226 VINP.n116 4.5005
R48739 VINP.n380 VINP.n116 4.5005
R48740 VINP.n225 VINP.n116 4.5005
R48741 VINP.n382 VINP.n116 4.5005
R48742 VINP.n224 VINP.n116 4.5005
R48743 VINP.n384 VINP.n116 4.5005
R48744 VINP.n223 VINP.n116 4.5005
R48745 VINP.n386 VINP.n116 4.5005
R48746 VINP.n222 VINP.n116 4.5005
R48747 VINP.n388 VINP.n116 4.5005
R48748 VINP.n221 VINP.n116 4.5005
R48749 VINP.n390 VINP.n116 4.5005
R48750 VINP.n220 VINP.n116 4.5005
R48751 VINP.n392 VINP.n116 4.5005
R48752 VINP.n219 VINP.n116 4.5005
R48753 VINP.n394 VINP.n116 4.5005
R48754 VINP.n218 VINP.n116 4.5005
R48755 VINP.n396 VINP.n116 4.5005
R48756 VINP.n217 VINP.n116 4.5005
R48757 VINP.n398 VINP.n116 4.5005
R48758 VINP.n216 VINP.n116 4.5005
R48759 VINP.n400 VINP.n116 4.5005
R48760 VINP.n215 VINP.n116 4.5005
R48761 VINP.n654 VINP.n116 4.5005
R48762 VINP.n656 VINP.n116 4.5005
R48763 VINP.n116 VINP.n0 4.5005
R48764 VINP.n278 VINP.n185 4.5005
R48765 VINP.n276 VINP.n185 4.5005
R48766 VINP.n280 VINP.n185 4.5005
R48767 VINP.n275 VINP.n185 4.5005
R48768 VINP.n282 VINP.n185 4.5005
R48769 VINP.n274 VINP.n185 4.5005
R48770 VINP.n284 VINP.n185 4.5005
R48771 VINP.n273 VINP.n185 4.5005
R48772 VINP.n286 VINP.n185 4.5005
R48773 VINP.n272 VINP.n185 4.5005
R48774 VINP.n288 VINP.n185 4.5005
R48775 VINP.n271 VINP.n185 4.5005
R48776 VINP.n290 VINP.n185 4.5005
R48777 VINP.n270 VINP.n185 4.5005
R48778 VINP.n292 VINP.n185 4.5005
R48779 VINP.n269 VINP.n185 4.5005
R48780 VINP.n294 VINP.n185 4.5005
R48781 VINP.n268 VINP.n185 4.5005
R48782 VINP.n296 VINP.n185 4.5005
R48783 VINP.n267 VINP.n185 4.5005
R48784 VINP.n298 VINP.n185 4.5005
R48785 VINP.n266 VINP.n185 4.5005
R48786 VINP.n300 VINP.n185 4.5005
R48787 VINP.n265 VINP.n185 4.5005
R48788 VINP.n302 VINP.n185 4.5005
R48789 VINP.n264 VINP.n185 4.5005
R48790 VINP.n304 VINP.n185 4.5005
R48791 VINP.n263 VINP.n185 4.5005
R48792 VINP.n306 VINP.n185 4.5005
R48793 VINP.n262 VINP.n185 4.5005
R48794 VINP.n308 VINP.n185 4.5005
R48795 VINP.n261 VINP.n185 4.5005
R48796 VINP.n310 VINP.n185 4.5005
R48797 VINP.n260 VINP.n185 4.5005
R48798 VINP.n312 VINP.n185 4.5005
R48799 VINP.n259 VINP.n185 4.5005
R48800 VINP.n314 VINP.n185 4.5005
R48801 VINP.n258 VINP.n185 4.5005
R48802 VINP.n316 VINP.n185 4.5005
R48803 VINP.n257 VINP.n185 4.5005
R48804 VINP.n318 VINP.n185 4.5005
R48805 VINP.n256 VINP.n185 4.5005
R48806 VINP.n320 VINP.n185 4.5005
R48807 VINP.n255 VINP.n185 4.5005
R48808 VINP.n322 VINP.n185 4.5005
R48809 VINP.n254 VINP.n185 4.5005
R48810 VINP.n324 VINP.n185 4.5005
R48811 VINP.n253 VINP.n185 4.5005
R48812 VINP.n326 VINP.n185 4.5005
R48813 VINP.n252 VINP.n185 4.5005
R48814 VINP.n328 VINP.n185 4.5005
R48815 VINP.n251 VINP.n185 4.5005
R48816 VINP.n330 VINP.n185 4.5005
R48817 VINP.n250 VINP.n185 4.5005
R48818 VINP.n332 VINP.n185 4.5005
R48819 VINP.n249 VINP.n185 4.5005
R48820 VINP.n334 VINP.n185 4.5005
R48821 VINP.n248 VINP.n185 4.5005
R48822 VINP.n336 VINP.n185 4.5005
R48823 VINP.n247 VINP.n185 4.5005
R48824 VINP.n338 VINP.n185 4.5005
R48825 VINP.n246 VINP.n185 4.5005
R48826 VINP.n340 VINP.n185 4.5005
R48827 VINP.n245 VINP.n185 4.5005
R48828 VINP.n342 VINP.n185 4.5005
R48829 VINP.n244 VINP.n185 4.5005
R48830 VINP.n344 VINP.n185 4.5005
R48831 VINP.n243 VINP.n185 4.5005
R48832 VINP.n346 VINP.n185 4.5005
R48833 VINP.n242 VINP.n185 4.5005
R48834 VINP.n348 VINP.n185 4.5005
R48835 VINP.n241 VINP.n185 4.5005
R48836 VINP.n350 VINP.n185 4.5005
R48837 VINP.n240 VINP.n185 4.5005
R48838 VINP.n352 VINP.n185 4.5005
R48839 VINP.n239 VINP.n185 4.5005
R48840 VINP.n354 VINP.n185 4.5005
R48841 VINP.n238 VINP.n185 4.5005
R48842 VINP.n356 VINP.n185 4.5005
R48843 VINP.n237 VINP.n185 4.5005
R48844 VINP.n358 VINP.n185 4.5005
R48845 VINP.n236 VINP.n185 4.5005
R48846 VINP.n360 VINP.n185 4.5005
R48847 VINP.n235 VINP.n185 4.5005
R48848 VINP.n362 VINP.n185 4.5005
R48849 VINP.n234 VINP.n185 4.5005
R48850 VINP.n364 VINP.n185 4.5005
R48851 VINP.n233 VINP.n185 4.5005
R48852 VINP.n366 VINP.n185 4.5005
R48853 VINP.n232 VINP.n185 4.5005
R48854 VINP.n368 VINP.n185 4.5005
R48855 VINP.n231 VINP.n185 4.5005
R48856 VINP.n370 VINP.n185 4.5005
R48857 VINP.n230 VINP.n185 4.5005
R48858 VINP.n372 VINP.n185 4.5005
R48859 VINP.n229 VINP.n185 4.5005
R48860 VINP.n374 VINP.n185 4.5005
R48861 VINP.n228 VINP.n185 4.5005
R48862 VINP.n376 VINP.n185 4.5005
R48863 VINP.n227 VINP.n185 4.5005
R48864 VINP.n378 VINP.n185 4.5005
R48865 VINP.n226 VINP.n185 4.5005
R48866 VINP.n380 VINP.n185 4.5005
R48867 VINP.n225 VINP.n185 4.5005
R48868 VINP.n382 VINP.n185 4.5005
R48869 VINP.n224 VINP.n185 4.5005
R48870 VINP.n384 VINP.n185 4.5005
R48871 VINP.n223 VINP.n185 4.5005
R48872 VINP.n386 VINP.n185 4.5005
R48873 VINP.n222 VINP.n185 4.5005
R48874 VINP.n388 VINP.n185 4.5005
R48875 VINP.n221 VINP.n185 4.5005
R48876 VINP.n390 VINP.n185 4.5005
R48877 VINP.n220 VINP.n185 4.5005
R48878 VINP.n392 VINP.n185 4.5005
R48879 VINP.n219 VINP.n185 4.5005
R48880 VINP.n394 VINP.n185 4.5005
R48881 VINP.n218 VINP.n185 4.5005
R48882 VINP.n396 VINP.n185 4.5005
R48883 VINP.n217 VINP.n185 4.5005
R48884 VINP.n398 VINP.n185 4.5005
R48885 VINP.n216 VINP.n185 4.5005
R48886 VINP.n400 VINP.n185 4.5005
R48887 VINP.n215 VINP.n185 4.5005
R48888 VINP.n654 VINP.n185 4.5005
R48889 VINP.n656 VINP.n185 4.5005
R48890 VINP.n185 VINP.n0 4.5005
R48891 VINP.n278 VINP.n115 4.5005
R48892 VINP.n276 VINP.n115 4.5005
R48893 VINP.n280 VINP.n115 4.5005
R48894 VINP.n275 VINP.n115 4.5005
R48895 VINP.n282 VINP.n115 4.5005
R48896 VINP.n274 VINP.n115 4.5005
R48897 VINP.n284 VINP.n115 4.5005
R48898 VINP.n273 VINP.n115 4.5005
R48899 VINP.n286 VINP.n115 4.5005
R48900 VINP.n272 VINP.n115 4.5005
R48901 VINP.n288 VINP.n115 4.5005
R48902 VINP.n271 VINP.n115 4.5005
R48903 VINP.n290 VINP.n115 4.5005
R48904 VINP.n270 VINP.n115 4.5005
R48905 VINP.n292 VINP.n115 4.5005
R48906 VINP.n269 VINP.n115 4.5005
R48907 VINP.n294 VINP.n115 4.5005
R48908 VINP.n268 VINP.n115 4.5005
R48909 VINP.n296 VINP.n115 4.5005
R48910 VINP.n267 VINP.n115 4.5005
R48911 VINP.n298 VINP.n115 4.5005
R48912 VINP.n266 VINP.n115 4.5005
R48913 VINP.n300 VINP.n115 4.5005
R48914 VINP.n265 VINP.n115 4.5005
R48915 VINP.n302 VINP.n115 4.5005
R48916 VINP.n264 VINP.n115 4.5005
R48917 VINP.n304 VINP.n115 4.5005
R48918 VINP.n263 VINP.n115 4.5005
R48919 VINP.n306 VINP.n115 4.5005
R48920 VINP.n262 VINP.n115 4.5005
R48921 VINP.n308 VINP.n115 4.5005
R48922 VINP.n261 VINP.n115 4.5005
R48923 VINP.n310 VINP.n115 4.5005
R48924 VINP.n260 VINP.n115 4.5005
R48925 VINP.n312 VINP.n115 4.5005
R48926 VINP.n259 VINP.n115 4.5005
R48927 VINP.n314 VINP.n115 4.5005
R48928 VINP.n258 VINP.n115 4.5005
R48929 VINP.n316 VINP.n115 4.5005
R48930 VINP.n257 VINP.n115 4.5005
R48931 VINP.n318 VINP.n115 4.5005
R48932 VINP.n256 VINP.n115 4.5005
R48933 VINP.n320 VINP.n115 4.5005
R48934 VINP.n255 VINP.n115 4.5005
R48935 VINP.n322 VINP.n115 4.5005
R48936 VINP.n254 VINP.n115 4.5005
R48937 VINP.n324 VINP.n115 4.5005
R48938 VINP.n253 VINP.n115 4.5005
R48939 VINP.n326 VINP.n115 4.5005
R48940 VINP.n252 VINP.n115 4.5005
R48941 VINP.n328 VINP.n115 4.5005
R48942 VINP.n251 VINP.n115 4.5005
R48943 VINP.n330 VINP.n115 4.5005
R48944 VINP.n250 VINP.n115 4.5005
R48945 VINP.n332 VINP.n115 4.5005
R48946 VINP.n249 VINP.n115 4.5005
R48947 VINP.n334 VINP.n115 4.5005
R48948 VINP.n248 VINP.n115 4.5005
R48949 VINP.n336 VINP.n115 4.5005
R48950 VINP.n247 VINP.n115 4.5005
R48951 VINP.n338 VINP.n115 4.5005
R48952 VINP.n246 VINP.n115 4.5005
R48953 VINP.n340 VINP.n115 4.5005
R48954 VINP.n245 VINP.n115 4.5005
R48955 VINP.n342 VINP.n115 4.5005
R48956 VINP.n244 VINP.n115 4.5005
R48957 VINP.n344 VINP.n115 4.5005
R48958 VINP.n243 VINP.n115 4.5005
R48959 VINP.n346 VINP.n115 4.5005
R48960 VINP.n242 VINP.n115 4.5005
R48961 VINP.n348 VINP.n115 4.5005
R48962 VINP.n241 VINP.n115 4.5005
R48963 VINP.n350 VINP.n115 4.5005
R48964 VINP.n240 VINP.n115 4.5005
R48965 VINP.n352 VINP.n115 4.5005
R48966 VINP.n239 VINP.n115 4.5005
R48967 VINP.n354 VINP.n115 4.5005
R48968 VINP.n238 VINP.n115 4.5005
R48969 VINP.n356 VINP.n115 4.5005
R48970 VINP.n237 VINP.n115 4.5005
R48971 VINP.n358 VINP.n115 4.5005
R48972 VINP.n236 VINP.n115 4.5005
R48973 VINP.n360 VINP.n115 4.5005
R48974 VINP.n235 VINP.n115 4.5005
R48975 VINP.n362 VINP.n115 4.5005
R48976 VINP.n234 VINP.n115 4.5005
R48977 VINP.n364 VINP.n115 4.5005
R48978 VINP.n233 VINP.n115 4.5005
R48979 VINP.n366 VINP.n115 4.5005
R48980 VINP.n232 VINP.n115 4.5005
R48981 VINP.n368 VINP.n115 4.5005
R48982 VINP.n231 VINP.n115 4.5005
R48983 VINP.n370 VINP.n115 4.5005
R48984 VINP.n230 VINP.n115 4.5005
R48985 VINP.n372 VINP.n115 4.5005
R48986 VINP.n229 VINP.n115 4.5005
R48987 VINP.n374 VINP.n115 4.5005
R48988 VINP.n228 VINP.n115 4.5005
R48989 VINP.n376 VINP.n115 4.5005
R48990 VINP.n227 VINP.n115 4.5005
R48991 VINP.n378 VINP.n115 4.5005
R48992 VINP.n226 VINP.n115 4.5005
R48993 VINP.n380 VINP.n115 4.5005
R48994 VINP.n225 VINP.n115 4.5005
R48995 VINP.n382 VINP.n115 4.5005
R48996 VINP.n224 VINP.n115 4.5005
R48997 VINP.n384 VINP.n115 4.5005
R48998 VINP.n223 VINP.n115 4.5005
R48999 VINP.n386 VINP.n115 4.5005
R49000 VINP.n222 VINP.n115 4.5005
R49001 VINP.n388 VINP.n115 4.5005
R49002 VINP.n221 VINP.n115 4.5005
R49003 VINP.n390 VINP.n115 4.5005
R49004 VINP.n220 VINP.n115 4.5005
R49005 VINP.n392 VINP.n115 4.5005
R49006 VINP.n219 VINP.n115 4.5005
R49007 VINP.n394 VINP.n115 4.5005
R49008 VINP.n218 VINP.n115 4.5005
R49009 VINP.n396 VINP.n115 4.5005
R49010 VINP.n217 VINP.n115 4.5005
R49011 VINP.n398 VINP.n115 4.5005
R49012 VINP.n216 VINP.n115 4.5005
R49013 VINP.n400 VINP.n115 4.5005
R49014 VINP.n215 VINP.n115 4.5005
R49015 VINP.n654 VINP.n115 4.5005
R49016 VINP.n656 VINP.n115 4.5005
R49017 VINP.n115 VINP.n0 4.5005
R49018 VINP.n278 VINP.n186 4.5005
R49019 VINP.n276 VINP.n186 4.5005
R49020 VINP.n280 VINP.n186 4.5005
R49021 VINP.n275 VINP.n186 4.5005
R49022 VINP.n282 VINP.n186 4.5005
R49023 VINP.n274 VINP.n186 4.5005
R49024 VINP.n284 VINP.n186 4.5005
R49025 VINP.n273 VINP.n186 4.5005
R49026 VINP.n286 VINP.n186 4.5005
R49027 VINP.n272 VINP.n186 4.5005
R49028 VINP.n288 VINP.n186 4.5005
R49029 VINP.n271 VINP.n186 4.5005
R49030 VINP.n290 VINP.n186 4.5005
R49031 VINP.n270 VINP.n186 4.5005
R49032 VINP.n292 VINP.n186 4.5005
R49033 VINP.n269 VINP.n186 4.5005
R49034 VINP.n294 VINP.n186 4.5005
R49035 VINP.n268 VINP.n186 4.5005
R49036 VINP.n296 VINP.n186 4.5005
R49037 VINP.n267 VINP.n186 4.5005
R49038 VINP.n298 VINP.n186 4.5005
R49039 VINP.n266 VINP.n186 4.5005
R49040 VINP.n300 VINP.n186 4.5005
R49041 VINP.n265 VINP.n186 4.5005
R49042 VINP.n302 VINP.n186 4.5005
R49043 VINP.n264 VINP.n186 4.5005
R49044 VINP.n304 VINP.n186 4.5005
R49045 VINP.n263 VINP.n186 4.5005
R49046 VINP.n306 VINP.n186 4.5005
R49047 VINP.n262 VINP.n186 4.5005
R49048 VINP.n308 VINP.n186 4.5005
R49049 VINP.n261 VINP.n186 4.5005
R49050 VINP.n310 VINP.n186 4.5005
R49051 VINP.n260 VINP.n186 4.5005
R49052 VINP.n312 VINP.n186 4.5005
R49053 VINP.n259 VINP.n186 4.5005
R49054 VINP.n314 VINP.n186 4.5005
R49055 VINP.n258 VINP.n186 4.5005
R49056 VINP.n316 VINP.n186 4.5005
R49057 VINP.n257 VINP.n186 4.5005
R49058 VINP.n318 VINP.n186 4.5005
R49059 VINP.n256 VINP.n186 4.5005
R49060 VINP.n320 VINP.n186 4.5005
R49061 VINP.n255 VINP.n186 4.5005
R49062 VINP.n322 VINP.n186 4.5005
R49063 VINP.n254 VINP.n186 4.5005
R49064 VINP.n324 VINP.n186 4.5005
R49065 VINP.n253 VINP.n186 4.5005
R49066 VINP.n326 VINP.n186 4.5005
R49067 VINP.n252 VINP.n186 4.5005
R49068 VINP.n328 VINP.n186 4.5005
R49069 VINP.n251 VINP.n186 4.5005
R49070 VINP.n330 VINP.n186 4.5005
R49071 VINP.n250 VINP.n186 4.5005
R49072 VINP.n332 VINP.n186 4.5005
R49073 VINP.n249 VINP.n186 4.5005
R49074 VINP.n334 VINP.n186 4.5005
R49075 VINP.n248 VINP.n186 4.5005
R49076 VINP.n336 VINP.n186 4.5005
R49077 VINP.n247 VINP.n186 4.5005
R49078 VINP.n338 VINP.n186 4.5005
R49079 VINP.n246 VINP.n186 4.5005
R49080 VINP.n340 VINP.n186 4.5005
R49081 VINP.n245 VINP.n186 4.5005
R49082 VINP.n342 VINP.n186 4.5005
R49083 VINP.n244 VINP.n186 4.5005
R49084 VINP.n344 VINP.n186 4.5005
R49085 VINP.n243 VINP.n186 4.5005
R49086 VINP.n346 VINP.n186 4.5005
R49087 VINP.n242 VINP.n186 4.5005
R49088 VINP.n348 VINP.n186 4.5005
R49089 VINP.n241 VINP.n186 4.5005
R49090 VINP.n350 VINP.n186 4.5005
R49091 VINP.n240 VINP.n186 4.5005
R49092 VINP.n352 VINP.n186 4.5005
R49093 VINP.n239 VINP.n186 4.5005
R49094 VINP.n354 VINP.n186 4.5005
R49095 VINP.n238 VINP.n186 4.5005
R49096 VINP.n356 VINP.n186 4.5005
R49097 VINP.n237 VINP.n186 4.5005
R49098 VINP.n358 VINP.n186 4.5005
R49099 VINP.n236 VINP.n186 4.5005
R49100 VINP.n360 VINP.n186 4.5005
R49101 VINP.n235 VINP.n186 4.5005
R49102 VINP.n362 VINP.n186 4.5005
R49103 VINP.n234 VINP.n186 4.5005
R49104 VINP.n364 VINP.n186 4.5005
R49105 VINP.n233 VINP.n186 4.5005
R49106 VINP.n366 VINP.n186 4.5005
R49107 VINP.n232 VINP.n186 4.5005
R49108 VINP.n368 VINP.n186 4.5005
R49109 VINP.n231 VINP.n186 4.5005
R49110 VINP.n370 VINP.n186 4.5005
R49111 VINP.n230 VINP.n186 4.5005
R49112 VINP.n372 VINP.n186 4.5005
R49113 VINP.n229 VINP.n186 4.5005
R49114 VINP.n374 VINP.n186 4.5005
R49115 VINP.n228 VINP.n186 4.5005
R49116 VINP.n376 VINP.n186 4.5005
R49117 VINP.n227 VINP.n186 4.5005
R49118 VINP.n378 VINP.n186 4.5005
R49119 VINP.n226 VINP.n186 4.5005
R49120 VINP.n380 VINP.n186 4.5005
R49121 VINP.n225 VINP.n186 4.5005
R49122 VINP.n382 VINP.n186 4.5005
R49123 VINP.n224 VINP.n186 4.5005
R49124 VINP.n384 VINP.n186 4.5005
R49125 VINP.n223 VINP.n186 4.5005
R49126 VINP.n386 VINP.n186 4.5005
R49127 VINP.n222 VINP.n186 4.5005
R49128 VINP.n388 VINP.n186 4.5005
R49129 VINP.n221 VINP.n186 4.5005
R49130 VINP.n390 VINP.n186 4.5005
R49131 VINP.n220 VINP.n186 4.5005
R49132 VINP.n392 VINP.n186 4.5005
R49133 VINP.n219 VINP.n186 4.5005
R49134 VINP.n394 VINP.n186 4.5005
R49135 VINP.n218 VINP.n186 4.5005
R49136 VINP.n396 VINP.n186 4.5005
R49137 VINP.n217 VINP.n186 4.5005
R49138 VINP.n398 VINP.n186 4.5005
R49139 VINP.n216 VINP.n186 4.5005
R49140 VINP.n400 VINP.n186 4.5005
R49141 VINP.n215 VINP.n186 4.5005
R49142 VINP.n654 VINP.n186 4.5005
R49143 VINP.n656 VINP.n186 4.5005
R49144 VINP.n186 VINP.n0 4.5005
R49145 VINP.n278 VINP.n114 4.5005
R49146 VINP.n276 VINP.n114 4.5005
R49147 VINP.n280 VINP.n114 4.5005
R49148 VINP.n275 VINP.n114 4.5005
R49149 VINP.n282 VINP.n114 4.5005
R49150 VINP.n274 VINP.n114 4.5005
R49151 VINP.n284 VINP.n114 4.5005
R49152 VINP.n273 VINP.n114 4.5005
R49153 VINP.n286 VINP.n114 4.5005
R49154 VINP.n272 VINP.n114 4.5005
R49155 VINP.n288 VINP.n114 4.5005
R49156 VINP.n271 VINP.n114 4.5005
R49157 VINP.n290 VINP.n114 4.5005
R49158 VINP.n270 VINP.n114 4.5005
R49159 VINP.n292 VINP.n114 4.5005
R49160 VINP.n269 VINP.n114 4.5005
R49161 VINP.n294 VINP.n114 4.5005
R49162 VINP.n268 VINP.n114 4.5005
R49163 VINP.n296 VINP.n114 4.5005
R49164 VINP.n267 VINP.n114 4.5005
R49165 VINP.n298 VINP.n114 4.5005
R49166 VINP.n266 VINP.n114 4.5005
R49167 VINP.n300 VINP.n114 4.5005
R49168 VINP.n265 VINP.n114 4.5005
R49169 VINP.n302 VINP.n114 4.5005
R49170 VINP.n264 VINP.n114 4.5005
R49171 VINP.n304 VINP.n114 4.5005
R49172 VINP.n263 VINP.n114 4.5005
R49173 VINP.n306 VINP.n114 4.5005
R49174 VINP.n262 VINP.n114 4.5005
R49175 VINP.n308 VINP.n114 4.5005
R49176 VINP.n261 VINP.n114 4.5005
R49177 VINP.n310 VINP.n114 4.5005
R49178 VINP.n260 VINP.n114 4.5005
R49179 VINP.n312 VINP.n114 4.5005
R49180 VINP.n259 VINP.n114 4.5005
R49181 VINP.n314 VINP.n114 4.5005
R49182 VINP.n258 VINP.n114 4.5005
R49183 VINP.n316 VINP.n114 4.5005
R49184 VINP.n257 VINP.n114 4.5005
R49185 VINP.n318 VINP.n114 4.5005
R49186 VINP.n256 VINP.n114 4.5005
R49187 VINP.n320 VINP.n114 4.5005
R49188 VINP.n255 VINP.n114 4.5005
R49189 VINP.n322 VINP.n114 4.5005
R49190 VINP.n254 VINP.n114 4.5005
R49191 VINP.n324 VINP.n114 4.5005
R49192 VINP.n253 VINP.n114 4.5005
R49193 VINP.n326 VINP.n114 4.5005
R49194 VINP.n252 VINP.n114 4.5005
R49195 VINP.n328 VINP.n114 4.5005
R49196 VINP.n251 VINP.n114 4.5005
R49197 VINP.n330 VINP.n114 4.5005
R49198 VINP.n250 VINP.n114 4.5005
R49199 VINP.n332 VINP.n114 4.5005
R49200 VINP.n249 VINP.n114 4.5005
R49201 VINP.n334 VINP.n114 4.5005
R49202 VINP.n248 VINP.n114 4.5005
R49203 VINP.n336 VINP.n114 4.5005
R49204 VINP.n247 VINP.n114 4.5005
R49205 VINP.n338 VINP.n114 4.5005
R49206 VINP.n246 VINP.n114 4.5005
R49207 VINP.n340 VINP.n114 4.5005
R49208 VINP.n245 VINP.n114 4.5005
R49209 VINP.n342 VINP.n114 4.5005
R49210 VINP.n244 VINP.n114 4.5005
R49211 VINP.n344 VINP.n114 4.5005
R49212 VINP.n243 VINP.n114 4.5005
R49213 VINP.n346 VINP.n114 4.5005
R49214 VINP.n242 VINP.n114 4.5005
R49215 VINP.n348 VINP.n114 4.5005
R49216 VINP.n241 VINP.n114 4.5005
R49217 VINP.n350 VINP.n114 4.5005
R49218 VINP.n240 VINP.n114 4.5005
R49219 VINP.n352 VINP.n114 4.5005
R49220 VINP.n239 VINP.n114 4.5005
R49221 VINP.n354 VINP.n114 4.5005
R49222 VINP.n238 VINP.n114 4.5005
R49223 VINP.n356 VINP.n114 4.5005
R49224 VINP.n237 VINP.n114 4.5005
R49225 VINP.n358 VINP.n114 4.5005
R49226 VINP.n236 VINP.n114 4.5005
R49227 VINP.n360 VINP.n114 4.5005
R49228 VINP.n235 VINP.n114 4.5005
R49229 VINP.n362 VINP.n114 4.5005
R49230 VINP.n234 VINP.n114 4.5005
R49231 VINP.n364 VINP.n114 4.5005
R49232 VINP.n233 VINP.n114 4.5005
R49233 VINP.n366 VINP.n114 4.5005
R49234 VINP.n232 VINP.n114 4.5005
R49235 VINP.n368 VINP.n114 4.5005
R49236 VINP.n231 VINP.n114 4.5005
R49237 VINP.n370 VINP.n114 4.5005
R49238 VINP.n230 VINP.n114 4.5005
R49239 VINP.n372 VINP.n114 4.5005
R49240 VINP.n229 VINP.n114 4.5005
R49241 VINP.n374 VINP.n114 4.5005
R49242 VINP.n228 VINP.n114 4.5005
R49243 VINP.n376 VINP.n114 4.5005
R49244 VINP.n227 VINP.n114 4.5005
R49245 VINP.n378 VINP.n114 4.5005
R49246 VINP.n226 VINP.n114 4.5005
R49247 VINP.n380 VINP.n114 4.5005
R49248 VINP.n225 VINP.n114 4.5005
R49249 VINP.n382 VINP.n114 4.5005
R49250 VINP.n224 VINP.n114 4.5005
R49251 VINP.n384 VINP.n114 4.5005
R49252 VINP.n223 VINP.n114 4.5005
R49253 VINP.n386 VINP.n114 4.5005
R49254 VINP.n222 VINP.n114 4.5005
R49255 VINP.n388 VINP.n114 4.5005
R49256 VINP.n221 VINP.n114 4.5005
R49257 VINP.n390 VINP.n114 4.5005
R49258 VINP.n220 VINP.n114 4.5005
R49259 VINP.n392 VINP.n114 4.5005
R49260 VINP.n219 VINP.n114 4.5005
R49261 VINP.n394 VINP.n114 4.5005
R49262 VINP.n218 VINP.n114 4.5005
R49263 VINP.n396 VINP.n114 4.5005
R49264 VINP.n217 VINP.n114 4.5005
R49265 VINP.n398 VINP.n114 4.5005
R49266 VINP.n216 VINP.n114 4.5005
R49267 VINP.n400 VINP.n114 4.5005
R49268 VINP.n215 VINP.n114 4.5005
R49269 VINP.n654 VINP.n114 4.5005
R49270 VINP.n656 VINP.n114 4.5005
R49271 VINP.n114 VINP.n0 4.5005
R49272 VINP.n278 VINP.n187 4.5005
R49273 VINP.n276 VINP.n187 4.5005
R49274 VINP.n280 VINP.n187 4.5005
R49275 VINP.n275 VINP.n187 4.5005
R49276 VINP.n282 VINP.n187 4.5005
R49277 VINP.n274 VINP.n187 4.5005
R49278 VINP.n284 VINP.n187 4.5005
R49279 VINP.n273 VINP.n187 4.5005
R49280 VINP.n286 VINP.n187 4.5005
R49281 VINP.n272 VINP.n187 4.5005
R49282 VINP.n288 VINP.n187 4.5005
R49283 VINP.n271 VINP.n187 4.5005
R49284 VINP.n290 VINP.n187 4.5005
R49285 VINP.n270 VINP.n187 4.5005
R49286 VINP.n292 VINP.n187 4.5005
R49287 VINP.n269 VINP.n187 4.5005
R49288 VINP.n294 VINP.n187 4.5005
R49289 VINP.n268 VINP.n187 4.5005
R49290 VINP.n296 VINP.n187 4.5005
R49291 VINP.n267 VINP.n187 4.5005
R49292 VINP.n298 VINP.n187 4.5005
R49293 VINP.n266 VINP.n187 4.5005
R49294 VINP.n300 VINP.n187 4.5005
R49295 VINP.n265 VINP.n187 4.5005
R49296 VINP.n302 VINP.n187 4.5005
R49297 VINP.n264 VINP.n187 4.5005
R49298 VINP.n304 VINP.n187 4.5005
R49299 VINP.n263 VINP.n187 4.5005
R49300 VINP.n306 VINP.n187 4.5005
R49301 VINP.n262 VINP.n187 4.5005
R49302 VINP.n308 VINP.n187 4.5005
R49303 VINP.n261 VINP.n187 4.5005
R49304 VINP.n310 VINP.n187 4.5005
R49305 VINP.n260 VINP.n187 4.5005
R49306 VINP.n312 VINP.n187 4.5005
R49307 VINP.n259 VINP.n187 4.5005
R49308 VINP.n314 VINP.n187 4.5005
R49309 VINP.n258 VINP.n187 4.5005
R49310 VINP.n316 VINP.n187 4.5005
R49311 VINP.n257 VINP.n187 4.5005
R49312 VINP.n318 VINP.n187 4.5005
R49313 VINP.n256 VINP.n187 4.5005
R49314 VINP.n320 VINP.n187 4.5005
R49315 VINP.n255 VINP.n187 4.5005
R49316 VINP.n322 VINP.n187 4.5005
R49317 VINP.n254 VINP.n187 4.5005
R49318 VINP.n324 VINP.n187 4.5005
R49319 VINP.n253 VINP.n187 4.5005
R49320 VINP.n326 VINP.n187 4.5005
R49321 VINP.n252 VINP.n187 4.5005
R49322 VINP.n328 VINP.n187 4.5005
R49323 VINP.n251 VINP.n187 4.5005
R49324 VINP.n330 VINP.n187 4.5005
R49325 VINP.n250 VINP.n187 4.5005
R49326 VINP.n332 VINP.n187 4.5005
R49327 VINP.n249 VINP.n187 4.5005
R49328 VINP.n334 VINP.n187 4.5005
R49329 VINP.n248 VINP.n187 4.5005
R49330 VINP.n336 VINP.n187 4.5005
R49331 VINP.n247 VINP.n187 4.5005
R49332 VINP.n338 VINP.n187 4.5005
R49333 VINP.n246 VINP.n187 4.5005
R49334 VINP.n340 VINP.n187 4.5005
R49335 VINP.n245 VINP.n187 4.5005
R49336 VINP.n342 VINP.n187 4.5005
R49337 VINP.n244 VINP.n187 4.5005
R49338 VINP.n344 VINP.n187 4.5005
R49339 VINP.n243 VINP.n187 4.5005
R49340 VINP.n346 VINP.n187 4.5005
R49341 VINP.n242 VINP.n187 4.5005
R49342 VINP.n348 VINP.n187 4.5005
R49343 VINP.n241 VINP.n187 4.5005
R49344 VINP.n350 VINP.n187 4.5005
R49345 VINP.n240 VINP.n187 4.5005
R49346 VINP.n352 VINP.n187 4.5005
R49347 VINP.n239 VINP.n187 4.5005
R49348 VINP.n354 VINP.n187 4.5005
R49349 VINP.n238 VINP.n187 4.5005
R49350 VINP.n356 VINP.n187 4.5005
R49351 VINP.n237 VINP.n187 4.5005
R49352 VINP.n358 VINP.n187 4.5005
R49353 VINP.n236 VINP.n187 4.5005
R49354 VINP.n360 VINP.n187 4.5005
R49355 VINP.n235 VINP.n187 4.5005
R49356 VINP.n362 VINP.n187 4.5005
R49357 VINP.n234 VINP.n187 4.5005
R49358 VINP.n364 VINP.n187 4.5005
R49359 VINP.n233 VINP.n187 4.5005
R49360 VINP.n366 VINP.n187 4.5005
R49361 VINP.n232 VINP.n187 4.5005
R49362 VINP.n368 VINP.n187 4.5005
R49363 VINP.n231 VINP.n187 4.5005
R49364 VINP.n370 VINP.n187 4.5005
R49365 VINP.n230 VINP.n187 4.5005
R49366 VINP.n372 VINP.n187 4.5005
R49367 VINP.n229 VINP.n187 4.5005
R49368 VINP.n374 VINP.n187 4.5005
R49369 VINP.n228 VINP.n187 4.5005
R49370 VINP.n376 VINP.n187 4.5005
R49371 VINP.n227 VINP.n187 4.5005
R49372 VINP.n378 VINP.n187 4.5005
R49373 VINP.n226 VINP.n187 4.5005
R49374 VINP.n380 VINP.n187 4.5005
R49375 VINP.n225 VINP.n187 4.5005
R49376 VINP.n382 VINP.n187 4.5005
R49377 VINP.n224 VINP.n187 4.5005
R49378 VINP.n384 VINP.n187 4.5005
R49379 VINP.n223 VINP.n187 4.5005
R49380 VINP.n386 VINP.n187 4.5005
R49381 VINP.n222 VINP.n187 4.5005
R49382 VINP.n388 VINP.n187 4.5005
R49383 VINP.n221 VINP.n187 4.5005
R49384 VINP.n390 VINP.n187 4.5005
R49385 VINP.n220 VINP.n187 4.5005
R49386 VINP.n392 VINP.n187 4.5005
R49387 VINP.n219 VINP.n187 4.5005
R49388 VINP.n394 VINP.n187 4.5005
R49389 VINP.n218 VINP.n187 4.5005
R49390 VINP.n396 VINP.n187 4.5005
R49391 VINP.n217 VINP.n187 4.5005
R49392 VINP.n398 VINP.n187 4.5005
R49393 VINP.n216 VINP.n187 4.5005
R49394 VINP.n400 VINP.n187 4.5005
R49395 VINP.n215 VINP.n187 4.5005
R49396 VINP.n654 VINP.n187 4.5005
R49397 VINP.n656 VINP.n187 4.5005
R49398 VINP.n187 VINP.n0 4.5005
R49399 VINP.n278 VINP.n113 4.5005
R49400 VINP.n276 VINP.n113 4.5005
R49401 VINP.n280 VINP.n113 4.5005
R49402 VINP.n275 VINP.n113 4.5005
R49403 VINP.n282 VINP.n113 4.5005
R49404 VINP.n274 VINP.n113 4.5005
R49405 VINP.n284 VINP.n113 4.5005
R49406 VINP.n273 VINP.n113 4.5005
R49407 VINP.n286 VINP.n113 4.5005
R49408 VINP.n272 VINP.n113 4.5005
R49409 VINP.n288 VINP.n113 4.5005
R49410 VINP.n271 VINP.n113 4.5005
R49411 VINP.n290 VINP.n113 4.5005
R49412 VINP.n270 VINP.n113 4.5005
R49413 VINP.n292 VINP.n113 4.5005
R49414 VINP.n269 VINP.n113 4.5005
R49415 VINP.n294 VINP.n113 4.5005
R49416 VINP.n268 VINP.n113 4.5005
R49417 VINP.n296 VINP.n113 4.5005
R49418 VINP.n267 VINP.n113 4.5005
R49419 VINP.n298 VINP.n113 4.5005
R49420 VINP.n266 VINP.n113 4.5005
R49421 VINP.n300 VINP.n113 4.5005
R49422 VINP.n265 VINP.n113 4.5005
R49423 VINP.n302 VINP.n113 4.5005
R49424 VINP.n264 VINP.n113 4.5005
R49425 VINP.n304 VINP.n113 4.5005
R49426 VINP.n263 VINP.n113 4.5005
R49427 VINP.n306 VINP.n113 4.5005
R49428 VINP.n262 VINP.n113 4.5005
R49429 VINP.n308 VINP.n113 4.5005
R49430 VINP.n261 VINP.n113 4.5005
R49431 VINP.n310 VINP.n113 4.5005
R49432 VINP.n260 VINP.n113 4.5005
R49433 VINP.n312 VINP.n113 4.5005
R49434 VINP.n259 VINP.n113 4.5005
R49435 VINP.n314 VINP.n113 4.5005
R49436 VINP.n258 VINP.n113 4.5005
R49437 VINP.n316 VINP.n113 4.5005
R49438 VINP.n257 VINP.n113 4.5005
R49439 VINP.n318 VINP.n113 4.5005
R49440 VINP.n256 VINP.n113 4.5005
R49441 VINP.n320 VINP.n113 4.5005
R49442 VINP.n255 VINP.n113 4.5005
R49443 VINP.n322 VINP.n113 4.5005
R49444 VINP.n254 VINP.n113 4.5005
R49445 VINP.n324 VINP.n113 4.5005
R49446 VINP.n253 VINP.n113 4.5005
R49447 VINP.n326 VINP.n113 4.5005
R49448 VINP.n252 VINP.n113 4.5005
R49449 VINP.n328 VINP.n113 4.5005
R49450 VINP.n251 VINP.n113 4.5005
R49451 VINP.n330 VINP.n113 4.5005
R49452 VINP.n250 VINP.n113 4.5005
R49453 VINP.n332 VINP.n113 4.5005
R49454 VINP.n249 VINP.n113 4.5005
R49455 VINP.n334 VINP.n113 4.5005
R49456 VINP.n248 VINP.n113 4.5005
R49457 VINP.n336 VINP.n113 4.5005
R49458 VINP.n247 VINP.n113 4.5005
R49459 VINP.n338 VINP.n113 4.5005
R49460 VINP.n246 VINP.n113 4.5005
R49461 VINP.n340 VINP.n113 4.5005
R49462 VINP.n245 VINP.n113 4.5005
R49463 VINP.n342 VINP.n113 4.5005
R49464 VINP.n244 VINP.n113 4.5005
R49465 VINP.n344 VINP.n113 4.5005
R49466 VINP.n243 VINP.n113 4.5005
R49467 VINP.n346 VINP.n113 4.5005
R49468 VINP.n242 VINP.n113 4.5005
R49469 VINP.n348 VINP.n113 4.5005
R49470 VINP.n241 VINP.n113 4.5005
R49471 VINP.n350 VINP.n113 4.5005
R49472 VINP.n240 VINP.n113 4.5005
R49473 VINP.n352 VINP.n113 4.5005
R49474 VINP.n239 VINP.n113 4.5005
R49475 VINP.n354 VINP.n113 4.5005
R49476 VINP.n238 VINP.n113 4.5005
R49477 VINP.n356 VINP.n113 4.5005
R49478 VINP.n237 VINP.n113 4.5005
R49479 VINP.n358 VINP.n113 4.5005
R49480 VINP.n236 VINP.n113 4.5005
R49481 VINP.n360 VINP.n113 4.5005
R49482 VINP.n235 VINP.n113 4.5005
R49483 VINP.n362 VINP.n113 4.5005
R49484 VINP.n234 VINP.n113 4.5005
R49485 VINP.n364 VINP.n113 4.5005
R49486 VINP.n233 VINP.n113 4.5005
R49487 VINP.n366 VINP.n113 4.5005
R49488 VINP.n232 VINP.n113 4.5005
R49489 VINP.n368 VINP.n113 4.5005
R49490 VINP.n231 VINP.n113 4.5005
R49491 VINP.n370 VINP.n113 4.5005
R49492 VINP.n230 VINP.n113 4.5005
R49493 VINP.n372 VINP.n113 4.5005
R49494 VINP.n229 VINP.n113 4.5005
R49495 VINP.n374 VINP.n113 4.5005
R49496 VINP.n228 VINP.n113 4.5005
R49497 VINP.n376 VINP.n113 4.5005
R49498 VINP.n227 VINP.n113 4.5005
R49499 VINP.n378 VINP.n113 4.5005
R49500 VINP.n226 VINP.n113 4.5005
R49501 VINP.n380 VINP.n113 4.5005
R49502 VINP.n225 VINP.n113 4.5005
R49503 VINP.n382 VINP.n113 4.5005
R49504 VINP.n224 VINP.n113 4.5005
R49505 VINP.n384 VINP.n113 4.5005
R49506 VINP.n223 VINP.n113 4.5005
R49507 VINP.n386 VINP.n113 4.5005
R49508 VINP.n222 VINP.n113 4.5005
R49509 VINP.n388 VINP.n113 4.5005
R49510 VINP.n221 VINP.n113 4.5005
R49511 VINP.n390 VINP.n113 4.5005
R49512 VINP.n220 VINP.n113 4.5005
R49513 VINP.n392 VINP.n113 4.5005
R49514 VINP.n219 VINP.n113 4.5005
R49515 VINP.n394 VINP.n113 4.5005
R49516 VINP.n218 VINP.n113 4.5005
R49517 VINP.n396 VINP.n113 4.5005
R49518 VINP.n217 VINP.n113 4.5005
R49519 VINP.n398 VINP.n113 4.5005
R49520 VINP.n216 VINP.n113 4.5005
R49521 VINP.n400 VINP.n113 4.5005
R49522 VINP.n215 VINP.n113 4.5005
R49523 VINP.n654 VINP.n113 4.5005
R49524 VINP.n656 VINP.n113 4.5005
R49525 VINP.n113 VINP.n0 4.5005
R49526 VINP.n278 VINP.n188 4.5005
R49527 VINP.n276 VINP.n188 4.5005
R49528 VINP.n280 VINP.n188 4.5005
R49529 VINP.n275 VINP.n188 4.5005
R49530 VINP.n282 VINP.n188 4.5005
R49531 VINP.n274 VINP.n188 4.5005
R49532 VINP.n284 VINP.n188 4.5005
R49533 VINP.n273 VINP.n188 4.5005
R49534 VINP.n286 VINP.n188 4.5005
R49535 VINP.n272 VINP.n188 4.5005
R49536 VINP.n288 VINP.n188 4.5005
R49537 VINP.n271 VINP.n188 4.5005
R49538 VINP.n290 VINP.n188 4.5005
R49539 VINP.n270 VINP.n188 4.5005
R49540 VINP.n292 VINP.n188 4.5005
R49541 VINP.n269 VINP.n188 4.5005
R49542 VINP.n294 VINP.n188 4.5005
R49543 VINP.n268 VINP.n188 4.5005
R49544 VINP.n296 VINP.n188 4.5005
R49545 VINP.n267 VINP.n188 4.5005
R49546 VINP.n298 VINP.n188 4.5005
R49547 VINP.n266 VINP.n188 4.5005
R49548 VINP.n300 VINP.n188 4.5005
R49549 VINP.n265 VINP.n188 4.5005
R49550 VINP.n302 VINP.n188 4.5005
R49551 VINP.n264 VINP.n188 4.5005
R49552 VINP.n304 VINP.n188 4.5005
R49553 VINP.n263 VINP.n188 4.5005
R49554 VINP.n306 VINP.n188 4.5005
R49555 VINP.n262 VINP.n188 4.5005
R49556 VINP.n308 VINP.n188 4.5005
R49557 VINP.n261 VINP.n188 4.5005
R49558 VINP.n310 VINP.n188 4.5005
R49559 VINP.n260 VINP.n188 4.5005
R49560 VINP.n312 VINP.n188 4.5005
R49561 VINP.n259 VINP.n188 4.5005
R49562 VINP.n314 VINP.n188 4.5005
R49563 VINP.n258 VINP.n188 4.5005
R49564 VINP.n316 VINP.n188 4.5005
R49565 VINP.n257 VINP.n188 4.5005
R49566 VINP.n318 VINP.n188 4.5005
R49567 VINP.n256 VINP.n188 4.5005
R49568 VINP.n320 VINP.n188 4.5005
R49569 VINP.n255 VINP.n188 4.5005
R49570 VINP.n322 VINP.n188 4.5005
R49571 VINP.n254 VINP.n188 4.5005
R49572 VINP.n324 VINP.n188 4.5005
R49573 VINP.n253 VINP.n188 4.5005
R49574 VINP.n326 VINP.n188 4.5005
R49575 VINP.n252 VINP.n188 4.5005
R49576 VINP.n328 VINP.n188 4.5005
R49577 VINP.n251 VINP.n188 4.5005
R49578 VINP.n330 VINP.n188 4.5005
R49579 VINP.n250 VINP.n188 4.5005
R49580 VINP.n332 VINP.n188 4.5005
R49581 VINP.n249 VINP.n188 4.5005
R49582 VINP.n334 VINP.n188 4.5005
R49583 VINP.n248 VINP.n188 4.5005
R49584 VINP.n336 VINP.n188 4.5005
R49585 VINP.n247 VINP.n188 4.5005
R49586 VINP.n338 VINP.n188 4.5005
R49587 VINP.n246 VINP.n188 4.5005
R49588 VINP.n340 VINP.n188 4.5005
R49589 VINP.n245 VINP.n188 4.5005
R49590 VINP.n342 VINP.n188 4.5005
R49591 VINP.n244 VINP.n188 4.5005
R49592 VINP.n344 VINP.n188 4.5005
R49593 VINP.n243 VINP.n188 4.5005
R49594 VINP.n346 VINP.n188 4.5005
R49595 VINP.n242 VINP.n188 4.5005
R49596 VINP.n348 VINP.n188 4.5005
R49597 VINP.n241 VINP.n188 4.5005
R49598 VINP.n350 VINP.n188 4.5005
R49599 VINP.n240 VINP.n188 4.5005
R49600 VINP.n352 VINP.n188 4.5005
R49601 VINP.n239 VINP.n188 4.5005
R49602 VINP.n354 VINP.n188 4.5005
R49603 VINP.n238 VINP.n188 4.5005
R49604 VINP.n356 VINP.n188 4.5005
R49605 VINP.n237 VINP.n188 4.5005
R49606 VINP.n358 VINP.n188 4.5005
R49607 VINP.n236 VINP.n188 4.5005
R49608 VINP.n360 VINP.n188 4.5005
R49609 VINP.n235 VINP.n188 4.5005
R49610 VINP.n362 VINP.n188 4.5005
R49611 VINP.n234 VINP.n188 4.5005
R49612 VINP.n364 VINP.n188 4.5005
R49613 VINP.n233 VINP.n188 4.5005
R49614 VINP.n366 VINP.n188 4.5005
R49615 VINP.n232 VINP.n188 4.5005
R49616 VINP.n368 VINP.n188 4.5005
R49617 VINP.n231 VINP.n188 4.5005
R49618 VINP.n370 VINP.n188 4.5005
R49619 VINP.n230 VINP.n188 4.5005
R49620 VINP.n372 VINP.n188 4.5005
R49621 VINP.n229 VINP.n188 4.5005
R49622 VINP.n374 VINP.n188 4.5005
R49623 VINP.n228 VINP.n188 4.5005
R49624 VINP.n376 VINP.n188 4.5005
R49625 VINP.n227 VINP.n188 4.5005
R49626 VINP.n378 VINP.n188 4.5005
R49627 VINP.n226 VINP.n188 4.5005
R49628 VINP.n380 VINP.n188 4.5005
R49629 VINP.n225 VINP.n188 4.5005
R49630 VINP.n382 VINP.n188 4.5005
R49631 VINP.n224 VINP.n188 4.5005
R49632 VINP.n384 VINP.n188 4.5005
R49633 VINP.n223 VINP.n188 4.5005
R49634 VINP.n386 VINP.n188 4.5005
R49635 VINP.n222 VINP.n188 4.5005
R49636 VINP.n388 VINP.n188 4.5005
R49637 VINP.n221 VINP.n188 4.5005
R49638 VINP.n390 VINP.n188 4.5005
R49639 VINP.n220 VINP.n188 4.5005
R49640 VINP.n392 VINP.n188 4.5005
R49641 VINP.n219 VINP.n188 4.5005
R49642 VINP.n394 VINP.n188 4.5005
R49643 VINP.n218 VINP.n188 4.5005
R49644 VINP.n396 VINP.n188 4.5005
R49645 VINP.n217 VINP.n188 4.5005
R49646 VINP.n398 VINP.n188 4.5005
R49647 VINP.n216 VINP.n188 4.5005
R49648 VINP.n400 VINP.n188 4.5005
R49649 VINP.n215 VINP.n188 4.5005
R49650 VINP.n654 VINP.n188 4.5005
R49651 VINP.n656 VINP.n188 4.5005
R49652 VINP.n188 VINP.n0 4.5005
R49653 VINP.n278 VINP.n112 4.5005
R49654 VINP.n276 VINP.n112 4.5005
R49655 VINP.n280 VINP.n112 4.5005
R49656 VINP.n275 VINP.n112 4.5005
R49657 VINP.n282 VINP.n112 4.5005
R49658 VINP.n274 VINP.n112 4.5005
R49659 VINP.n284 VINP.n112 4.5005
R49660 VINP.n273 VINP.n112 4.5005
R49661 VINP.n286 VINP.n112 4.5005
R49662 VINP.n272 VINP.n112 4.5005
R49663 VINP.n288 VINP.n112 4.5005
R49664 VINP.n271 VINP.n112 4.5005
R49665 VINP.n290 VINP.n112 4.5005
R49666 VINP.n270 VINP.n112 4.5005
R49667 VINP.n292 VINP.n112 4.5005
R49668 VINP.n269 VINP.n112 4.5005
R49669 VINP.n294 VINP.n112 4.5005
R49670 VINP.n268 VINP.n112 4.5005
R49671 VINP.n296 VINP.n112 4.5005
R49672 VINP.n267 VINP.n112 4.5005
R49673 VINP.n298 VINP.n112 4.5005
R49674 VINP.n266 VINP.n112 4.5005
R49675 VINP.n300 VINP.n112 4.5005
R49676 VINP.n265 VINP.n112 4.5005
R49677 VINP.n302 VINP.n112 4.5005
R49678 VINP.n264 VINP.n112 4.5005
R49679 VINP.n304 VINP.n112 4.5005
R49680 VINP.n263 VINP.n112 4.5005
R49681 VINP.n306 VINP.n112 4.5005
R49682 VINP.n262 VINP.n112 4.5005
R49683 VINP.n308 VINP.n112 4.5005
R49684 VINP.n261 VINP.n112 4.5005
R49685 VINP.n310 VINP.n112 4.5005
R49686 VINP.n260 VINP.n112 4.5005
R49687 VINP.n312 VINP.n112 4.5005
R49688 VINP.n259 VINP.n112 4.5005
R49689 VINP.n314 VINP.n112 4.5005
R49690 VINP.n258 VINP.n112 4.5005
R49691 VINP.n316 VINP.n112 4.5005
R49692 VINP.n257 VINP.n112 4.5005
R49693 VINP.n318 VINP.n112 4.5005
R49694 VINP.n256 VINP.n112 4.5005
R49695 VINP.n320 VINP.n112 4.5005
R49696 VINP.n255 VINP.n112 4.5005
R49697 VINP.n322 VINP.n112 4.5005
R49698 VINP.n254 VINP.n112 4.5005
R49699 VINP.n324 VINP.n112 4.5005
R49700 VINP.n253 VINP.n112 4.5005
R49701 VINP.n326 VINP.n112 4.5005
R49702 VINP.n252 VINP.n112 4.5005
R49703 VINP.n328 VINP.n112 4.5005
R49704 VINP.n251 VINP.n112 4.5005
R49705 VINP.n330 VINP.n112 4.5005
R49706 VINP.n250 VINP.n112 4.5005
R49707 VINP.n332 VINP.n112 4.5005
R49708 VINP.n249 VINP.n112 4.5005
R49709 VINP.n334 VINP.n112 4.5005
R49710 VINP.n248 VINP.n112 4.5005
R49711 VINP.n336 VINP.n112 4.5005
R49712 VINP.n247 VINP.n112 4.5005
R49713 VINP.n338 VINP.n112 4.5005
R49714 VINP.n246 VINP.n112 4.5005
R49715 VINP.n340 VINP.n112 4.5005
R49716 VINP.n245 VINP.n112 4.5005
R49717 VINP.n342 VINP.n112 4.5005
R49718 VINP.n244 VINP.n112 4.5005
R49719 VINP.n344 VINP.n112 4.5005
R49720 VINP.n243 VINP.n112 4.5005
R49721 VINP.n346 VINP.n112 4.5005
R49722 VINP.n242 VINP.n112 4.5005
R49723 VINP.n348 VINP.n112 4.5005
R49724 VINP.n241 VINP.n112 4.5005
R49725 VINP.n350 VINP.n112 4.5005
R49726 VINP.n240 VINP.n112 4.5005
R49727 VINP.n352 VINP.n112 4.5005
R49728 VINP.n239 VINP.n112 4.5005
R49729 VINP.n354 VINP.n112 4.5005
R49730 VINP.n238 VINP.n112 4.5005
R49731 VINP.n356 VINP.n112 4.5005
R49732 VINP.n237 VINP.n112 4.5005
R49733 VINP.n358 VINP.n112 4.5005
R49734 VINP.n236 VINP.n112 4.5005
R49735 VINP.n360 VINP.n112 4.5005
R49736 VINP.n235 VINP.n112 4.5005
R49737 VINP.n362 VINP.n112 4.5005
R49738 VINP.n234 VINP.n112 4.5005
R49739 VINP.n364 VINP.n112 4.5005
R49740 VINP.n233 VINP.n112 4.5005
R49741 VINP.n366 VINP.n112 4.5005
R49742 VINP.n232 VINP.n112 4.5005
R49743 VINP.n368 VINP.n112 4.5005
R49744 VINP.n231 VINP.n112 4.5005
R49745 VINP.n370 VINP.n112 4.5005
R49746 VINP.n230 VINP.n112 4.5005
R49747 VINP.n372 VINP.n112 4.5005
R49748 VINP.n229 VINP.n112 4.5005
R49749 VINP.n374 VINP.n112 4.5005
R49750 VINP.n228 VINP.n112 4.5005
R49751 VINP.n376 VINP.n112 4.5005
R49752 VINP.n227 VINP.n112 4.5005
R49753 VINP.n378 VINP.n112 4.5005
R49754 VINP.n226 VINP.n112 4.5005
R49755 VINP.n380 VINP.n112 4.5005
R49756 VINP.n225 VINP.n112 4.5005
R49757 VINP.n382 VINP.n112 4.5005
R49758 VINP.n224 VINP.n112 4.5005
R49759 VINP.n384 VINP.n112 4.5005
R49760 VINP.n223 VINP.n112 4.5005
R49761 VINP.n386 VINP.n112 4.5005
R49762 VINP.n222 VINP.n112 4.5005
R49763 VINP.n388 VINP.n112 4.5005
R49764 VINP.n221 VINP.n112 4.5005
R49765 VINP.n390 VINP.n112 4.5005
R49766 VINP.n220 VINP.n112 4.5005
R49767 VINP.n392 VINP.n112 4.5005
R49768 VINP.n219 VINP.n112 4.5005
R49769 VINP.n394 VINP.n112 4.5005
R49770 VINP.n218 VINP.n112 4.5005
R49771 VINP.n396 VINP.n112 4.5005
R49772 VINP.n217 VINP.n112 4.5005
R49773 VINP.n398 VINP.n112 4.5005
R49774 VINP.n216 VINP.n112 4.5005
R49775 VINP.n400 VINP.n112 4.5005
R49776 VINP.n215 VINP.n112 4.5005
R49777 VINP.n654 VINP.n112 4.5005
R49778 VINP.n656 VINP.n112 4.5005
R49779 VINP.n112 VINP.n0 4.5005
R49780 VINP.n278 VINP.n189 4.5005
R49781 VINP.n276 VINP.n189 4.5005
R49782 VINP.n280 VINP.n189 4.5005
R49783 VINP.n275 VINP.n189 4.5005
R49784 VINP.n282 VINP.n189 4.5005
R49785 VINP.n274 VINP.n189 4.5005
R49786 VINP.n284 VINP.n189 4.5005
R49787 VINP.n273 VINP.n189 4.5005
R49788 VINP.n286 VINP.n189 4.5005
R49789 VINP.n272 VINP.n189 4.5005
R49790 VINP.n288 VINP.n189 4.5005
R49791 VINP.n271 VINP.n189 4.5005
R49792 VINP.n290 VINP.n189 4.5005
R49793 VINP.n270 VINP.n189 4.5005
R49794 VINP.n292 VINP.n189 4.5005
R49795 VINP.n269 VINP.n189 4.5005
R49796 VINP.n294 VINP.n189 4.5005
R49797 VINP.n268 VINP.n189 4.5005
R49798 VINP.n296 VINP.n189 4.5005
R49799 VINP.n267 VINP.n189 4.5005
R49800 VINP.n298 VINP.n189 4.5005
R49801 VINP.n266 VINP.n189 4.5005
R49802 VINP.n300 VINP.n189 4.5005
R49803 VINP.n265 VINP.n189 4.5005
R49804 VINP.n302 VINP.n189 4.5005
R49805 VINP.n264 VINP.n189 4.5005
R49806 VINP.n304 VINP.n189 4.5005
R49807 VINP.n263 VINP.n189 4.5005
R49808 VINP.n306 VINP.n189 4.5005
R49809 VINP.n262 VINP.n189 4.5005
R49810 VINP.n308 VINP.n189 4.5005
R49811 VINP.n261 VINP.n189 4.5005
R49812 VINP.n310 VINP.n189 4.5005
R49813 VINP.n260 VINP.n189 4.5005
R49814 VINP.n312 VINP.n189 4.5005
R49815 VINP.n259 VINP.n189 4.5005
R49816 VINP.n314 VINP.n189 4.5005
R49817 VINP.n258 VINP.n189 4.5005
R49818 VINP.n316 VINP.n189 4.5005
R49819 VINP.n257 VINP.n189 4.5005
R49820 VINP.n318 VINP.n189 4.5005
R49821 VINP.n256 VINP.n189 4.5005
R49822 VINP.n320 VINP.n189 4.5005
R49823 VINP.n255 VINP.n189 4.5005
R49824 VINP.n322 VINP.n189 4.5005
R49825 VINP.n254 VINP.n189 4.5005
R49826 VINP.n324 VINP.n189 4.5005
R49827 VINP.n253 VINP.n189 4.5005
R49828 VINP.n326 VINP.n189 4.5005
R49829 VINP.n252 VINP.n189 4.5005
R49830 VINP.n328 VINP.n189 4.5005
R49831 VINP.n251 VINP.n189 4.5005
R49832 VINP.n330 VINP.n189 4.5005
R49833 VINP.n250 VINP.n189 4.5005
R49834 VINP.n332 VINP.n189 4.5005
R49835 VINP.n249 VINP.n189 4.5005
R49836 VINP.n334 VINP.n189 4.5005
R49837 VINP.n248 VINP.n189 4.5005
R49838 VINP.n336 VINP.n189 4.5005
R49839 VINP.n247 VINP.n189 4.5005
R49840 VINP.n338 VINP.n189 4.5005
R49841 VINP.n246 VINP.n189 4.5005
R49842 VINP.n340 VINP.n189 4.5005
R49843 VINP.n245 VINP.n189 4.5005
R49844 VINP.n342 VINP.n189 4.5005
R49845 VINP.n244 VINP.n189 4.5005
R49846 VINP.n344 VINP.n189 4.5005
R49847 VINP.n243 VINP.n189 4.5005
R49848 VINP.n346 VINP.n189 4.5005
R49849 VINP.n242 VINP.n189 4.5005
R49850 VINP.n348 VINP.n189 4.5005
R49851 VINP.n241 VINP.n189 4.5005
R49852 VINP.n350 VINP.n189 4.5005
R49853 VINP.n240 VINP.n189 4.5005
R49854 VINP.n352 VINP.n189 4.5005
R49855 VINP.n239 VINP.n189 4.5005
R49856 VINP.n354 VINP.n189 4.5005
R49857 VINP.n238 VINP.n189 4.5005
R49858 VINP.n356 VINP.n189 4.5005
R49859 VINP.n237 VINP.n189 4.5005
R49860 VINP.n358 VINP.n189 4.5005
R49861 VINP.n236 VINP.n189 4.5005
R49862 VINP.n360 VINP.n189 4.5005
R49863 VINP.n235 VINP.n189 4.5005
R49864 VINP.n362 VINP.n189 4.5005
R49865 VINP.n234 VINP.n189 4.5005
R49866 VINP.n364 VINP.n189 4.5005
R49867 VINP.n233 VINP.n189 4.5005
R49868 VINP.n366 VINP.n189 4.5005
R49869 VINP.n232 VINP.n189 4.5005
R49870 VINP.n368 VINP.n189 4.5005
R49871 VINP.n231 VINP.n189 4.5005
R49872 VINP.n370 VINP.n189 4.5005
R49873 VINP.n230 VINP.n189 4.5005
R49874 VINP.n372 VINP.n189 4.5005
R49875 VINP.n229 VINP.n189 4.5005
R49876 VINP.n374 VINP.n189 4.5005
R49877 VINP.n228 VINP.n189 4.5005
R49878 VINP.n376 VINP.n189 4.5005
R49879 VINP.n227 VINP.n189 4.5005
R49880 VINP.n378 VINP.n189 4.5005
R49881 VINP.n226 VINP.n189 4.5005
R49882 VINP.n380 VINP.n189 4.5005
R49883 VINP.n225 VINP.n189 4.5005
R49884 VINP.n382 VINP.n189 4.5005
R49885 VINP.n224 VINP.n189 4.5005
R49886 VINP.n384 VINP.n189 4.5005
R49887 VINP.n223 VINP.n189 4.5005
R49888 VINP.n386 VINP.n189 4.5005
R49889 VINP.n222 VINP.n189 4.5005
R49890 VINP.n388 VINP.n189 4.5005
R49891 VINP.n221 VINP.n189 4.5005
R49892 VINP.n390 VINP.n189 4.5005
R49893 VINP.n220 VINP.n189 4.5005
R49894 VINP.n392 VINP.n189 4.5005
R49895 VINP.n219 VINP.n189 4.5005
R49896 VINP.n394 VINP.n189 4.5005
R49897 VINP.n218 VINP.n189 4.5005
R49898 VINP.n396 VINP.n189 4.5005
R49899 VINP.n217 VINP.n189 4.5005
R49900 VINP.n398 VINP.n189 4.5005
R49901 VINP.n216 VINP.n189 4.5005
R49902 VINP.n400 VINP.n189 4.5005
R49903 VINP.n215 VINP.n189 4.5005
R49904 VINP.n654 VINP.n189 4.5005
R49905 VINP.n656 VINP.n189 4.5005
R49906 VINP.n189 VINP.n0 4.5005
R49907 VINP.n278 VINP.n111 4.5005
R49908 VINP.n276 VINP.n111 4.5005
R49909 VINP.n280 VINP.n111 4.5005
R49910 VINP.n275 VINP.n111 4.5005
R49911 VINP.n282 VINP.n111 4.5005
R49912 VINP.n274 VINP.n111 4.5005
R49913 VINP.n284 VINP.n111 4.5005
R49914 VINP.n273 VINP.n111 4.5005
R49915 VINP.n286 VINP.n111 4.5005
R49916 VINP.n272 VINP.n111 4.5005
R49917 VINP.n288 VINP.n111 4.5005
R49918 VINP.n271 VINP.n111 4.5005
R49919 VINP.n290 VINP.n111 4.5005
R49920 VINP.n270 VINP.n111 4.5005
R49921 VINP.n292 VINP.n111 4.5005
R49922 VINP.n269 VINP.n111 4.5005
R49923 VINP.n294 VINP.n111 4.5005
R49924 VINP.n268 VINP.n111 4.5005
R49925 VINP.n296 VINP.n111 4.5005
R49926 VINP.n267 VINP.n111 4.5005
R49927 VINP.n298 VINP.n111 4.5005
R49928 VINP.n266 VINP.n111 4.5005
R49929 VINP.n300 VINP.n111 4.5005
R49930 VINP.n265 VINP.n111 4.5005
R49931 VINP.n302 VINP.n111 4.5005
R49932 VINP.n264 VINP.n111 4.5005
R49933 VINP.n304 VINP.n111 4.5005
R49934 VINP.n263 VINP.n111 4.5005
R49935 VINP.n306 VINP.n111 4.5005
R49936 VINP.n262 VINP.n111 4.5005
R49937 VINP.n308 VINP.n111 4.5005
R49938 VINP.n261 VINP.n111 4.5005
R49939 VINP.n310 VINP.n111 4.5005
R49940 VINP.n260 VINP.n111 4.5005
R49941 VINP.n312 VINP.n111 4.5005
R49942 VINP.n259 VINP.n111 4.5005
R49943 VINP.n314 VINP.n111 4.5005
R49944 VINP.n258 VINP.n111 4.5005
R49945 VINP.n316 VINP.n111 4.5005
R49946 VINP.n257 VINP.n111 4.5005
R49947 VINP.n318 VINP.n111 4.5005
R49948 VINP.n256 VINP.n111 4.5005
R49949 VINP.n320 VINP.n111 4.5005
R49950 VINP.n255 VINP.n111 4.5005
R49951 VINP.n322 VINP.n111 4.5005
R49952 VINP.n254 VINP.n111 4.5005
R49953 VINP.n324 VINP.n111 4.5005
R49954 VINP.n253 VINP.n111 4.5005
R49955 VINP.n326 VINP.n111 4.5005
R49956 VINP.n252 VINP.n111 4.5005
R49957 VINP.n328 VINP.n111 4.5005
R49958 VINP.n251 VINP.n111 4.5005
R49959 VINP.n330 VINP.n111 4.5005
R49960 VINP.n250 VINP.n111 4.5005
R49961 VINP.n332 VINP.n111 4.5005
R49962 VINP.n249 VINP.n111 4.5005
R49963 VINP.n334 VINP.n111 4.5005
R49964 VINP.n248 VINP.n111 4.5005
R49965 VINP.n336 VINP.n111 4.5005
R49966 VINP.n247 VINP.n111 4.5005
R49967 VINP.n338 VINP.n111 4.5005
R49968 VINP.n246 VINP.n111 4.5005
R49969 VINP.n340 VINP.n111 4.5005
R49970 VINP.n245 VINP.n111 4.5005
R49971 VINP.n342 VINP.n111 4.5005
R49972 VINP.n244 VINP.n111 4.5005
R49973 VINP.n344 VINP.n111 4.5005
R49974 VINP.n243 VINP.n111 4.5005
R49975 VINP.n346 VINP.n111 4.5005
R49976 VINP.n242 VINP.n111 4.5005
R49977 VINP.n348 VINP.n111 4.5005
R49978 VINP.n241 VINP.n111 4.5005
R49979 VINP.n350 VINP.n111 4.5005
R49980 VINP.n240 VINP.n111 4.5005
R49981 VINP.n352 VINP.n111 4.5005
R49982 VINP.n239 VINP.n111 4.5005
R49983 VINP.n354 VINP.n111 4.5005
R49984 VINP.n238 VINP.n111 4.5005
R49985 VINP.n356 VINP.n111 4.5005
R49986 VINP.n237 VINP.n111 4.5005
R49987 VINP.n358 VINP.n111 4.5005
R49988 VINP.n236 VINP.n111 4.5005
R49989 VINP.n360 VINP.n111 4.5005
R49990 VINP.n235 VINP.n111 4.5005
R49991 VINP.n362 VINP.n111 4.5005
R49992 VINP.n234 VINP.n111 4.5005
R49993 VINP.n364 VINP.n111 4.5005
R49994 VINP.n233 VINP.n111 4.5005
R49995 VINP.n366 VINP.n111 4.5005
R49996 VINP.n232 VINP.n111 4.5005
R49997 VINP.n368 VINP.n111 4.5005
R49998 VINP.n231 VINP.n111 4.5005
R49999 VINP.n370 VINP.n111 4.5005
R50000 VINP.n230 VINP.n111 4.5005
R50001 VINP.n372 VINP.n111 4.5005
R50002 VINP.n229 VINP.n111 4.5005
R50003 VINP.n374 VINP.n111 4.5005
R50004 VINP.n228 VINP.n111 4.5005
R50005 VINP.n376 VINP.n111 4.5005
R50006 VINP.n227 VINP.n111 4.5005
R50007 VINP.n378 VINP.n111 4.5005
R50008 VINP.n226 VINP.n111 4.5005
R50009 VINP.n380 VINP.n111 4.5005
R50010 VINP.n225 VINP.n111 4.5005
R50011 VINP.n382 VINP.n111 4.5005
R50012 VINP.n224 VINP.n111 4.5005
R50013 VINP.n384 VINP.n111 4.5005
R50014 VINP.n223 VINP.n111 4.5005
R50015 VINP.n386 VINP.n111 4.5005
R50016 VINP.n222 VINP.n111 4.5005
R50017 VINP.n388 VINP.n111 4.5005
R50018 VINP.n221 VINP.n111 4.5005
R50019 VINP.n390 VINP.n111 4.5005
R50020 VINP.n220 VINP.n111 4.5005
R50021 VINP.n392 VINP.n111 4.5005
R50022 VINP.n219 VINP.n111 4.5005
R50023 VINP.n394 VINP.n111 4.5005
R50024 VINP.n218 VINP.n111 4.5005
R50025 VINP.n396 VINP.n111 4.5005
R50026 VINP.n217 VINP.n111 4.5005
R50027 VINP.n398 VINP.n111 4.5005
R50028 VINP.n216 VINP.n111 4.5005
R50029 VINP.n400 VINP.n111 4.5005
R50030 VINP.n215 VINP.n111 4.5005
R50031 VINP.n654 VINP.n111 4.5005
R50032 VINP.n656 VINP.n111 4.5005
R50033 VINP.n111 VINP.n0 4.5005
R50034 VINP.n278 VINP.n190 4.5005
R50035 VINP.n276 VINP.n190 4.5005
R50036 VINP.n280 VINP.n190 4.5005
R50037 VINP.n275 VINP.n190 4.5005
R50038 VINP.n282 VINP.n190 4.5005
R50039 VINP.n274 VINP.n190 4.5005
R50040 VINP.n284 VINP.n190 4.5005
R50041 VINP.n273 VINP.n190 4.5005
R50042 VINP.n286 VINP.n190 4.5005
R50043 VINP.n272 VINP.n190 4.5005
R50044 VINP.n288 VINP.n190 4.5005
R50045 VINP.n271 VINP.n190 4.5005
R50046 VINP.n290 VINP.n190 4.5005
R50047 VINP.n270 VINP.n190 4.5005
R50048 VINP.n292 VINP.n190 4.5005
R50049 VINP.n269 VINP.n190 4.5005
R50050 VINP.n294 VINP.n190 4.5005
R50051 VINP.n268 VINP.n190 4.5005
R50052 VINP.n296 VINP.n190 4.5005
R50053 VINP.n267 VINP.n190 4.5005
R50054 VINP.n298 VINP.n190 4.5005
R50055 VINP.n266 VINP.n190 4.5005
R50056 VINP.n300 VINP.n190 4.5005
R50057 VINP.n265 VINP.n190 4.5005
R50058 VINP.n302 VINP.n190 4.5005
R50059 VINP.n264 VINP.n190 4.5005
R50060 VINP.n304 VINP.n190 4.5005
R50061 VINP.n263 VINP.n190 4.5005
R50062 VINP.n306 VINP.n190 4.5005
R50063 VINP.n262 VINP.n190 4.5005
R50064 VINP.n308 VINP.n190 4.5005
R50065 VINP.n261 VINP.n190 4.5005
R50066 VINP.n310 VINP.n190 4.5005
R50067 VINP.n260 VINP.n190 4.5005
R50068 VINP.n312 VINP.n190 4.5005
R50069 VINP.n259 VINP.n190 4.5005
R50070 VINP.n314 VINP.n190 4.5005
R50071 VINP.n258 VINP.n190 4.5005
R50072 VINP.n316 VINP.n190 4.5005
R50073 VINP.n257 VINP.n190 4.5005
R50074 VINP.n318 VINP.n190 4.5005
R50075 VINP.n256 VINP.n190 4.5005
R50076 VINP.n320 VINP.n190 4.5005
R50077 VINP.n255 VINP.n190 4.5005
R50078 VINP.n322 VINP.n190 4.5005
R50079 VINP.n254 VINP.n190 4.5005
R50080 VINP.n324 VINP.n190 4.5005
R50081 VINP.n253 VINP.n190 4.5005
R50082 VINP.n326 VINP.n190 4.5005
R50083 VINP.n252 VINP.n190 4.5005
R50084 VINP.n328 VINP.n190 4.5005
R50085 VINP.n251 VINP.n190 4.5005
R50086 VINP.n330 VINP.n190 4.5005
R50087 VINP.n250 VINP.n190 4.5005
R50088 VINP.n332 VINP.n190 4.5005
R50089 VINP.n249 VINP.n190 4.5005
R50090 VINP.n334 VINP.n190 4.5005
R50091 VINP.n248 VINP.n190 4.5005
R50092 VINP.n336 VINP.n190 4.5005
R50093 VINP.n247 VINP.n190 4.5005
R50094 VINP.n338 VINP.n190 4.5005
R50095 VINP.n246 VINP.n190 4.5005
R50096 VINP.n340 VINP.n190 4.5005
R50097 VINP.n245 VINP.n190 4.5005
R50098 VINP.n342 VINP.n190 4.5005
R50099 VINP.n244 VINP.n190 4.5005
R50100 VINP.n344 VINP.n190 4.5005
R50101 VINP.n243 VINP.n190 4.5005
R50102 VINP.n346 VINP.n190 4.5005
R50103 VINP.n242 VINP.n190 4.5005
R50104 VINP.n348 VINP.n190 4.5005
R50105 VINP.n241 VINP.n190 4.5005
R50106 VINP.n350 VINP.n190 4.5005
R50107 VINP.n240 VINP.n190 4.5005
R50108 VINP.n352 VINP.n190 4.5005
R50109 VINP.n239 VINP.n190 4.5005
R50110 VINP.n354 VINP.n190 4.5005
R50111 VINP.n238 VINP.n190 4.5005
R50112 VINP.n356 VINP.n190 4.5005
R50113 VINP.n237 VINP.n190 4.5005
R50114 VINP.n358 VINP.n190 4.5005
R50115 VINP.n236 VINP.n190 4.5005
R50116 VINP.n360 VINP.n190 4.5005
R50117 VINP.n235 VINP.n190 4.5005
R50118 VINP.n362 VINP.n190 4.5005
R50119 VINP.n234 VINP.n190 4.5005
R50120 VINP.n364 VINP.n190 4.5005
R50121 VINP.n233 VINP.n190 4.5005
R50122 VINP.n366 VINP.n190 4.5005
R50123 VINP.n232 VINP.n190 4.5005
R50124 VINP.n368 VINP.n190 4.5005
R50125 VINP.n231 VINP.n190 4.5005
R50126 VINP.n370 VINP.n190 4.5005
R50127 VINP.n230 VINP.n190 4.5005
R50128 VINP.n372 VINP.n190 4.5005
R50129 VINP.n229 VINP.n190 4.5005
R50130 VINP.n374 VINP.n190 4.5005
R50131 VINP.n228 VINP.n190 4.5005
R50132 VINP.n376 VINP.n190 4.5005
R50133 VINP.n227 VINP.n190 4.5005
R50134 VINP.n378 VINP.n190 4.5005
R50135 VINP.n226 VINP.n190 4.5005
R50136 VINP.n380 VINP.n190 4.5005
R50137 VINP.n225 VINP.n190 4.5005
R50138 VINP.n382 VINP.n190 4.5005
R50139 VINP.n224 VINP.n190 4.5005
R50140 VINP.n384 VINP.n190 4.5005
R50141 VINP.n223 VINP.n190 4.5005
R50142 VINP.n386 VINP.n190 4.5005
R50143 VINP.n222 VINP.n190 4.5005
R50144 VINP.n388 VINP.n190 4.5005
R50145 VINP.n221 VINP.n190 4.5005
R50146 VINP.n390 VINP.n190 4.5005
R50147 VINP.n220 VINP.n190 4.5005
R50148 VINP.n392 VINP.n190 4.5005
R50149 VINP.n219 VINP.n190 4.5005
R50150 VINP.n394 VINP.n190 4.5005
R50151 VINP.n218 VINP.n190 4.5005
R50152 VINP.n396 VINP.n190 4.5005
R50153 VINP.n217 VINP.n190 4.5005
R50154 VINP.n398 VINP.n190 4.5005
R50155 VINP.n216 VINP.n190 4.5005
R50156 VINP.n400 VINP.n190 4.5005
R50157 VINP.n215 VINP.n190 4.5005
R50158 VINP.n654 VINP.n190 4.5005
R50159 VINP.n656 VINP.n190 4.5005
R50160 VINP.n190 VINP.n0 4.5005
R50161 VINP.n278 VINP.n110 4.5005
R50162 VINP.n276 VINP.n110 4.5005
R50163 VINP.n280 VINP.n110 4.5005
R50164 VINP.n275 VINP.n110 4.5005
R50165 VINP.n282 VINP.n110 4.5005
R50166 VINP.n274 VINP.n110 4.5005
R50167 VINP.n284 VINP.n110 4.5005
R50168 VINP.n273 VINP.n110 4.5005
R50169 VINP.n286 VINP.n110 4.5005
R50170 VINP.n272 VINP.n110 4.5005
R50171 VINP.n288 VINP.n110 4.5005
R50172 VINP.n271 VINP.n110 4.5005
R50173 VINP.n290 VINP.n110 4.5005
R50174 VINP.n270 VINP.n110 4.5005
R50175 VINP.n292 VINP.n110 4.5005
R50176 VINP.n269 VINP.n110 4.5005
R50177 VINP.n294 VINP.n110 4.5005
R50178 VINP.n268 VINP.n110 4.5005
R50179 VINP.n296 VINP.n110 4.5005
R50180 VINP.n267 VINP.n110 4.5005
R50181 VINP.n298 VINP.n110 4.5005
R50182 VINP.n266 VINP.n110 4.5005
R50183 VINP.n300 VINP.n110 4.5005
R50184 VINP.n265 VINP.n110 4.5005
R50185 VINP.n302 VINP.n110 4.5005
R50186 VINP.n264 VINP.n110 4.5005
R50187 VINP.n304 VINP.n110 4.5005
R50188 VINP.n263 VINP.n110 4.5005
R50189 VINP.n306 VINP.n110 4.5005
R50190 VINP.n262 VINP.n110 4.5005
R50191 VINP.n308 VINP.n110 4.5005
R50192 VINP.n261 VINP.n110 4.5005
R50193 VINP.n310 VINP.n110 4.5005
R50194 VINP.n260 VINP.n110 4.5005
R50195 VINP.n312 VINP.n110 4.5005
R50196 VINP.n259 VINP.n110 4.5005
R50197 VINP.n314 VINP.n110 4.5005
R50198 VINP.n258 VINP.n110 4.5005
R50199 VINP.n316 VINP.n110 4.5005
R50200 VINP.n257 VINP.n110 4.5005
R50201 VINP.n318 VINP.n110 4.5005
R50202 VINP.n256 VINP.n110 4.5005
R50203 VINP.n320 VINP.n110 4.5005
R50204 VINP.n255 VINP.n110 4.5005
R50205 VINP.n322 VINP.n110 4.5005
R50206 VINP.n254 VINP.n110 4.5005
R50207 VINP.n324 VINP.n110 4.5005
R50208 VINP.n253 VINP.n110 4.5005
R50209 VINP.n326 VINP.n110 4.5005
R50210 VINP.n252 VINP.n110 4.5005
R50211 VINP.n328 VINP.n110 4.5005
R50212 VINP.n251 VINP.n110 4.5005
R50213 VINP.n330 VINP.n110 4.5005
R50214 VINP.n250 VINP.n110 4.5005
R50215 VINP.n332 VINP.n110 4.5005
R50216 VINP.n249 VINP.n110 4.5005
R50217 VINP.n334 VINP.n110 4.5005
R50218 VINP.n248 VINP.n110 4.5005
R50219 VINP.n336 VINP.n110 4.5005
R50220 VINP.n247 VINP.n110 4.5005
R50221 VINP.n338 VINP.n110 4.5005
R50222 VINP.n246 VINP.n110 4.5005
R50223 VINP.n340 VINP.n110 4.5005
R50224 VINP.n245 VINP.n110 4.5005
R50225 VINP.n342 VINP.n110 4.5005
R50226 VINP.n244 VINP.n110 4.5005
R50227 VINP.n344 VINP.n110 4.5005
R50228 VINP.n243 VINP.n110 4.5005
R50229 VINP.n346 VINP.n110 4.5005
R50230 VINP.n242 VINP.n110 4.5005
R50231 VINP.n348 VINP.n110 4.5005
R50232 VINP.n241 VINP.n110 4.5005
R50233 VINP.n350 VINP.n110 4.5005
R50234 VINP.n240 VINP.n110 4.5005
R50235 VINP.n352 VINP.n110 4.5005
R50236 VINP.n239 VINP.n110 4.5005
R50237 VINP.n354 VINP.n110 4.5005
R50238 VINP.n238 VINP.n110 4.5005
R50239 VINP.n356 VINP.n110 4.5005
R50240 VINP.n237 VINP.n110 4.5005
R50241 VINP.n358 VINP.n110 4.5005
R50242 VINP.n236 VINP.n110 4.5005
R50243 VINP.n360 VINP.n110 4.5005
R50244 VINP.n235 VINP.n110 4.5005
R50245 VINP.n362 VINP.n110 4.5005
R50246 VINP.n234 VINP.n110 4.5005
R50247 VINP.n364 VINP.n110 4.5005
R50248 VINP.n233 VINP.n110 4.5005
R50249 VINP.n366 VINP.n110 4.5005
R50250 VINP.n232 VINP.n110 4.5005
R50251 VINP.n368 VINP.n110 4.5005
R50252 VINP.n231 VINP.n110 4.5005
R50253 VINP.n370 VINP.n110 4.5005
R50254 VINP.n230 VINP.n110 4.5005
R50255 VINP.n372 VINP.n110 4.5005
R50256 VINP.n229 VINP.n110 4.5005
R50257 VINP.n374 VINP.n110 4.5005
R50258 VINP.n228 VINP.n110 4.5005
R50259 VINP.n376 VINP.n110 4.5005
R50260 VINP.n227 VINP.n110 4.5005
R50261 VINP.n378 VINP.n110 4.5005
R50262 VINP.n226 VINP.n110 4.5005
R50263 VINP.n380 VINP.n110 4.5005
R50264 VINP.n225 VINP.n110 4.5005
R50265 VINP.n382 VINP.n110 4.5005
R50266 VINP.n224 VINP.n110 4.5005
R50267 VINP.n384 VINP.n110 4.5005
R50268 VINP.n223 VINP.n110 4.5005
R50269 VINP.n386 VINP.n110 4.5005
R50270 VINP.n222 VINP.n110 4.5005
R50271 VINP.n388 VINP.n110 4.5005
R50272 VINP.n221 VINP.n110 4.5005
R50273 VINP.n390 VINP.n110 4.5005
R50274 VINP.n220 VINP.n110 4.5005
R50275 VINP.n392 VINP.n110 4.5005
R50276 VINP.n219 VINP.n110 4.5005
R50277 VINP.n394 VINP.n110 4.5005
R50278 VINP.n218 VINP.n110 4.5005
R50279 VINP.n396 VINP.n110 4.5005
R50280 VINP.n217 VINP.n110 4.5005
R50281 VINP.n398 VINP.n110 4.5005
R50282 VINP.n216 VINP.n110 4.5005
R50283 VINP.n400 VINP.n110 4.5005
R50284 VINP.n215 VINP.n110 4.5005
R50285 VINP.n654 VINP.n110 4.5005
R50286 VINP.n656 VINP.n110 4.5005
R50287 VINP.n110 VINP.n0 4.5005
R50288 VINP.n278 VINP.n191 4.5005
R50289 VINP.n276 VINP.n191 4.5005
R50290 VINP.n280 VINP.n191 4.5005
R50291 VINP.n275 VINP.n191 4.5005
R50292 VINP.n282 VINP.n191 4.5005
R50293 VINP.n274 VINP.n191 4.5005
R50294 VINP.n284 VINP.n191 4.5005
R50295 VINP.n273 VINP.n191 4.5005
R50296 VINP.n286 VINP.n191 4.5005
R50297 VINP.n272 VINP.n191 4.5005
R50298 VINP.n288 VINP.n191 4.5005
R50299 VINP.n271 VINP.n191 4.5005
R50300 VINP.n290 VINP.n191 4.5005
R50301 VINP.n270 VINP.n191 4.5005
R50302 VINP.n292 VINP.n191 4.5005
R50303 VINP.n269 VINP.n191 4.5005
R50304 VINP.n294 VINP.n191 4.5005
R50305 VINP.n268 VINP.n191 4.5005
R50306 VINP.n296 VINP.n191 4.5005
R50307 VINP.n267 VINP.n191 4.5005
R50308 VINP.n298 VINP.n191 4.5005
R50309 VINP.n266 VINP.n191 4.5005
R50310 VINP.n300 VINP.n191 4.5005
R50311 VINP.n265 VINP.n191 4.5005
R50312 VINP.n302 VINP.n191 4.5005
R50313 VINP.n264 VINP.n191 4.5005
R50314 VINP.n304 VINP.n191 4.5005
R50315 VINP.n263 VINP.n191 4.5005
R50316 VINP.n306 VINP.n191 4.5005
R50317 VINP.n262 VINP.n191 4.5005
R50318 VINP.n308 VINP.n191 4.5005
R50319 VINP.n261 VINP.n191 4.5005
R50320 VINP.n310 VINP.n191 4.5005
R50321 VINP.n260 VINP.n191 4.5005
R50322 VINP.n312 VINP.n191 4.5005
R50323 VINP.n259 VINP.n191 4.5005
R50324 VINP.n314 VINP.n191 4.5005
R50325 VINP.n258 VINP.n191 4.5005
R50326 VINP.n316 VINP.n191 4.5005
R50327 VINP.n257 VINP.n191 4.5005
R50328 VINP.n318 VINP.n191 4.5005
R50329 VINP.n256 VINP.n191 4.5005
R50330 VINP.n320 VINP.n191 4.5005
R50331 VINP.n255 VINP.n191 4.5005
R50332 VINP.n322 VINP.n191 4.5005
R50333 VINP.n254 VINP.n191 4.5005
R50334 VINP.n324 VINP.n191 4.5005
R50335 VINP.n253 VINP.n191 4.5005
R50336 VINP.n326 VINP.n191 4.5005
R50337 VINP.n252 VINP.n191 4.5005
R50338 VINP.n328 VINP.n191 4.5005
R50339 VINP.n251 VINP.n191 4.5005
R50340 VINP.n330 VINP.n191 4.5005
R50341 VINP.n250 VINP.n191 4.5005
R50342 VINP.n332 VINP.n191 4.5005
R50343 VINP.n249 VINP.n191 4.5005
R50344 VINP.n334 VINP.n191 4.5005
R50345 VINP.n248 VINP.n191 4.5005
R50346 VINP.n336 VINP.n191 4.5005
R50347 VINP.n247 VINP.n191 4.5005
R50348 VINP.n338 VINP.n191 4.5005
R50349 VINP.n246 VINP.n191 4.5005
R50350 VINP.n340 VINP.n191 4.5005
R50351 VINP.n245 VINP.n191 4.5005
R50352 VINP.n342 VINP.n191 4.5005
R50353 VINP.n244 VINP.n191 4.5005
R50354 VINP.n344 VINP.n191 4.5005
R50355 VINP.n243 VINP.n191 4.5005
R50356 VINP.n346 VINP.n191 4.5005
R50357 VINP.n242 VINP.n191 4.5005
R50358 VINP.n348 VINP.n191 4.5005
R50359 VINP.n241 VINP.n191 4.5005
R50360 VINP.n350 VINP.n191 4.5005
R50361 VINP.n240 VINP.n191 4.5005
R50362 VINP.n352 VINP.n191 4.5005
R50363 VINP.n239 VINP.n191 4.5005
R50364 VINP.n354 VINP.n191 4.5005
R50365 VINP.n238 VINP.n191 4.5005
R50366 VINP.n356 VINP.n191 4.5005
R50367 VINP.n237 VINP.n191 4.5005
R50368 VINP.n358 VINP.n191 4.5005
R50369 VINP.n236 VINP.n191 4.5005
R50370 VINP.n360 VINP.n191 4.5005
R50371 VINP.n235 VINP.n191 4.5005
R50372 VINP.n362 VINP.n191 4.5005
R50373 VINP.n234 VINP.n191 4.5005
R50374 VINP.n364 VINP.n191 4.5005
R50375 VINP.n233 VINP.n191 4.5005
R50376 VINP.n366 VINP.n191 4.5005
R50377 VINP.n232 VINP.n191 4.5005
R50378 VINP.n368 VINP.n191 4.5005
R50379 VINP.n231 VINP.n191 4.5005
R50380 VINP.n370 VINP.n191 4.5005
R50381 VINP.n230 VINP.n191 4.5005
R50382 VINP.n372 VINP.n191 4.5005
R50383 VINP.n229 VINP.n191 4.5005
R50384 VINP.n374 VINP.n191 4.5005
R50385 VINP.n228 VINP.n191 4.5005
R50386 VINP.n376 VINP.n191 4.5005
R50387 VINP.n227 VINP.n191 4.5005
R50388 VINP.n378 VINP.n191 4.5005
R50389 VINP.n226 VINP.n191 4.5005
R50390 VINP.n380 VINP.n191 4.5005
R50391 VINP.n225 VINP.n191 4.5005
R50392 VINP.n382 VINP.n191 4.5005
R50393 VINP.n224 VINP.n191 4.5005
R50394 VINP.n384 VINP.n191 4.5005
R50395 VINP.n223 VINP.n191 4.5005
R50396 VINP.n386 VINP.n191 4.5005
R50397 VINP.n222 VINP.n191 4.5005
R50398 VINP.n388 VINP.n191 4.5005
R50399 VINP.n221 VINP.n191 4.5005
R50400 VINP.n390 VINP.n191 4.5005
R50401 VINP.n220 VINP.n191 4.5005
R50402 VINP.n392 VINP.n191 4.5005
R50403 VINP.n219 VINP.n191 4.5005
R50404 VINP.n394 VINP.n191 4.5005
R50405 VINP.n218 VINP.n191 4.5005
R50406 VINP.n396 VINP.n191 4.5005
R50407 VINP.n217 VINP.n191 4.5005
R50408 VINP.n398 VINP.n191 4.5005
R50409 VINP.n216 VINP.n191 4.5005
R50410 VINP.n400 VINP.n191 4.5005
R50411 VINP.n215 VINP.n191 4.5005
R50412 VINP.n654 VINP.n191 4.5005
R50413 VINP.n656 VINP.n191 4.5005
R50414 VINP.n191 VINP.n0 4.5005
R50415 VINP.n278 VINP.n109 4.5005
R50416 VINP.n276 VINP.n109 4.5005
R50417 VINP.n280 VINP.n109 4.5005
R50418 VINP.n275 VINP.n109 4.5005
R50419 VINP.n282 VINP.n109 4.5005
R50420 VINP.n274 VINP.n109 4.5005
R50421 VINP.n284 VINP.n109 4.5005
R50422 VINP.n273 VINP.n109 4.5005
R50423 VINP.n286 VINP.n109 4.5005
R50424 VINP.n272 VINP.n109 4.5005
R50425 VINP.n288 VINP.n109 4.5005
R50426 VINP.n271 VINP.n109 4.5005
R50427 VINP.n290 VINP.n109 4.5005
R50428 VINP.n270 VINP.n109 4.5005
R50429 VINP.n292 VINP.n109 4.5005
R50430 VINP.n269 VINP.n109 4.5005
R50431 VINP.n294 VINP.n109 4.5005
R50432 VINP.n268 VINP.n109 4.5005
R50433 VINP.n296 VINP.n109 4.5005
R50434 VINP.n267 VINP.n109 4.5005
R50435 VINP.n298 VINP.n109 4.5005
R50436 VINP.n266 VINP.n109 4.5005
R50437 VINP.n300 VINP.n109 4.5005
R50438 VINP.n265 VINP.n109 4.5005
R50439 VINP.n302 VINP.n109 4.5005
R50440 VINP.n264 VINP.n109 4.5005
R50441 VINP.n304 VINP.n109 4.5005
R50442 VINP.n263 VINP.n109 4.5005
R50443 VINP.n306 VINP.n109 4.5005
R50444 VINP.n262 VINP.n109 4.5005
R50445 VINP.n308 VINP.n109 4.5005
R50446 VINP.n261 VINP.n109 4.5005
R50447 VINP.n310 VINP.n109 4.5005
R50448 VINP.n260 VINP.n109 4.5005
R50449 VINP.n312 VINP.n109 4.5005
R50450 VINP.n259 VINP.n109 4.5005
R50451 VINP.n314 VINP.n109 4.5005
R50452 VINP.n258 VINP.n109 4.5005
R50453 VINP.n316 VINP.n109 4.5005
R50454 VINP.n257 VINP.n109 4.5005
R50455 VINP.n318 VINP.n109 4.5005
R50456 VINP.n256 VINP.n109 4.5005
R50457 VINP.n320 VINP.n109 4.5005
R50458 VINP.n255 VINP.n109 4.5005
R50459 VINP.n322 VINP.n109 4.5005
R50460 VINP.n254 VINP.n109 4.5005
R50461 VINP.n324 VINP.n109 4.5005
R50462 VINP.n253 VINP.n109 4.5005
R50463 VINP.n326 VINP.n109 4.5005
R50464 VINP.n252 VINP.n109 4.5005
R50465 VINP.n328 VINP.n109 4.5005
R50466 VINP.n251 VINP.n109 4.5005
R50467 VINP.n330 VINP.n109 4.5005
R50468 VINP.n250 VINP.n109 4.5005
R50469 VINP.n332 VINP.n109 4.5005
R50470 VINP.n249 VINP.n109 4.5005
R50471 VINP.n334 VINP.n109 4.5005
R50472 VINP.n248 VINP.n109 4.5005
R50473 VINP.n336 VINP.n109 4.5005
R50474 VINP.n247 VINP.n109 4.5005
R50475 VINP.n338 VINP.n109 4.5005
R50476 VINP.n246 VINP.n109 4.5005
R50477 VINP.n340 VINP.n109 4.5005
R50478 VINP.n245 VINP.n109 4.5005
R50479 VINP.n342 VINP.n109 4.5005
R50480 VINP.n244 VINP.n109 4.5005
R50481 VINP.n344 VINP.n109 4.5005
R50482 VINP.n243 VINP.n109 4.5005
R50483 VINP.n346 VINP.n109 4.5005
R50484 VINP.n242 VINP.n109 4.5005
R50485 VINP.n348 VINP.n109 4.5005
R50486 VINP.n241 VINP.n109 4.5005
R50487 VINP.n350 VINP.n109 4.5005
R50488 VINP.n240 VINP.n109 4.5005
R50489 VINP.n352 VINP.n109 4.5005
R50490 VINP.n239 VINP.n109 4.5005
R50491 VINP.n354 VINP.n109 4.5005
R50492 VINP.n238 VINP.n109 4.5005
R50493 VINP.n356 VINP.n109 4.5005
R50494 VINP.n237 VINP.n109 4.5005
R50495 VINP.n358 VINP.n109 4.5005
R50496 VINP.n236 VINP.n109 4.5005
R50497 VINP.n360 VINP.n109 4.5005
R50498 VINP.n235 VINP.n109 4.5005
R50499 VINP.n362 VINP.n109 4.5005
R50500 VINP.n234 VINP.n109 4.5005
R50501 VINP.n364 VINP.n109 4.5005
R50502 VINP.n233 VINP.n109 4.5005
R50503 VINP.n366 VINP.n109 4.5005
R50504 VINP.n232 VINP.n109 4.5005
R50505 VINP.n368 VINP.n109 4.5005
R50506 VINP.n231 VINP.n109 4.5005
R50507 VINP.n370 VINP.n109 4.5005
R50508 VINP.n230 VINP.n109 4.5005
R50509 VINP.n372 VINP.n109 4.5005
R50510 VINP.n229 VINP.n109 4.5005
R50511 VINP.n374 VINP.n109 4.5005
R50512 VINP.n228 VINP.n109 4.5005
R50513 VINP.n376 VINP.n109 4.5005
R50514 VINP.n227 VINP.n109 4.5005
R50515 VINP.n378 VINP.n109 4.5005
R50516 VINP.n226 VINP.n109 4.5005
R50517 VINP.n380 VINP.n109 4.5005
R50518 VINP.n225 VINP.n109 4.5005
R50519 VINP.n382 VINP.n109 4.5005
R50520 VINP.n224 VINP.n109 4.5005
R50521 VINP.n384 VINP.n109 4.5005
R50522 VINP.n223 VINP.n109 4.5005
R50523 VINP.n386 VINP.n109 4.5005
R50524 VINP.n222 VINP.n109 4.5005
R50525 VINP.n388 VINP.n109 4.5005
R50526 VINP.n221 VINP.n109 4.5005
R50527 VINP.n390 VINP.n109 4.5005
R50528 VINP.n220 VINP.n109 4.5005
R50529 VINP.n392 VINP.n109 4.5005
R50530 VINP.n219 VINP.n109 4.5005
R50531 VINP.n394 VINP.n109 4.5005
R50532 VINP.n218 VINP.n109 4.5005
R50533 VINP.n396 VINP.n109 4.5005
R50534 VINP.n217 VINP.n109 4.5005
R50535 VINP.n398 VINP.n109 4.5005
R50536 VINP.n216 VINP.n109 4.5005
R50537 VINP.n400 VINP.n109 4.5005
R50538 VINP.n215 VINP.n109 4.5005
R50539 VINP.n654 VINP.n109 4.5005
R50540 VINP.n656 VINP.n109 4.5005
R50541 VINP.n109 VINP.n0 4.5005
R50542 VINP.n278 VINP.n192 4.5005
R50543 VINP.n276 VINP.n192 4.5005
R50544 VINP.n280 VINP.n192 4.5005
R50545 VINP.n275 VINP.n192 4.5005
R50546 VINP.n282 VINP.n192 4.5005
R50547 VINP.n274 VINP.n192 4.5005
R50548 VINP.n284 VINP.n192 4.5005
R50549 VINP.n273 VINP.n192 4.5005
R50550 VINP.n286 VINP.n192 4.5005
R50551 VINP.n272 VINP.n192 4.5005
R50552 VINP.n288 VINP.n192 4.5005
R50553 VINP.n271 VINP.n192 4.5005
R50554 VINP.n290 VINP.n192 4.5005
R50555 VINP.n270 VINP.n192 4.5005
R50556 VINP.n292 VINP.n192 4.5005
R50557 VINP.n269 VINP.n192 4.5005
R50558 VINP.n294 VINP.n192 4.5005
R50559 VINP.n268 VINP.n192 4.5005
R50560 VINP.n296 VINP.n192 4.5005
R50561 VINP.n267 VINP.n192 4.5005
R50562 VINP.n298 VINP.n192 4.5005
R50563 VINP.n266 VINP.n192 4.5005
R50564 VINP.n300 VINP.n192 4.5005
R50565 VINP.n265 VINP.n192 4.5005
R50566 VINP.n302 VINP.n192 4.5005
R50567 VINP.n264 VINP.n192 4.5005
R50568 VINP.n304 VINP.n192 4.5005
R50569 VINP.n263 VINP.n192 4.5005
R50570 VINP.n306 VINP.n192 4.5005
R50571 VINP.n262 VINP.n192 4.5005
R50572 VINP.n308 VINP.n192 4.5005
R50573 VINP.n261 VINP.n192 4.5005
R50574 VINP.n310 VINP.n192 4.5005
R50575 VINP.n260 VINP.n192 4.5005
R50576 VINP.n312 VINP.n192 4.5005
R50577 VINP.n259 VINP.n192 4.5005
R50578 VINP.n314 VINP.n192 4.5005
R50579 VINP.n258 VINP.n192 4.5005
R50580 VINP.n316 VINP.n192 4.5005
R50581 VINP.n257 VINP.n192 4.5005
R50582 VINP.n318 VINP.n192 4.5005
R50583 VINP.n256 VINP.n192 4.5005
R50584 VINP.n320 VINP.n192 4.5005
R50585 VINP.n255 VINP.n192 4.5005
R50586 VINP.n322 VINP.n192 4.5005
R50587 VINP.n254 VINP.n192 4.5005
R50588 VINP.n324 VINP.n192 4.5005
R50589 VINP.n253 VINP.n192 4.5005
R50590 VINP.n326 VINP.n192 4.5005
R50591 VINP.n252 VINP.n192 4.5005
R50592 VINP.n328 VINP.n192 4.5005
R50593 VINP.n251 VINP.n192 4.5005
R50594 VINP.n330 VINP.n192 4.5005
R50595 VINP.n250 VINP.n192 4.5005
R50596 VINP.n332 VINP.n192 4.5005
R50597 VINP.n249 VINP.n192 4.5005
R50598 VINP.n334 VINP.n192 4.5005
R50599 VINP.n248 VINP.n192 4.5005
R50600 VINP.n336 VINP.n192 4.5005
R50601 VINP.n247 VINP.n192 4.5005
R50602 VINP.n338 VINP.n192 4.5005
R50603 VINP.n246 VINP.n192 4.5005
R50604 VINP.n340 VINP.n192 4.5005
R50605 VINP.n245 VINP.n192 4.5005
R50606 VINP.n342 VINP.n192 4.5005
R50607 VINP.n244 VINP.n192 4.5005
R50608 VINP.n344 VINP.n192 4.5005
R50609 VINP.n243 VINP.n192 4.5005
R50610 VINP.n346 VINP.n192 4.5005
R50611 VINP.n242 VINP.n192 4.5005
R50612 VINP.n348 VINP.n192 4.5005
R50613 VINP.n241 VINP.n192 4.5005
R50614 VINP.n350 VINP.n192 4.5005
R50615 VINP.n240 VINP.n192 4.5005
R50616 VINP.n352 VINP.n192 4.5005
R50617 VINP.n239 VINP.n192 4.5005
R50618 VINP.n354 VINP.n192 4.5005
R50619 VINP.n238 VINP.n192 4.5005
R50620 VINP.n356 VINP.n192 4.5005
R50621 VINP.n237 VINP.n192 4.5005
R50622 VINP.n358 VINP.n192 4.5005
R50623 VINP.n236 VINP.n192 4.5005
R50624 VINP.n360 VINP.n192 4.5005
R50625 VINP.n235 VINP.n192 4.5005
R50626 VINP.n362 VINP.n192 4.5005
R50627 VINP.n234 VINP.n192 4.5005
R50628 VINP.n364 VINP.n192 4.5005
R50629 VINP.n233 VINP.n192 4.5005
R50630 VINP.n366 VINP.n192 4.5005
R50631 VINP.n232 VINP.n192 4.5005
R50632 VINP.n368 VINP.n192 4.5005
R50633 VINP.n231 VINP.n192 4.5005
R50634 VINP.n370 VINP.n192 4.5005
R50635 VINP.n230 VINP.n192 4.5005
R50636 VINP.n372 VINP.n192 4.5005
R50637 VINP.n229 VINP.n192 4.5005
R50638 VINP.n374 VINP.n192 4.5005
R50639 VINP.n228 VINP.n192 4.5005
R50640 VINP.n376 VINP.n192 4.5005
R50641 VINP.n227 VINP.n192 4.5005
R50642 VINP.n378 VINP.n192 4.5005
R50643 VINP.n226 VINP.n192 4.5005
R50644 VINP.n380 VINP.n192 4.5005
R50645 VINP.n225 VINP.n192 4.5005
R50646 VINP.n382 VINP.n192 4.5005
R50647 VINP.n224 VINP.n192 4.5005
R50648 VINP.n384 VINP.n192 4.5005
R50649 VINP.n223 VINP.n192 4.5005
R50650 VINP.n386 VINP.n192 4.5005
R50651 VINP.n222 VINP.n192 4.5005
R50652 VINP.n388 VINP.n192 4.5005
R50653 VINP.n221 VINP.n192 4.5005
R50654 VINP.n390 VINP.n192 4.5005
R50655 VINP.n220 VINP.n192 4.5005
R50656 VINP.n392 VINP.n192 4.5005
R50657 VINP.n219 VINP.n192 4.5005
R50658 VINP.n394 VINP.n192 4.5005
R50659 VINP.n218 VINP.n192 4.5005
R50660 VINP.n396 VINP.n192 4.5005
R50661 VINP.n217 VINP.n192 4.5005
R50662 VINP.n398 VINP.n192 4.5005
R50663 VINP.n216 VINP.n192 4.5005
R50664 VINP.n400 VINP.n192 4.5005
R50665 VINP.n215 VINP.n192 4.5005
R50666 VINP.n654 VINP.n192 4.5005
R50667 VINP.n656 VINP.n192 4.5005
R50668 VINP.n192 VINP.n0 4.5005
R50669 VINP.n278 VINP.n108 4.5005
R50670 VINP.n276 VINP.n108 4.5005
R50671 VINP.n280 VINP.n108 4.5005
R50672 VINP.n275 VINP.n108 4.5005
R50673 VINP.n282 VINP.n108 4.5005
R50674 VINP.n274 VINP.n108 4.5005
R50675 VINP.n284 VINP.n108 4.5005
R50676 VINP.n273 VINP.n108 4.5005
R50677 VINP.n286 VINP.n108 4.5005
R50678 VINP.n272 VINP.n108 4.5005
R50679 VINP.n288 VINP.n108 4.5005
R50680 VINP.n271 VINP.n108 4.5005
R50681 VINP.n290 VINP.n108 4.5005
R50682 VINP.n270 VINP.n108 4.5005
R50683 VINP.n292 VINP.n108 4.5005
R50684 VINP.n269 VINP.n108 4.5005
R50685 VINP.n294 VINP.n108 4.5005
R50686 VINP.n268 VINP.n108 4.5005
R50687 VINP.n296 VINP.n108 4.5005
R50688 VINP.n267 VINP.n108 4.5005
R50689 VINP.n298 VINP.n108 4.5005
R50690 VINP.n266 VINP.n108 4.5005
R50691 VINP.n300 VINP.n108 4.5005
R50692 VINP.n265 VINP.n108 4.5005
R50693 VINP.n302 VINP.n108 4.5005
R50694 VINP.n264 VINP.n108 4.5005
R50695 VINP.n304 VINP.n108 4.5005
R50696 VINP.n263 VINP.n108 4.5005
R50697 VINP.n306 VINP.n108 4.5005
R50698 VINP.n262 VINP.n108 4.5005
R50699 VINP.n308 VINP.n108 4.5005
R50700 VINP.n261 VINP.n108 4.5005
R50701 VINP.n310 VINP.n108 4.5005
R50702 VINP.n260 VINP.n108 4.5005
R50703 VINP.n312 VINP.n108 4.5005
R50704 VINP.n259 VINP.n108 4.5005
R50705 VINP.n314 VINP.n108 4.5005
R50706 VINP.n258 VINP.n108 4.5005
R50707 VINP.n316 VINP.n108 4.5005
R50708 VINP.n257 VINP.n108 4.5005
R50709 VINP.n318 VINP.n108 4.5005
R50710 VINP.n256 VINP.n108 4.5005
R50711 VINP.n320 VINP.n108 4.5005
R50712 VINP.n255 VINP.n108 4.5005
R50713 VINP.n322 VINP.n108 4.5005
R50714 VINP.n254 VINP.n108 4.5005
R50715 VINP.n324 VINP.n108 4.5005
R50716 VINP.n253 VINP.n108 4.5005
R50717 VINP.n326 VINP.n108 4.5005
R50718 VINP.n252 VINP.n108 4.5005
R50719 VINP.n328 VINP.n108 4.5005
R50720 VINP.n251 VINP.n108 4.5005
R50721 VINP.n330 VINP.n108 4.5005
R50722 VINP.n250 VINP.n108 4.5005
R50723 VINP.n332 VINP.n108 4.5005
R50724 VINP.n249 VINP.n108 4.5005
R50725 VINP.n334 VINP.n108 4.5005
R50726 VINP.n248 VINP.n108 4.5005
R50727 VINP.n336 VINP.n108 4.5005
R50728 VINP.n247 VINP.n108 4.5005
R50729 VINP.n338 VINP.n108 4.5005
R50730 VINP.n246 VINP.n108 4.5005
R50731 VINP.n340 VINP.n108 4.5005
R50732 VINP.n245 VINP.n108 4.5005
R50733 VINP.n342 VINP.n108 4.5005
R50734 VINP.n244 VINP.n108 4.5005
R50735 VINP.n344 VINP.n108 4.5005
R50736 VINP.n243 VINP.n108 4.5005
R50737 VINP.n346 VINP.n108 4.5005
R50738 VINP.n242 VINP.n108 4.5005
R50739 VINP.n348 VINP.n108 4.5005
R50740 VINP.n241 VINP.n108 4.5005
R50741 VINP.n350 VINP.n108 4.5005
R50742 VINP.n240 VINP.n108 4.5005
R50743 VINP.n352 VINP.n108 4.5005
R50744 VINP.n239 VINP.n108 4.5005
R50745 VINP.n354 VINP.n108 4.5005
R50746 VINP.n238 VINP.n108 4.5005
R50747 VINP.n356 VINP.n108 4.5005
R50748 VINP.n237 VINP.n108 4.5005
R50749 VINP.n358 VINP.n108 4.5005
R50750 VINP.n236 VINP.n108 4.5005
R50751 VINP.n360 VINP.n108 4.5005
R50752 VINP.n235 VINP.n108 4.5005
R50753 VINP.n362 VINP.n108 4.5005
R50754 VINP.n234 VINP.n108 4.5005
R50755 VINP.n364 VINP.n108 4.5005
R50756 VINP.n233 VINP.n108 4.5005
R50757 VINP.n366 VINP.n108 4.5005
R50758 VINP.n232 VINP.n108 4.5005
R50759 VINP.n368 VINP.n108 4.5005
R50760 VINP.n231 VINP.n108 4.5005
R50761 VINP.n370 VINP.n108 4.5005
R50762 VINP.n230 VINP.n108 4.5005
R50763 VINP.n372 VINP.n108 4.5005
R50764 VINP.n229 VINP.n108 4.5005
R50765 VINP.n374 VINP.n108 4.5005
R50766 VINP.n228 VINP.n108 4.5005
R50767 VINP.n376 VINP.n108 4.5005
R50768 VINP.n227 VINP.n108 4.5005
R50769 VINP.n378 VINP.n108 4.5005
R50770 VINP.n226 VINP.n108 4.5005
R50771 VINP.n380 VINP.n108 4.5005
R50772 VINP.n225 VINP.n108 4.5005
R50773 VINP.n382 VINP.n108 4.5005
R50774 VINP.n224 VINP.n108 4.5005
R50775 VINP.n384 VINP.n108 4.5005
R50776 VINP.n223 VINP.n108 4.5005
R50777 VINP.n386 VINP.n108 4.5005
R50778 VINP.n222 VINP.n108 4.5005
R50779 VINP.n388 VINP.n108 4.5005
R50780 VINP.n221 VINP.n108 4.5005
R50781 VINP.n390 VINP.n108 4.5005
R50782 VINP.n220 VINP.n108 4.5005
R50783 VINP.n392 VINP.n108 4.5005
R50784 VINP.n219 VINP.n108 4.5005
R50785 VINP.n394 VINP.n108 4.5005
R50786 VINP.n218 VINP.n108 4.5005
R50787 VINP.n396 VINP.n108 4.5005
R50788 VINP.n217 VINP.n108 4.5005
R50789 VINP.n398 VINP.n108 4.5005
R50790 VINP.n216 VINP.n108 4.5005
R50791 VINP.n400 VINP.n108 4.5005
R50792 VINP.n215 VINP.n108 4.5005
R50793 VINP.n654 VINP.n108 4.5005
R50794 VINP.n656 VINP.n108 4.5005
R50795 VINP.n108 VINP.n0 4.5005
R50796 VINP.n278 VINP.n193 4.5005
R50797 VINP.n276 VINP.n193 4.5005
R50798 VINP.n280 VINP.n193 4.5005
R50799 VINP.n275 VINP.n193 4.5005
R50800 VINP.n282 VINP.n193 4.5005
R50801 VINP.n274 VINP.n193 4.5005
R50802 VINP.n284 VINP.n193 4.5005
R50803 VINP.n273 VINP.n193 4.5005
R50804 VINP.n286 VINP.n193 4.5005
R50805 VINP.n272 VINP.n193 4.5005
R50806 VINP.n288 VINP.n193 4.5005
R50807 VINP.n271 VINP.n193 4.5005
R50808 VINP.n290 VINP.n193 4.5005
R50809 VINP.n270 VINP.n193 4.5005
R50810 VINP.n292 VINP.n193 4.5005
R50811 VINP.n269 VINP.n193 4.5005
R50812 VINP.n294 VINP.n193 4.5005
R50813 VINP.n268 VINP.n193 4.5005
R50814 VINP.n296 VINP.n193 4.5005
R50815 VINP.n267 VINP.n193 4.5005
R50816 VINP.n298 VINP.n193 4.5005
R50817 VINP.n266 VINP.n193 4.5005
R50818 VINP.n300 VINP.n193 4.5005
R50819 VINP.n265 VINP.n193 4.5005
R50820 VINP.n302 VINP.n193 4.5005
R50821 VINP.n264 VINP.n193 4.5005
R50822 VINP.n304 VINP.n193 4.5005
R50823 VINP.n263 VINP.n193 4.5005
R50824 VINP.n306 VINP.n193 4.5005
R50825 VINP.n262 VINP.n193 4.5005
R50826 VINP.n308 VINP.n193 4.5005
R50827 VINP.n261 VINP.n193 4.5005
R50828 VINP.n310 VINP.n193 4.5005
R50829 VINP.n260 VINP.n193 4.5005
R50830 VINP.n312 VINP.n193 4.5005
R50831 VINP.n259 VINP.n193 4.5005
R50832 VINP.n314 VINP.n193 4.5005
R50833 VINP.n258 VINP.n193 4.5005
R50834 VINP.n316 VINP.n193 4.5005
R50835 VINP.n257 VINP.n193 4.5005
R50836 VINP.n318 VINP.n193 4.5005
R50837 VINP.n256 VINP.n193 4.5005
R50838 VINP.n320 VINP.n193 4.5005
R50839 VINP.n255 VINP.n193 4.5005
R50840 VINP.n322 VINP.n193 4.5005
R50841 VINP.n254 VINP.n193 4.5005
R50842 VINP.n324 VINP.n193 4.5005
R50843 VINP.n253 VINP.n193 4.5005
R50844 VINP.n326 VINP.n193 4.5005
R50845 VINP.n252 VINP.n193 4.5005
R50846 VINP.n328 VINP.n193 4.5005
R50847 VINP.n251 VINP.n193 4.5005
R50848 VINP.n330 VINP.n193 4.5005
R50849 VINP.n250 VINP.n193 4.5005
R50850 VINP.n332 VINP.n193 4.5005
R50851 VINP.n249 VINP.n193 4.5005
R50852 VINP.n334 VINP.n193 4.5005
R50853 VINP.n248 VINP.n193 4.5005
R50854 VINP.n336 VINP.n193 4.5005
R50855 VINP.n247 VINP.n193 4.5005
R50856 VINP.n338 VINP.n193 4.5005
R50857 VINP.n246 VINP.n193 4.5005
R50858 VINP.n340 VINP.n193 4.5005
R50859 VINP.n245 VINP.n193 4.5005
R50860 VINP.n342 VINP.n193 4.5005
R50861 VINP.n244 VINP.n193 4.5005
R50862 VINP.n344 VINP.n193 4.5005
R50863 VINP.n243 VINP.n193 4.5005
R50864 VINP.n346 VINP.n193 4.5005
R50865 VINP.n242 VINP.n193 4.5005
R50866 VINP.n348 VINP.n193 4.5005
R50867 VINP.n241 VINP.n193 4.5005
R50868 VINP.n350 VINP.n193 4.5005
R50869 VINP.n240 VINP.n193 4.5005
R50870 VINP.n352 VINP.n193 4.5005
R50871 VINP.n239 VINP.n193 4.5005
R50872 VINP.n354 VINP.n193 4.5005
R50873 VINP.n238 VINP.n193 4.5005
R50874 VINP.n356 VINP.n193 4.5005
R50875 VINP.n237 VINP.n193 4.5005
R50876 VINP.n358 VINP.n193 4.5005
R50877 VINP.n236 VINP.n193 4.5005
R50878 VINP.n360 VINP.n193 4.5005
R50879 VINP.n235 VINP.n193 4.5005
R50880 VINP.n362 VINP.n193 4.5005
R50881 VINP.n234 VINP.n193 4.5005
R50882 VINP.n364 VINP.n193 4.5005
R50883 VINP.n233 VINP.n193 4.5005
R50884 VINP.n366 VINP.n193 4.5005
R50885 VINP.n232 VINP.n193 4.5005
R50886 VINP.n368 VINP.n193 4.5005
R50887 VINP.n231 VINP.n193 4.5005
R50888 VINP.n370 VINP.n193 4.5005
R50889 VINP.n230 VINP.n193 4.5005
R50890 VINP.n372 VINP.n193 4.5005
R50891 VINP.n229 VINP.n193 4.5005
R50892 VINP.n374 VINP.n193 4.5005
R50893 VINP.n228 VINP.n193 4.5005
R50894 VINP.n376 VINP.n193 4.5005
R50895 VINP.n227 VINP.n193 4.5005
R50896 VINP.n378 VINP.n193 4.5005
R50897 VINP.n226 VINP.n193 4.5005
R50898 VINP.n380 VINP.n193 4.5005
R50899 VINP.n225 VINP.n193 4.5005
R50900 VINP.n382 VINP.n193 4.5005
R50901 VINP.n224 VINP.n193 4.5005
R50902 VINP.n384 VINP.n193 4.5005
R50903 VINP.n223 VINP.n193 4.5005
R50904 VINP.n386 VINP.n193 4.5005
R50905 VINP.n222 VINP.n193 4.5005
R50906 VINP.n388 VINP.n193 4.5005
R50907 VINP.n221 VINP.n193 4.5005
R50908 VINP.n390 VINP.n193 4.5005
R50909 VINP.n220 VINP.n193 4.5005
R50910 VINP.n392 VINP.n193 4.5005
R50911 VINP.n219 VINP.n193 4.5005
R50912 VINP.n394 VINP.n193 4.5005
R50913 VINP.n218 VINP.n193 4.5005
R50914 VINP.n396 VINP.n193 4.5005
R50915 VINP.n217 VINP.n193 4.5005
R50916 VINP.n398 VINP.n193 4.5005
R50917 VINP.n216 VINP.n193 4.5005
R50918 VINP.n400 VINP.n193 4.5005
R50919 VINP.n215 VINP.n193 4.5005
R50920 VINP.n654 VINP.n193 4.5005
R50921 VINP.n656 VINP.n193 4.5005
R50922 VINP.n193 VINP.n0 4.5005
R50923 VINP.n278 VINP.n107 4.5005
R50924 VINP.n276 VINP.n107 4.5005
R50925 VINP.n280 VINP.n107 4.5005
R50926 VINP.n275 VINP.n107 4.5005
R50927 VINP.n282 VINP.n107 4.5005
R50928 VINP.n274 VINP.n107 4.5005
R50929 VINP.n284 VINP.n107 4.5005
R50930 VINP.n273 VINP.n107 4.5005
R50931 VINP.n286 VINP.n107 4.5005
R50932 VINP.n272 VINP.n107 4.5005
R50933 VINP.n288 VINP.n107 4.5005
R50934 VINP.n271 VINP.n107 4.5005
R50935 VINP.n290 VINP.n107 4.5005
R50936 VINP.n270 VINP.n107 4.5005
R50937 VINP.n292 VINP.n107 4.5005
R50938 VINP.n269 VINP.n107 4.5005
R50939 VINP.n294 VINP.n107 4.5005
R50940 VINP.n268 VINP.n107 4.5005
R50941 VINP.n296 VINP.n107 4.5005
R50942 VINP.n267 VINP.n107 4.5005
R50943 VINP.n298 VINP.n107 4.5005
R50944 VINP.n266 VINP.n107 4.5005
R50945 VINP.n300 VINP.n107 4.5005
R50946 VINP.n265 VINP.n107 4.5005
R50947 VINP.n302 VINP.n107 4.5005
R50948 VINP.n264 VINP.n107 4.5005
R50949 VINP.n304 VINP.n107 4.5005
R50950 VINP.n263 VINP.n107 4.5005
R50951 VINP.n306 VINP.n107 4.5005
R50952 VINP.n262 VINP.n107 4.5005
R50953 VINP.n308 VINP.n107 4.5005
R50954 VINP.n261 VINP.n107 4.5005
R50955 VINP.n310 VINP.n107 4.5005
R50956 VINP.n260 VINP.n107 4.5005
R50957 VINP.n312 VINP.n107 4.5005
R50958 VINP.n259 VINP.n107 4.5005
R50959 VINP.n314 VINP.n107 4.5005
R50960 VINP.n258 VINP.n107 4.5005
R50961 VINP.n316 VINP.n107 4.5005
R50962 VINP.n257 VINP.n107 4.5005
R50963 VINP.n318 VINP.n107 4.5005
R50964 VINP.n256 VINP.n107 4.5005
R50965 VINP.n320 VINP.n107 4.5005
R50966 VINP.n255 VINP.n107 4.5005
R50967 VINP.n322 VINP.n107 4.5005
R50968 VINP.n254 VINP.n107 4.5005
R50969 VINP.n324 VINP.n107 4.5005
R50970 VINP.n253 VINP.n107 4.5005
R50971 VINP.n326 VINP.n107 4.5005
R50972 VINP.n252 VINP.n107 4.5005
R50973 VINP.n328 VINP.n107 4.5005
R50974 VINP.n251 VINP.n107 4.5005
R50975 VINP.n330 VINP.n107 4.5005
R50976 VINP.n250 VINP.n107 4.5005
R50977 VINP.n332 VINP.n107 4.5005
R50978 VINP.n249 VINP.n107 4.5005
R50979 VINP.n334 VINP.n107 4.5005
R50980 VINP.n248 VINP.n107 4.5005
R50981 VINP.n336 VINP.n107 4.5005
R50982 VINP.n247 VINP.n107 4.5005
R50983 VINP.n338 VINP.n107 4.5005
R50984 VINP.n246 VINP.n107 4.5005
R50985 VINP.n340 VINP.n107 4.5005
R50986 VINP.n245 VINP.n107 4.5005
R50987 VINP.n342 VINP.n107 4.5005
R50988 VINP.n244 VINP.n107 4.5005
R50989 VINP.n344 VINP.n107 4.5005
R50990 VINP.n243 VINP.n107 4.5005
R50991 VINP.n346 VINP.n107 4.5005
R50992 VINP.n242 VINP.n107 4.5005
R50993 VINP.n348 VINP.n107 4.5005
R50994 VINP.n241 VINP.n107 4.5005
R50995 VINP.n350 VINP.n107 4.5005
R50996 VINP.n240 VINP.n107 4.5005
R50997 VINP.n352 VINP.n107 4.5005
R50998 VINP.n239 VINP.n107 4.5005
R50999 VINP.n354 VINP.n107 4.5005
R51000 VINP.n238 VINP.n107 4.5005
R51001 VINP.n356 VINP.n107 4.5005
R51002 VINP.n237 VINP.n107 4.5005
R51003 VINP.n358 VINP.n107 4.5005
R51004 VINP.n236 VINP.n107 4.5005
R51005 VINP.n360 VINP.n107 4.5005
R51006 VINP.n235 VINP.n107 4.5005
R51007 VINP.n362 VINP.n107 4.5005
R51008 VINP.n234 VINP.n107 4.5005
R51009 VINP.n364 VINP.n107 4.5005
R51010 VINP.n233 VINP.n107 4.5005
R51011 VINP.n366 VINP.n107 4.5005
R51012 VINP.n232 VINP.n107 4.5005
R51013 VINP.n368 VINP.n107 4.5005
R51014 VINP.n231 VINP.n107 4.5005
R51015 VINP.n370 VINP.n107 4.5005
R51016 VINP.n230 VINP.n107 4.5005
R51017 VINP.n372 VINP.n107 4.5005
R51018 VINP.n229 VINP.n107 4.5005
R51019 VINP.n374 VINP.n107 4.5005
R51020 VINP.n228 VINP.n107 4.5005
R51021 VINP.n376 VINP.n107 4.5005
R51022 VINP.n227 VINP.n107 4.5005
R51023 VINP.n378 VINP.n107 4.5005
R51024 VINP.n226 VINP.n107 4.5005
R51025 VINP.n380 VINP.n107 4.5005
R51026 VINP.n225 VINP.n107 4.5005
R51027 VINP.n382 VINP.n107 4.5005
R51028 VINP.n224 VINP.n107 4.5005
R51029 VINP.n384 VINP.n107 4.5005
R51030 VINP.n223 VINP.n107 4.5005
R51031 VINP.n386 VINP.n107 4.5005
R51032 VINP.n222 VINP.n107 4.5005
R51033 VINP.n388 VINP.n107 4.5005
R51034 VINP.n221 VINP.n107 4.5005
R51035 VINP.n390 VINP.n107 4.5005
R51036 VINP.n220 VINP.n107 4.5005
R51037 VINP.n392 VINP.n107 4.5005
R51038 VINP.n219 VINP.n107 4.5005
R51039 VINP.n394 VINP.n107 4.5005
R51040 VINP.n218 VINP.n107 4.5005
R51041 VINP.n396 VINP.n107 4.5005
R51042 VINP.n217 VINP.n107 4.5005
R51043 VINP.n398 VINP.n107 4.5005
R51044 VINP.n216 VINP.n107 4.5005
R51045 VINP.n400 VINP.n107 4.5005
R51046 VINP.n215 VINP.n107 4.5005
R51047 VINP.n654 VINP.n107 4.5005
R51048 VINP.n656 VINP.n107 4.5005
R51049 VINP.n107 VINP.n0 4.5005
R51050 VINP.n278 VINP.n194 4.5005
R51051 VINP.n276 VINP.n194 4.5005
R51052 VINP.n280 VINP.n194 4.5005
R51053 VINP.n275 VINP.n194 4.5005
R51054 VINP.n282 VINP.n194 4.5005
R51055 VINP.n274 VINP.n194 4.5005
R51056 VINP.n284 VINP.n194 4.5005
R51057 VINP.n273 VINP.n194 4.5005
R51058 VINP.n286 VINP.n194 4.5005
R51059 VINP.n272 VINP.n194 4.5005
R51060 VINP.n288 VINP.n194 4.5005
R51061 VINP.n271 VINP.n194 4.5005
R51062 VINP.n290 VINP.n194 4.5005
R51063 VINP.n270 VINP.n194 4.5005
R51064 VINP.n292 VINP.n194 4.5005
R51065 VINP.n269 VINP.n194 4.5005
R51066 VINP.n294 VINP.n194 4.5005
R51067 VINP.n268 VINP.n194 4.5005
R51068 VINP.n296 VINP.n194 4.5005
R51069 VINP.n267 VINP.n194 4.5005
R51070 VINP.n298 VINP.n194 4.5005
R51071 VINP.n266 VINP.n194 4.5005
R51072 VINP.n300 VINP.n194 4.5005
R51073 VINP.n265 VINP.n194 4.5005
R51074 VINP.n302 VINP.n194 4.5005
R51075 VINP.n264 VINP.n194 4.5005
R51076 VINP.n304 VINP.n194 4.5005
R51077 VINP.n263 VINP.n194 4.5005
R51078 VINP.n306 VINP.n194 4.5005
R51079 VINP.n262 VINP.n194 4.5005
R51080 VINP.n308 VINP.n194 4.5005
R51081 VINP.n261 VINP.n194 4.5005
R51082 VINP.n310 VINP.n194 4.5005
R51083 VINP.n260 VINP.n194 4.5005
R51084 VINP.n312 VINP.n194 4.5005
R51085 VINP.n259 VINP.n194 4.5005
R51086 VINP.n314 VINP.n194 4.5005
R51087 VINP.n258 VINP.n194 4.5005
R51088 VINP.n316 VINP.n194 4.5005
R51089 VINP.n257 VINP.n194 4.5005
R51090 VINP.n318 VINP.n194 4.5005
R51091 VINP.n256 VINP.n194 4.5005
R51092 VINP.n320 VINP.n194 4.5005
R51093 VINP.n255 VINP.n194 4.5005
R51094 VINP.n322 VINP.n194 4.5005
R51095 VINP.n254 VINP.n194 4.5005
R51096 VINP.n324 VINP.n194 4.5005
R51097 VINP.n253 VINP.n194 4.5005
R51098 VINP.n326 VINP.n194 4.5005
R51099 VINP.n252 VINP.n194 4.5005
R51100 VINP.n328 VINP.n194 4.5005
R51101 VINP.n251 VINP.n194 4.5005
R51102 VINP.n330 VINP.n194 4.5005
R51103 VINP.n250 VINP.n194 4.5005
R51104 VINP.n332 VINP.n194 4.5005
R51105 VINP.n249 VINP.n194 4.5005
R51106 VINP.n334 VINP.n194 4.5005
R51107 VINP.n248 VINP.n194 4.5005
R51108 VINP.n336 VINP.n194 4.5005
R51109 VINP.n247 VINP.n194 4.5005
R51110 VINP.n338 VINP.n194 4.5005
R51111 VINP.n246 VINP.n194 4.5005
R51112 VINP.n340 VINP.n194 4.5005
R51113 VINP.n245 VINP.n194 4.5005
R51114 VINP.n342 VINP.n194 4.5005
R51115 VINP.n244 VINP.n194 4.5005
R51116 VINP.n344 VINP.n194 4.5005
R51117 VINP.n243 VINP.n194 4.5005
R51118 VINP.n346 VINP.n194 4.5005
R51119 VINP.n242 VINP.n194 4.5005
R51120 VINP.n348 VINP.n194 4.5005
R51121 VINP.n241 VINP.n194 4.5005
R51122 VINP.n350 VINP.n194 4.5005
R51123 VINP.n240 VINP.n194 4.5005
R51124 VINP.n352 VINP.n194 4.5005
R51125 VINP.n239 VINP.n194 4.5005
R51126 VINP.n354 VINP.n194 4.5005
R51127 VINP.n238 VINP.n194 4.5005
R51128 VINP.n356 VINP.n194 4.5005
R51129 VINP.n237 VINP.n194 4.5005
R51130 VINP.n358 VINP.n194 4.5005
R51131 VINP.n236 VINP.n194 4.5005
R51132 VINP.n360 VINP.n194 4.5005
R51133 VINP.n235 VINP.n194 4.5005
R51134 VINP.n362 VINP.n194 4.5005
R51135 VINP.n234 VINP.n194 4.5005
R51136 VINP.n364 VINP.n194 4.5005
R51137 VINP.n233 VINP.n194 4.5005
R51138 VINP.n366 VINP.n194 4.5005
R51139 VINP.n232 VINP.n194 4.5005
R51140 VINP.n368 VINP.n194 4.5005
R51141 VINP.n231 VINP.n194 4.5005
R51142 VINP.n370 VINP.n194 4.5005
R51143 VINP.n230 VINP.n194 4.5005
R51144 VINP.n372 VINP.n194 4.5005
R51145 VINP.n229 VINP.n194 4.5005
R51146 VINP.n374 VINP.n194 4.5005
R51147 VINP.n228 VINP.n194 4.5005
R51148 VINP.n376 VINP.n194 4.5005
R51149 VINP.n227 VINP.n194 4.5005
R51150 VINP.n378 VINP.n194 4.5005
R51151 VINP.n226 VINP.n194 4.5005
R51152 VINP.n380 VINP.n194 4.5005
R51153 VINP.n225 VINP.n194 4.5005
R51154 VINP.n382 VINP.n194 4.5005
R51155 VINP.n224 VINP.n194 4.5005
R51156 VINP.n384 VINP.n194 4.5005
R51157 VINP.n223 VINP.n194 4.5005
R51158 VINP.n386 VINP.n194 4.5005
R51159 VINP.n222 VINP.n194 4.5005
R51160 VINP.n388 VINP.n194 4.5005
R51161 VINP.n221 VINP.n194 4.5005
R51162 VINP.n390 VINP.n194 4.5005
R51163 VINP.n220 VINP.n194 4.5005
R51164 VINP.n392 VINP.n194 4.5005
R51165 VINP.n219 VINP.n194 4.5005
R51166 VINP.n394 VINP.n194 4.5005
R51167 VINP.n218 VINP.n194 4.5005
R51168 VINP.n396 VINP.n194 4.5005
R51169 VINP.n217 VINP.n194 4.5005
R51170 VINP.n398 VINP.n194 4.5005
R51171 VINP.n216 VINP.n194 4.5005
R51172 VINP.n400 VINP.n194 4.5005
R51173 VINP.n215 VINP.n194 4.5005
R51174 VINP.n654 VINP.n194 4.5005
R51175 VINP.n656 VINP.n194 4.5005
R51176 VINP.n194 VINP.n0 4.5005
R51177 VINP.n278 VINP.n106 4.5005
R51178 VINP.n276 VINP.n106 4.5005
R51179 VINP.n280 VINP.n106 4.5005
R51180 VINP.n275 VINP.n106 4.5005
R51181 VINP.n282 VINP.n106 4.5005
R51182 VINP.n274 VINP.n106 4.5005
R51183 VINP.n284 VINP.n106 4.5005
R51184 VINP.n273 VINP.n106 4.5005
R51185 VINP.n286 VINP.n106 4.5005
R51186 VINP.n272 VINP.n106 4.5005
R51187 VINP.n288 VINP.n106 4.5005
R51188 VINP.n271 VINP.n106 4.5005
R51189 VINP.n290 VINP.n106 4.5005
R51190 VINP.n270 VINP.n106 4.5005
R51191 VINP.n292 VINP.n106 4.5005
R51192 VINP.n269 VINP.n106 4.5005
R51193 VINP.n294 VINP.n106 4.5005
R51194 VINP.n268 VINP.n106 4.5005
R51195 VINP.n296 VINP.n106 4.5005
R51196 VINP.n267 VINP.n106 4.5005
R51197 VINP.n298 VINP.n106 4.5005
R51198 VINP.n266 VINP.n106 4.5005
R51199 VINP.n300 VINP.n106 4.5005
R51200 VINP.n265 VINP.n106 4.5005
R51201 VINP.n302 VINP.n106 4.5005
R51202 VINP.n264 VINP.n106 4.5005
R51203 VINP.n304 VINP.n106 4.5005
R51204 VINP.n263 VINP.n106 4.5005
R51205 VINP.n306 VINP.n106 4.5005
R51206 VINP.n262 VINP.n106 4.5005
R51207 VINP.n308 VINP.n106 4.5005
R51208 VINP.n261 VINP.n106 4.5005
R51209 VINP.n310 VINP.n106 4.5005
R51210 VINP.n260 VINP.n106 4.5005
R51211 VINP.n312 VINP.n106 4.5005
R51212 VINP.n259 VINP.n106 4.5005
R51213 VINP.n314 VINP.n106 4.5005
R51214 VINP.n258 VINP.n106 4.5005
R51215 VINP.n316 VINP.n106 4.5005
R51216 VINP.n257 VINP.n106 4.5005
R51217 VINP.n318 VINP.n106 4.5005
R51218 VINP.n256 VINP.n106 4.5005
R51219 VINP.n320 VINP.n106 4.5005
R51220 VINP.n255 VINP.n106 4.5005
R51221 VINP.n322 VINP.n106 4.5005
R51222 VINP.n254 VINP.n106 4.5005
R51223 VINP.n324 VINP.n106 4.5005
R51224 VINP.n253 VINP.n106 4.5005
R51225 VINP.n326 VINP.n106 4.5005
R51226 VINP.n252 VINP.n106 4.5005
R51227 VINP.n328 VINP.n106 4.5005
R51228 VINP.n251 VINP.n106 4.5005
R51229 VINP.n330 VINP.n106 4.5005
R51230 VINP.n250 VINP.n106 4.5005
R51231 VINP.n332 VINP.n106 4.5005
R51232 VINP.n249 VINP.n106 4.5005
R51233 VINP.n334 VINP.n106 4.5005
R51234 VINP.n248 VINP.n106 4.5005
R51235 VINP.n336 VINP.n106 4.5005
R51236 VINP.n247 VINP.n106 4.5005
R51237 VINP.n338 VINP.n106 4.5005
R51238 VINP.n246 VINP.n106 4.5005
R51239 VINP.n340 VINP.n106 4.5005
R51240 VINP.n245 VINP.n106 4.5005
R51241 VINP.n342 VINP.n106 4.5005
R51242 VINP.n244 VINP.n106 4.5005
R51243 VINP.n344 VINP.n106 4.5005
R51244 VINP.n243 VINP.n106 4.5005
R51245 VINP.n346 VINP.n106 4.5005
R51246 VINP.n242 VINP.n106 4.5005
R51247 VINP.n348 VINP.n106 4.5005
R51248 VINP.n241 VINP.n106 4.5005
R51249 VINP.n350 VINP.n106 4.5005
R51250 VINP.n240 VINP.n106 4.5005
R51251 VINP.n352 VINP.n106 4.5005
R51252 VINP.n239 VINP.n106 4.5005
R51253 VINP.n354 VINP.n106 4.5005
R51254 VINP.n238 VINP.n106 4.5005
R51255 VINP.n356 VINP.n106 4.5005
R51256 VINP.n237 VINP.n106 4.5005
R51257 VINP.n358 VINP.n106 4.5005
R51258 VINP.n236 VINP.n106 4.5005
R51259 VINP.n360 VINP.n106 4.5005
R51260 VINP.n235 VINP.n106 4.5005
R51261 VINP.n362 VINP.n106 4.5005
R51262 VINP.n234 VINP.n106 4.5005
R51263 VINP.n364 VINP.n106 4.5005
R51264 VINP.n233 VINP.n106 4.5005
R51265 VINP.n366 VINP.n106 4.5005
R51266 VINP.n232 VINP.n106 4.5005
R51267 VINP.n368 VINP.n106 4.5005
R51268 VINP.n231 VINP.n106 4.5005
R51269 VINP.n370 VINP.n106 4.5005
R51270 VINP.n230 VINP.n106 4.5005
R51271 VINP.n372 VINP.n106 4.5005
R51272 VINP.n229 VINP.n106 4.5005
R51273 VINP.n374 VINP.n106 4.5005
R51274 VINP.n228 VINP.n106 4.5005
R51275 VINP.n376 VINP.n106 4.5005
R51276 VINP.n227 VINP.n106 4.5005
R51277 VINP.n378 VINP.n106 4.5005
R51278 VINP.n226 VINP.n106 4.5005
R51279 VINP.n380 VINP.n106 4.5005
R51280 VINP.n225 VINP.n106 4.5005
R51281 VINP.n382 VINP.n106 4.5005
R51282 VINP.n224 VINP.n106 4.5005
R51283 VINP.n384 VINP.n106 4.5005
R51284 VINP.n223 VINP.n106 4.5005
R51285 VINP.n386 VINP.n106 4.5005
R51286 VINP.n222 VINP.n106 4.5005
R51287 VINP.n388 VINP.n106 4.5005
R51288 VINP.n221 VINP.n106 4.5005
R51289 VINP.n390 VINP.n106 4.5005
R51290 VINP.n220 VINP.n106 4.5005
R51291 VINP.n392 VINP.n106 4.5005
R51292 VINP.n219 VINP.n106 4.5005
R51293 VINP.n394 VINP.n106 4.5005
R51294 VINP.n218 VINP.n106 4.5005
R51295 VINP.n396 VINP.n106 4.5005
R51296 VINP.n217 VINP.n106 4.5005
R51297 VINP.n398 VINP.n106 4.5005
R51298 VINP.n216 VINP.n106 4.5005
R51299 VINP.n400 VINP.n106 4.5005
R51300 VINP.n215 VINP.n106 4.5005
R51301 VINP.n654 VINP.n106 4.5005
R51302 VINP.n656 VINP.n106 4.5005
R51303 VINP.n106 VINP.n0 4.5005
R51304 VINP.n278 VINP.n195 4.5005
R51305 VINP.n276 VINP.n195 4.5005
R51306 VINP.n280 VINP.n195 4.5005
R51307 VINP.n275 VINP.n195 4.5005
R51308 VINP.n282 VINP.n195 4.5005
R51309 VINP.n274 VINP.n195 4.5005
R51310 VINP.n284 VINP.n195 4.5005
R51311 VINP.n273 VINP.n195 4.5005
R51312 VINP.n286 VINP.n195 4.5005
R51313 VINP.n272 VINP.n195 4.5005
R51314 VINP.n288 VINP.n195 4.5005
R51315 VINP.n271 VINP.n195 4.5005
R51316 VINP.n290 VINP.n195 4.5005
R51317 VINP.n270 VINP.n195 4.5005
R51318 VINP.n292 VINP.n195 4.5005
R51319 VINP.n269 VINP.n195 4.5005
R51320 VINP.n294 VINP.n195 4.5005
R51321 VINP.n268 VINP.n195 4.5005
R51322 VINP.n296 VINP.n195 4.5005
R51323 VINP.n267 VINP.n195 4.5005
R51324 VINP.n298 VINP.n195 4.5005
R51325 VINP.n266 VINP.n195 4.5005
R51326 VINP.n300 VINP.n195 4.5005
R51327 VINP.n265 VINP.n195 4.5005
R51328 VINP.n302 VINP.n195 4.5005
R51329 VINP.n264 VINP.n195 4.5005
R51330 VINP.n304 VINP.n195 4.5005
R51331 VINP.n263 VINP.n195 4.5005
R51332 VINP.n306 VINP.n195 4.5005
R51333 VINP.n262 VINP.n195 4.5005
R51334 VINP.n308 VINP.n195 4.5005
R51335 VINP.n261 VINP.n195 4.5005
R51336 VINP.n310 VINP.n195 4.5005
R51337 VINP.n260 VINP.n195 4.5005
R51338 VINP.n312 VINP.n195 4.5005
R51339 VINP.n259 VINP.n195 4.5005
R51340 VINP.n314 VINP.n195 4.5005
R51341 VINP.n258 VINP.n195 4.5005
R51342 VINP.n316 VINP.n195 4.5005
R51343 VINP.n257 VINP.n195 4.5005
R51344 VINP.n318 VINP.n195 4.5005
R51345 VINP.n256 VINP.n195 4.5005
R51346 VINP.n320 VINP.n195 4.5005
R51347 VINP.n255 VINP.n195 4.5005
R51348 VINP.n322 VINP.n195 4.5005
R51349 VINP.n254 VINP.n195 4.5005
R51350 VINP.n324 VINP.n195 4.5005
R51351 VINP.n253 VINP.n195 4.5005
R51352 VINP.n326 VINP.n195 4.5005
R51353 VINP.n252 VINP.n195 4.5005
R51354 VINP.n328 VINP.n195 4.5005
R51355 VINP.n251 VINP.n195 4.5005
R51356 VINP.n330 VINP.n195 4.5005
R51357 VINP.n250 VINP.n195 4.5005
R51358 VINP.n332 VINP.n195 4.5005
R51359 VINP.n249 VINP.n195 4.5005
R51360 VINP.n334 VINP.n195 4.5005
R51361 VINP.n248 VINP.n195 4.5005
R51362 VINP.n336 VINP.n195 4.5005
R51363 VINP.n247 VINP.n195 4.5005
R51364 VINP.n338 VINP.n195 4.5005
R51365 VINP.n246 VINP.n195 4.5005
R51366 VINP.n340 VINP.n195 4.5005
R51367 VINP.n245 VINP.n195 4.5005
R51368 VINP.n342 VINP.n195 4.5005
R51369 VINP.n244 VINP.n195 4.5005
R51370 VINP.n344 VINP.n195 4.5005
R51371 VINP.n243 VINP.n195 4.5005
R51372 VINP.n346 VINP.n195 4.5005
R51373 VINP.n242 VINP.n195 4.5005
R51374 VINP.n348 VINP.n195 4.5005
R51375 VINP.n241 VINP.n195 4.5005
R51376 VINP.n350 VINP.n195 4.5005
R51377 VINP.n240 VINP.n195 4.5005
R51378 VINP.n352 VINP.n195 4.5005
R51379 VINP.n239 VINP.n195 4.5005
R51380 VINP.n354 VINP.n195 4.5005
R51381 VINP.n238 VINP.n195 4.5005
R51382 VINP.n356 VINP.n195 4.5005
R51383 VINP.n237 VINP.n195 4.5005
R51384 VINP.n358 VINP.n195 4.5005
R51385 VINP.n236 VINP.n195 4.5005
R51386 VINP.n360 VINP.n195 4.5005
R51387 VINP.n235 VINP.n195 4.5005
R51388 VINP.n362 VINP.n195 4.5005
R51389 VINP.n234 VINP.n195 4.5005
R51390 VINP.n364 VINP.n195 4.5005
R51391 VINP.n233 VINP.n195 4.5005
R51392 VINP.n366 VINP.n195 4.5005
R51393 VINP.n232 VINP.n195 4.5005
R51394 VINP.n368 VINP.n195 4.5005
R51395 VINP.n231 VINP.n195 4.5005
R51396 VINP.n370 VINP.n195 4.5005
R51397 VINP.n230 VINP.n195 4.5005
R51398 VINP.n372 VINP.n195 4.5005
R51399 VINP.n229 VINP.n195 4.5005
R51400 VINP.n374 VINP.n195 4.5005
R51401 VINP.n228 VINP.n195 4.5005
R51402 VINP.n376 VINP.n195 4.5005
R51403 VINP.n227 VINP.n195 4.5005
R51404 VINP.n378 VINP.n195 4.5005
R51405 VINP.n226 VINP.n195 4.5005
R51406 VINP.n380 VINP.n195 4.5005
R51407 VINP.n225 VINP.n195 4.5005
R51408 VINP.n382 VINP.n195 4.5005
R51409 VINP.n224 VINP.n195 4.5005
R51410 VINP.n384 VINP.n195 4.5005
R51411 VINP.n223 VINP.n195 4.5005
R51412 VINP.n386 VINP.n195 4.5005
R51413 VINP.n222 VINP.n195 4.5005
R51414 VINP.n388 VINP.n195 4.5005
R51415 VINP.n221 VINP.n195 4.5005
R51416 VINP.n390 VINP.n195 4.5005
R51417 VINP.n220 VINP.n195 4.5005
R51418 VINP.n392 VINP.n195 4.5005
R51419 VINP.n219 VINP.n195 4.5005
R51420 VINP.n394 VINP.n195 4.5005
R51421 VINP.n218 VINP.n195 4.5005
R51422 VINP.n396 VINP.n195 4.5005
R51423 VINP.n217 VINP.n195 4.5005
R51424 VINP.n398 VINP.n195 4.5005
R51425 VINP.n216 VINP.n195 4.5005
R51426 VINP.n400 VINP.n195 4.5005
R51427 VINP.n215 VINP.n195 4.5005
R51428 VINP.n654 VINP.n195 4.5005
R51429 VINP.n656 VINP.n195 4.5005
R51430 VINP.n195 VINP.n0 4.5005
R51431 VINP.n278 VINP.n105 4.5005
R51432 VINP.n276 VINP.n105 4.5005
R51433 VINP.n280 VINP.n105 4.5005
R51434 VINP.n275 VINP.n105 4.5005
R51435 VINP.n282 VINP.n105 4.5005
R51436 VINP.n274 VINP.n105 4.5005
R51437 VINP.n284 VINP.n105 4.5005
R51438 VINP.n273 VINP.n105 4.5005
R51439 VINP.n286 VINP.n105 4.5005
R51440 VINP.n272 VINP.n105 4.5005
R51441 VINP.n288 VINP.n105 4.5005
R51442 VINP.n271 VINP.n105 4.5005
R51443 VINP.n290 VINP.n105 4.5005
R51444 VINP.n270 VINP.n105 4.5005
R51445 VINP.n292 VINP.n105 4.5005
R51446 VINP.n269 VINP.n105 4.5005
R51447 VINP.n294 VINP.n105 4.5005
R51448 VINP.n268 VINP.n105 4.5005
R51449 VINP.n296 VINP.n105 4.5005
R51450 VINP.n267 VINP.n105 4.5005
R51451 VINP.n298 VINP.n105 4.5005
R51452 VINP.n266 VINP.n105 4.5005
R51453 VINP.n300 VINP.n105 4.5005
R51454 VINP.n265 VINP.n105 4.5005
R51455 VINP.n302 VINP.n105 4.5005
R51456 VINP.n264 VINP.n105 4.5005
R51457 VINP.n304 VINP.n105 4.5005
R51458 VINP.n263 VINP.n105 4.5005
R51459 VINP.n306 VINP.n105 4.5005
R51460 VINP.n262 VINP.n105 4.5005
R51461 VINP.n308 VINP.n105 4.5005
R51462 VINP.n261 VINP.n105 4.5005
R51463 VINP.n310 VINP.n105 4.5005
R51464 VINP.n260 VINP.n105 4.5005
R51465 VINP.n312 VINP.n105 4.5005
R51466 VINP.n259 VINP.n105 4.5005
R51467 VINP.n314 VINP.n105 4.5005
R51468 VINP.n258 VINP.n105 4.5005
R51469 VINP.n316 VINP.n105 4.5005
R51470 VINP.n257 VINP.n105 4.5005
R51471 VINP.n318 VINP.n105 4.5005
R51472 VINP.n256 VINP.n105 4.5005
R51473 VINP.n320 VINP.n105 4.5005
R51474 VINP.n255 VINP.n105 4.5005
R51475 VINP.n322 VINP.n105 4.5005
R51476 VINP.n254 VINP.n105 4.5005
R51477 VINP.n324 VINP.n105 4.5005
R51478 VINP.n253 VINP.n105 4.5005
R51479 VINP.n326 VINP.n105 4.5005
R51480 VINP.n252 VINP.n105 4.5005
R51481 VINP.n328 VINP.n105 4.5005
R51482 VINP.n251 VINP.n105 4.5005
R51483 VINP.n330 VINP.n105 4.5005
R51484 VINP.n250 VINP.n105 4.5005
R51485 VINP.n332 VINP.n105 4.5005
R51486 VINP.n249 VINP.n105 4.5005
R51487 VINP.n334 VINP.n105 4.5005
R51488 VINP.n248 VINP.n105 4.5005
R51489 VINP.n336 VINP.n105 4.5005
R51490 VINP.n247 VINP.n105 4.5005
R51491 VINP.n338 VINP.n105 4.5005
R51492 VINP.n246 VINP.n105 4.5005
R51493 VINP.n340 VINP.n105 4.5005
R51494 VINP.n245 VINP.n105 4.5005
R51495 VINP.n342 VINP.n105 4.5005
R51496 VINP.n244 VINP.n105 4.5005
R51497 VINP.n344 VINP.n105 4.5005
R51498 VINP.n243 VINP.n105 4.5005
R51499 VINP.n346 VINP.n105 4.5005
R51500 VINP.n242 VINP.n105 4.5005
R51501 VINP.n348 VINP.n105 4.5005
R51502 VINP.n241 VINP.n105 4.5005
R51503 VINP.n350 VINP.n105 4.5005
R51504 VINP.n240 VINP.n105 4.5005
R51505 VINP.n352 VINP.n105 4.5005
R51506 VINP.n239 VINP.n105 4.5005
R51507 VINP.n354 VINP.n105 4.5005
R51508 VINP.n238 VINP.n105 4.5005
R51509 VINP.n356 VINP.n105 4.5005
R51510 VINP.n237 VINP.n105 4.5005
R51511 VINP.n358 VINP.n105 4.5005
R51512 VINP.n236 VINP.n105 4.5005
R51513 VINP.n360 VINP.n105 4.5005
R51514 VINP.n235 VINP.n105 4.5005
R51515 VINP.n362 VINP.n105 4.5005
R51516 VINP.n234 VINP.n105 4.5005
R51517 VINP.n364 VINP.n105 4.5005
R51518 VINP.n233 VINP.n105 4.5005
R51519 VINP.n366 VINP.n105 4.5005
R51520 VINP.n232 VINP.n105 4.5005
R51521 VINP.n368 VINP.n105 4.5005
R51522 VINP.n231 VINP.n105 4.5005
R51523 VINP.n370 VINP.n105 4.5005
R51524 VINP.n230 VINP.n105 4.5005
R51525 VINP.n372 VINP.n105 4.5005
R51526 VINP.n229 VINP.n105 4.5005
R51527 VINP.n374 VINP.n105 4.5005
R51528 VINP.n228 VINP.n105 4.5005
R51529 VINP.n376 VINP.n105 4.5005
R51530 VINP.n227 VINP.n105 4.5005
R51531 VINP.n378 VINP.n105 4.5005
R51532 VINP.n226 VINP.n105 4.5005
R51533 VINP.n380 VINP.n105 4.5005
R51534 VINP.n225 VINP.n105 4.5005
R51535 VINP.n382 VINP.n105 4.5005
R51536 VINP.n224 VINP.n105 4.5005
R51537 VINP.n384 VINP.n105 4.5005
R51538 VINP.n223 VINP.n105 4.5005
R51539 VINP.n386 VINP.n105 4.5005
R51540 VINP.n222 VINP.n105 4.5005
R51541 VINP.n388 VINP.n105 4.5005
R51542 VINP.n221 VINP.n105 4.5005
R51543 VINP.n390 VINP.n105 4.5005
R51544 VINP.n220 VINP.n105 4.5005
R51545 VINP.n392 VINP.n105 4.5005
R51546 VINP.n219 VINP.n105 4.5005
R51547 VINP.n394 VINP.n105 4.5005
R51548 VINP.n218 VINP.n105 4.5005
R51549 VINP.n396 VINP.n105 4.5005
R51550 VINP.n217 VINP.n105 4.5005
R51551 VINP.n398 VINP.n105 4.5005
R51552 VINP.n216 VINP.n105 4.5005
R51553 VINP.n400 VINP.n105 4.5005
R51554 VINP.n215 VINP.n105 4.5005
R51555 VINP.n654 VINP.n105 4.5005
R51556 VINP.n656 VINP.n105 4.5005
R51557 VINP.n105 VINP.n0 4.5005
R51558 VINP.n278 VINP.n196 4.5005
R51559 VINP.n276 VINP.n196 4.5005
R51560 VINP.n280 VINP.n196 4.5005
R51561 VINP.n275 VINP.n196 4.5005
R51562 VINP.n282 VINP.n196 4.5005
R51563 VINP.n274 VINP.n196 4.5005
R51564 VINP.n284 VINP.n196 4.5005
R51565 VINP.n273 VINP.n196 4.5005
R51566 VINP.n286 VINP.n196 4.5005
R51567 VINP.n272 VINP.n196 4.5005
R51568 VINP.n288 VINP.n196 4.5005
R51569 VINP.n271 VINP.n196 4.5005
R51570 VINP.n290 VINP.n196 4.5005
R51571 VINP.n270 VINP.n196 4.5005
R51572 VINP.n292 VINP.n196 4.5005
R51573 VINP.n269 VINP.n196 4.5005
R51574 VINP.n294 VINP.n196 4.5005
R51575 VINP.n268 VINP.n196 4.5005
R51576 VINP.n296 VINP.n196 4.5005
R51577 VINP.n267 VINP.n196 4.5005
R51578 VINP.n298 VINP.n196 4.5005
R51579 VINP.n266 VINP.n196 4.5005
R51580 VINP.n300 VINP.n196 4.5005
R51581 VINP.n265 VINP.n196 4.5005
R51582 VINP.n302 VINP.n196 4.5005
R51583 VINP.n264 VINP.n196 4.5005
R51584 VINP.n304 VINP.n196 4.5005
R51585 VINP.n263 VINP.n196 4.5005
R51586 VINP.n306 VINP.n196 4.5005
R51587 VINP.n262 VINP.n196 4.5005
R51588 VINP.n308 VINP.n196 4.5005
R51589 VINP.n261 VINP.n196 4.5005
R51590 VINP.n310 VINP.n196 4.5005
R51591 VINP.n260 VINP.n196 4.5005
R51592 VINP.n312 VINP.n196 4.5005
R51593 VINP.n259 VINP.n196 4.5005
R51594 VINP.n314 VINP.n196 4.5005
R51595 VINP.n258 VINP.n196 4.5005
R51596 VINP.n316 VINP.n196 4.5005
R51597 VINP.n257 VINP.n196 4.5005
R51598 VINP.n318 VINP.n196 4.5005
R51599 VINP.n256 VINP.n196 4.5005
R51600 VINP.n320 VINP.n196 4.5005
R51601 VINP.n255 VINP.n196 4.5005
R51602 VINP.n322 VINP.n196 4.5005
R51603 VINP.n254 VINP.n196 4.5005
R51604 VINP.n324 VINP.n196 4.5005
R51605 VINP.n253 VINP.n196 4.5005
R51606 VINP.n326 VINP.n196 4.5005
R51607 VINP.n252 VINP.n196 4.5005
R51608 VINP.n328 VINP.n196 4.5005
R51609 VINP.n251 VINP.n196 4.5005
R51610 VINP.n330 VINP.n196 4.5005
R51611 VINP.n250 VINP.n196 4.5005
R51612 VINP.n332 VINP.n196 4.5005
R51613 VINP.n249 VINP.n196 4.5005
R51614 VINP.n334 VINP.n196 4.5005
R51615 VINP.n248 VINP.n196 4.5005
R51616 VINP.n336 VINP.n196 4.5005
R51617 VINP.n247 VINP.n196 4.5005
R51618 VINP.n338 VINP.n196 4.5005
R51619 VINP.n246 VINP.n196 4.5005
R51620 VINP.n340 VINP.n196 4.5005
R51621 VINP.n245 VINP.n196 4.5005
R51622 VINP.n342 VINP.n196 4.5005
R51623 VINP.n244 VINP.n196 4.5005
R51624 VINP.n344 VINP.n196 4.5005
R51625 VINP.n243 VINP.n196 4.5005
R51626 VINP.n346 VINP.n196 4.5005
R51627 VINP.n242 VINP.n196 4.5005
R51628 VINP.n348 VINP.n196 4.5005
R51629 VINP.n241 VINP.n196 4.5005
R51630 VINP.n350 VINP.n196 4.5005
R51631 VINP.n240 VINP.n196 4.5005
R51632 VINP.n352 VINP.n196 4.5005
R51633 VINP.n239 VINP.n196 4.5005
R51634 VINP.n354 VINP.n196 4.5005
R51635 VINP.n238 VINP.n196 4.5005
R51636 VINP.n356 VINP.n196 4.5005
R51637 VINP.n237 VINP.n196 4.5005
R51638 VINP.n358 VINP.n196 4.5005
R51639 VINP.n236 VINP.n196 4.5005
R51640 VINP.n360 VINP.n196 4.5005
R51641 VINP.n235 VINP.n196 4.5005
R51642 VINP.n362 VINP.n196 4.5005
R51643 VINP.n234 VINP.n196 4.5005
R51644 VINP.n364 VINP.n196 4.5005
R51645 VINP.n233 VINP.n196 4.5005
R51646 VINP.n366 VINP.n196 4.5005
R51647 VINP.n232 VINP.n196 4.5005
R51648 VINP.n368 VINP.n196 4.5005
R51649 VINP.n231 VINP.n196 4.5005
R51650 VINP.n370 VINP.n196 4.5005
R51651 VINP.n230 VINP.n196 4.5005
R51652 VINP.n372 VINP.n196 4.5005
R51653 VINP.n229 VINP.n196 4.5005
R51654 VINP.n374 VINP.n196 4.5005
R51655 VINP.n228 VINP.n196 4.5005
R51656 VINP.n376 VINP.n196 4.5005
R51657 VINP.n227 VINP.n196 4.5005
R51658 VINP.n378 VINP.n196 4.5005
R51659 VINP.n226 VINP.n196 4.5005
R51660 VINP.n380 VINP.n196 4.5005
R51661 VINP.n225 VINP.n196 4.5005
R51662 VINP.n382 VINP.n196 4.5005
R51663 VINP.n224 VINP.n196 4.5005
R51664 VINP.n384 VINP.n196 4.5005
R51665 VINP.n223 VINP.n196 4.5005
R51666 VINP.n386 VINP.n196 4.5005
R51667 VINP.n222 VINP.n196 4.5005
R51668 VINP.n388 VINP.n196 4.5005
R51669 VINP.n221 VINP.n196 4.5005
R51670 VINP.n390 VINP.n196 4.5005
R51671 VINP.n220 VINP.n196 4.5005
R51672 VINP.n392 VINP.n196 4.5005
R51673 VINP.n219 VINP.n196 4.5005
R51674 VINP.n394 VINP.n196 4.5005
R51675 VINP.n218 VINP.n196 4.5005
R51676 VINP.n396 VINP.n196 4.5005
R51677 VINP.n217 VINP.n196 4.5005
R51678 VINP.n398 VINP.n196 4.5005
R51679 VINP.n216 VINP.n196 4.5005
R51680 VINP.n400 VINP.n196 4.5005
R51681 VINP.n215 VINP.n196 4.5005
R51682 VINP.n654 VINP.n196 4.5005
R51683 VINP.n656 VINP.n196 4.5005
R51684 VINP.n196 VINP.n0 4.5005
R51685 VINP.n278 VINP.n104 4.5005
R51686 VINP.n276 VINP.n104 4.5005
R51687 VINP.n280 VINP.n104 4.5005
R51688 VINP.n275 VINP.n104 4.5005
R51689 VINP.n282 VINP.n104 4.5005
R51690 VINP.n274 VINP.n104 4.5005
R51691 VINP.n284 VINP.n104 4.5005
R51692 VINP.n273 VINP.n104 4.5005
R51693 VINP.n286 VINP.n104 4.5005
R51694 VINP.n272 VINP.n104 4.5005
R51695 VINP.n288 VINP.n104 4.5005
R51696 VINP.n271 VINP.n104 4.5005
R51697 VINP.n290 VINP.n104 4.5005
R51698 VINP.n270 VINP.n104 4.5005
R51699 VINP.n292 VINP.n104 4.5005
R51700 VINP.n269 VINP.n104 4.5005
R51701 VINP.n294 VINP.n104 4.5005
R51702 VINP.n268 VINP.n104 4.5005
R51703 VINP.n296 VINP.n104 4.5005
R51704 VINP.n267 VINP.n104 4.5005
R51705 VINP.n298 VINP.n104 4.5005
R51706 VINP.n266 VINP.n104 4.5005
R51707 VINP.n300 VINP.n104 4.5005
R51708 VINP.n265 VINP.n104 4.5005
R51709 VINP.n302 VINP.n104 4.5005
R51710 VINP.n264 VINP.n104 4.5005
R51711 VINP.n304 VINP.n104 4.5005
R51712 VINP.n263 VINP.n104 4.5005
R51713 VINP.n306 VINP.n104 4.5005
R51714 VINP.n262 VINP.n104 4.5005
R51715 VINP.n308 VINP.n104 4.5005
R51716 VINP.n261 VINP.n104 4.5005
R51717 VINP.n310 VINP.n104 4.5005
R51718 VINP.n260 VINP.n104 4.5005
R51719 VINP.n312 VINP.n104 4.5005
R51720 VINP.n259 VINP.n104 4.5005
R51721 VINP.n314 VINP.n104 4.5005
R51722 VINP.n258 VINP.n104 4.5005
R51723 VINP.n316 VINP.n104 4.5005
R51724 VINP.n257 VINP.n104 4.5005
R51725 VINP.n318 VINP.n104 4.5005
R51726 VINP.n256 VINP.n104 4.5005
R51727 VINP.n320 VINP.n104 4.5005
R51728 VINP.n255 VINP.n104 4.5005
R51729 VINP.n322 VINP.n104 4.5005
R51730 VINP.n254 VINP.n104 4.5005
R51731 VINP.n324 VINP.n104 4.5005
R51732 VINP.n253 VINP.n104 4.5005
R51733 VINP.n326 VINP.n104 4.5005
R51734 VINP.n252 VINP.n104 4.5005
R51735 VINP.n328 VINP.n104 4.5005
R51736 VINP.n251 VINP.n104 4.5005
R51737 VINP.n330 VINP.n104 4.5005
R51738 VINP.n250 VINP.n104 4.5005
R51739 VINP.n332 VINP.n104 4.5005
R51740 VINP.n249 VINP.n104 4.5005
R51741 VINP.n334 VINP.n104 4.5005
R51742 VINP.n248 VINP.n104 4.5005
R51743 VINP.n336 VINP.n104 4.5005
R51744 VINP.n247 VINP.n104 4.5005
R51745 VINP.n338 VINP.n104 4.5005
R51746 VINP.n246 VINP.n104 4.5005
R51747 VINP.n340 VINP.n104 4.5005
R51748 VINP.n245 VINP.n104 4.5005
R51749 VINP.n342 VINP.n104 4.5005
R51750 VINP.n244 VINP.n104 4.5005
R51751 VINP.n344 VINP.n104 4.5005
R51752 VINP.n243 VINP.n104 4.5005
R51753 VINP.n346 VINP.n104 4.5005
R51754 VINP.n242 VINP.n104 4.5005
R51755 VINP.n348 VINP.n104 4.5005
R51756 VINP.n241 VINP.n104 4.5005
R51757 VINP.n350 VINP.n104 4.5005
R51758 VINP.n240 VINP.n104 4.5005
R51759 VINP.n352 VINP.n104 4.5005
R51760 VINP.n239 VINP.n104 4.5005
R51761 VINP.n354 VINP.n104 4.5005
R51762 VINP.n238 VINP.n104 4.5005
R51763 VINP.n356 VINP.n104 4.5005
R51764 VINP.n237 VINP.n104 4.5005
R51765 VINP.n358 VINP.n104 4.5005
R51766 VINP.n236 VINP.n104 4.5005
R51767 VINP.n360 VINP.n104 4.5005
R51768 VINP.n235 VINP.n104 4.5005
R51769 VINP.n362 VINP.n104 4.5005
R51770 VINP.n234 VINP.n104 4.5005
R51771 VINP.n364 VINP.n104 4.5005
R51772 VINP.n233 VINP.n104 4.5005
R51773 VINP.n366 VINP.n104 4.5005
R51774 VINP.n232 VINP.n104 4.5005
R51775 VINP.n368 VINP.n104 4.5005
R51776 VINP.n231 VINP.n104 4.5005
R51777 VINP.n370 VINP.n104 4.5005
R51778 VINP.n230 VINP.n104 4.5005
R51779 VINP.n372 VINP.n104 4.5005
R51780 VINP.n229 VINP.n104 4.5005
R51781 VINP.n374 VINP.n104 4.5005
R51782 VINP.n228 VINP.n104 4.5005
R51783 VINP.n376 VINP.n104 4.5005
R51784 VINP.n227 VINP.n104 4.5005
R51785 VINP.n378 VINP.n104 4.5005
R51786 VINP.n226 VINP.n104 4.5005
R51787 VINP.n380 VINP.n104 4.5005
R51788 VINP.n225 VINP.n104 4.5005
R51789 VINP.n382 VINP.n104 4.5005
R51790 VINP.n224 VINP.n104 4.5005
R51791 VINP.n384 VINP.n104 4.5005
R51792 VINP.n223 VINP.n104 4.5005
R51793 VINP.n386 VINP.n104 4.5005
R51794 VINP.n222 VINP.n104 4.5005
R51795 VINP.n388 VINP.n104 4.5005
R51796 VINP.n221 VINP.n104 4.5005
R51797 VINP.n390 VINP.n104 4.5005
R51798 VINP.n220 VINP.n104 4.5005
R51799 VINP.n392 VINP.n104 4.5005
R51800 VINP.n219 VINP.n104 4.5005
R51801 VINP.n394 VINP.n104 4.5005
R51802 VINP.n218 VINP.n104 4.5005
R51803 VINP.n396 VINP.n104 4.5005
R51804 VINP.n217 VINP.n104 4.5005
R51805 VINP.n398 VINP.n104 4.5005
R51806 VINP.n216 VINP.n104 4.5005
R51807 VINP.n400 VINP.n104 4.5005
R51808 VINP.n215 VINP.n104 4.5005
R51809 VINP.n654 VINP.n104 4.5005
R51810 VINP.n656 VINP.n104 4.5005
R51811 VINP.n104 VINP.n0 4.5005
R51812 VINP.n278 VINP.n197 4.5005
R51813 VINP.n276 VINP.n197 4.5005
R51814 VINP.n280 VINP.n197 4.5005
R51815 VINP.n275 VINP.n197 4.5005
R51816 VINP.n282 VINP.n197 4.5005
R51817 VINP.n274 VINP.n197 4.5005
R51818 VINP.n284 VINP.n197 4.5005
R51819 VINP.n273 VINP.n197 4.5005
R51820 VINP.n286 VINP.n197 4.5005
R51821 VINP.n272 VINP.n197 4.5005
R51822 VINP.n288 VINP.n197 4.5005
R51823 VINP.n271 VINP.n197 4.5005
R51824 VINP.n290 VINP.n197 4.5005
R51825 VINP.n270 VINP.n197 4.5005
R51826 VINP.n292 VINP.n197 4.5005
R51827 VINP.n269 VINP.n197 4.5005
R51828 VINP.n294 VINP.n197 4.5005
R51829 VINP.n268 VINP.n197 4.5005
R51830 VINP.n296 VINP.n197 4.5005
R51831 VINP.n267 VINP.n197 4.5005
R51832 VINP.n298 VINP.n197 4.5005
R51833 VINP.n266 VINP.n197 4.5005
R51834 VINP.n300 VINP.n197 4.5005
R51835 VINP.n265 VINP.n197 4.5005
R51836 VINP.n302 VINP.n197 4.5005
R51837 VINP.n264 VINP.n197 4.5005
R51838 VINP.n304 VINP.n197 4.5005
R51839 VINP.n263 VINP.n197 4.5005
R51840 VINP.n306 VINP.n197 4.5005
R51841 VINP.n262 VINP.n197 4.5005
R51842 VINP.n308 VINP.n197 4.5005
R51843 VINP.n261 VINP.n197 4.5005
R51844 VINP.n310 VINP.n197 4.5005
R51845 VINP.n260 VINP.n197 4.5005
R51846 VINP.n312 VINP.n197 4.5005
R51847 VINP.n259 VINP.n197 4.5005
R51848 VINP.n314 VINP.n197 4.5005
R51849 VINP.n258 VINP.n197 4.5005
R51850 VINP.n316 VINP.n197 4.5005
R51851 VINP.n257 VINP.n197 4.5005
R51852 VINP.n318 VINP.n197 4.5005
R51853 VINP.n256 VINP.n197 4.5005
R51854 VINP.n320 VINP.n197 4.5005
R51855 VINP.n255 VINP.n197 4.5005
R51856 VINP.n322 VINP.n197 4.5005
R51857 VINP.n254 VINP.n197 4.5005
R51858 VINP.n324 VINP.n197 4.5005
R51859 VINP.n253 VINP.n197 4.5005
R51860 VINP.n326 VINP.n197 4.5005
R51861 VINP.n252 VINP.n197 4.5005
R51862 VINP.n328 VINP.n197 4.5005
R51863 VINP.n251 VINP.n197 4.5005
R51864 VINP.n330 VINP.n197 4.5005
R51865 VINP.n250 VINP.n197 4.5005
R51866 VINP.n332 VINP.n197 4.5005
R51867 VINP.n249 VINP.n197 4.5005
R51868 VINP.n334 VINP.n197 4.5005
R51869 VINP.n248 VINP.n197 4.5005
R51870 VINP.n336 VINP.n197 4.5005
R51871 VINP.n247 VINP.n197 4.5005
R51872 VINP.n338 VINP.n197 4.5005
R51873 VINP.n246 VINP.n197 4.5005
R51874 VINP.n340 VINP.n197 4.5005
R51875 VINP.n245 VINP.n197 4.5005
R51876 VINP.n342 VINP.n197 4.5005
R51877 VINP.n244 VINP.n197 4.5005
R51878 VINP.n344 VINP.n197 4.5005
R51879 VINP.n243 VINP.n197 4.5005
R51880 VINP.n346 VINP.n197 4.5005
R51881 VINP.n242 VINP.n197 4.5005
R51882 VINP.n348 VINP.n197 4.5005
R51883 VINP.n241 VINP.n197 4.5005
R51884 VINP.n350 VINP.n197 4.5005
R51885 VINP.n240 VINP.n197 4.5005
R51886 VINP.n352 VINP.n197 4.5005
R51887 VINP.n239 VINP.n197 4.5005
R51888 VINP.n354 VINP.n197 4.5005
R51889 VINP.n238 VINP.n197 4.5005
R51890 VINP.n356 VINP.n197 4.5005
R51891 VINP.n237 VINP.n197 4.5005
R51892 VINP.n358 VINP.n197 4.5005
R51893 VINP.n236 VINP.n197 4.5005
R51894 VINP.n360 VINP.n197 4.5005
R51895 VINP.n235 VINP.n197 4.5005
R51896 VINP.n362 VINP.n197 4.5005
R51897 VINP.n234 VINP.n197 4.5005
R51898 VINP.n364 VINP.n197 4.5005
R51899 VINP.n233 VINP.n197 4.5005
R51900 VINP.n366 VINP.n197 4.5005
R51901 VINP.n232 VINP.n197 4.5005
R51902 VINP.n368 VINP.n197 4.5005
R51903 VINP.n231 VINP.n197 4.5005
R51904 VINP.n370 VINP.n197 4.5005
R51905 VINP.n230 VINP.n197 4.5005
R51906 VINP.n372 VINP.n197 4.5005
R51907 VINP.n229 VINP.n197 4.5005
R51908 VINP.n374 VINP.n197 4.5005
R51909 VINP.n228 VINP.n197 4.5005
R51910 VINP.n376 VINP.n197 4.5005
R51911 VINP.n227 VINP.n197 4.5005
R51912 VINP.n378 VINP.n197 4.5005
R51913 VINP.n226 VINP.n197 4.5005
R51914 VINP.n380 VINP.n197 4.5005
R51915 VINP.n225 VINP.n197 4.5005
R51916 VINP.n382 VINP.n197 4.5005
R51917 VINP.n224 VINP.n197 4.5005
R51918 VINP.n384 VINP.n197 4.5005
R51919 VINP.n223 VINP.n197 4.5005
R51920 VINP.n386 VINP.n197 4.5005
R51921 VINP.n222 VINP.n197 4.5005
R51922 VINP.n388 VINP.n197 4.5005
R51923 VINP.n221 VINP.n197 4.5005
R51924 VINP.n390 VINP.n197 4.5005
R51925 VINP.n220 VINP.n197 4.5005
R51926 VINP.n392 VINP.n197 4.5005
R51927 VINP.n219 VINP.n197 4.5005
R51928 VINP.n394 VINP.n197 4.5005
R51929 VINP.n218 VINP.n197 4.5005
R51930 VINP.n396 VINP.n197 4.5005
R51931 VINP.n217 VINP.n197 4.5005
R51932 VINP.n398 VINP.n197 4.5005
R51933 VINP.n216 VINP.n197 4.5005
R51934 VINP.n400 VINP.n197 4.5005
R51935 VINP.n215 VINP.n197 4.5005
R51936 VINP.n654 VINP.n197 4.5005
R51937 VINP.n656 VINP.n197 4.5005
R51938 VINP.n197 VINP.n0 4.5005
R51939 VINP.n278 VINP.n103 4.5005
R51940 VINP.n276 VINP.n103 4.5005
R51941 VINP.n280 VINP.n103 4.5005
R51942 VINP.n275 VINP.n103 4.5005
R51943 VINP.n282 VINP.n103 4.5005
R51944 VINP.n274 VINP.n103 4.5005
R51945 VINP.n284 VINP.n103 4.5005
R51946 VINP.n273 VINP.n103 4.5005
R51947 VINP.n286 VINP.n103 4.5005
R51948 VINP.n272 VINP.n103 4.5005
R51949 VINP.n288 VINP.n103 4.5005
R51950 VINP.n271 VINP.n103 4.5005
R51951 VINP.n290 VINP.n103 4.5005
R51952 VINP.n270 VINP.n103 4.5005
R51953 VINP.n292 VINP.n103 4.5005
R51954 VINP.n269 VINP.n103 4.5005
R51955 VINP.n294 VINP.n103 4.5005
R51956 VINP.n268 VINP.n103 4.5005
R51957 VINP.n296 VINP.n103 4.5005
R51958 VINP.n267 VINP.n103 4.5005
R51959 VINP.n298 VINP.n103 4.5005
R51960 VINP.n266 VINP.n103 4.5005
R51961 VINP.n300 VINP.n103 4.5005
R51962 VINP.n265 VINP.n103 4.5005
R51963 VINP.n302 VINP.n103 4.5005
R51964 VINP.n264 VINP.n103 4.5005
R51965 VINP.n304 VINP.n103 4.5005
R51966 VINP.n263 VINP.n103 4.5005
R51967 VINP.n306 VINP.n103 4.5005
R51968 VINP.n262 VINP.n103 4.5005
R51969 VINP.n308 VINP.n103 4.5005
R51970 VINP.n261 VINP.n103 4.5005
R51971 VINP.n310 VINP.n103 4.5005
R51972 VINP.n260 VINP.n103 4.5005
R51973 VINP.n312 VINP.n103 4.5005
R51974 VINP.n259 VINP.n103 4.5005
R51975 VINP.n314 VINP.n103 4.5005
R51976 VINP.n258 VINP.n103 4.5005
R51977 VINP.n316 VINP.n103 4.5005
R51978 VINP.n257 VINP.n103 4.5005
R51979 VINP.n318 VINP.n103 4.5005
R51980 VINP.n256 VINP.n103 4.5005
R51981 VINP.n320 VINP.n103 4.5005
R51982 VINP.n255 VINP.n103 4.5005
R51983 VINP.n322 VINP.n103 4.5005
R51984 VINP.n254 VINP.n103 4.5005
R51985 VINP.n324 VINP.n103 4.5005
R51986 VINP.n253 VINP.n103 4.5005
R51987 VINP.n326 VINP.n103 4.5005
R51988 VINP.n252 VINP.n103 4.5005
R51989 VINP.n328 VINP.n103 4.5005
R51990 VINP.n251 VINP.n103 4.5005
R51991 VINP.n330 VINP.n103 4.5005
R51992 VINP.n250 VINP.n103 4.5005
R51993 VINP.n332 VINP.n103 4.5005
R51994 VINP.n249 VINP.n103 4.5005
R51995 VINP.n334 VINP.n103 4.5005
R51996 VINP.n248 VINP.n103 4.5005
R51997 VINP.n336 VINP.n103 4.5005
R51998 VINP.n247 VINP.n103 4.5005
R51999 VINP.n338 VINP.n103 4.5005
R52000 VINP.n246 VINP.n103 4.5005
R52001 VINP.n340 VINP.n103 4.5005
R52002 VINP.n245 VINP.n103 4.5005
R52003 VINP.n342 VINP.n103 4.5005
R52004 VINP.n244 VINP.n103 4.5005
R52005 VINP.n344 VINP.n103 4.5005
R52006 VINP.n243 VINP.n103 4.5005
R52007 VINP.n346 VINP.n103 4.5005
R52008 VINP.n242 VINP.n103 4.5005
R52009 VINP.n348 VINP.n103 4.5005
R52010 VINP.n241 VINP.n103 4.5005
R52011 VINP.n350 VINP.n103 4.5005
R52012 VINP.n240 VINP.n103 4.5005
R52013 VINP.n352 VINP.n103 4.5005
R52014 VINP.n239 VINP.n103 4.5005
R52015 VINP.n354 VINP.n103 4.5005
R52016 VINP.n238 VINP.n103 4.5005
R52017 VINP.n356 VINP.n103 4.5005
R52018 VINP.n237 VINP.n103 4.5005
R52019 VINP.n358 VINP.n103 4.5005
R52020 VINP.n236 VINP.n103 4.5005
R52021 VINP.n360 VINP.n103 4.5005
R52022 VINP.n235 VINP.n103 4.5005
R52023 VINP.n362 VINP.n103 4.5005
R52024 VINP.n234 VINP.n103 4.5005
R52025 VINP.n364 VINP.n103 4.5005
R52026 VINP.n233 VINP.n103 4.5005
R52027 VINP.n366 VINP.n103 4.5005
R52028 VINP.n232 VINP.n103 4.5005
R52029 VINP.n368 VINP.n103 4.5005
R52030 VINP.n231 VINP.n103 4.5005
R52031 VINP.n370 VINP.n103 4.5005
R52032 VINP.n230 VINP.n103 4.5005
R52033 VINP.n372 VINP.n103 4.5005
R52034 VINP.n229 VINP.n103 4.5005
R52035 VINP.n374 VINP.n103 4.5005
R52036 VINP.n228 VINP.n103 4.5005
R52037 VINP.n376 VINP.n103 4.5005
R52038 VINP.n227 VINP.n103 4.5005
R52039 VINP.n378 VINP.n103 4.5005
R52040 VINP.n226 VINP.n103 4.5005
R52041 VINP.n380 VINP.n103 4.5005
R52042 VINP.n225 VINP.n103 4.5005
R52043 VINP.n382 VINP.n103 4.5005
R52044 VINP.n224 VINP.n103 4.5005
R52045 VINP.n384 VINP.n103 4.5005
R52046 VINP.n223 VINP.n103 4.5005
R52047 VINP.n386 VINP.n103 4.5005
R52048 VINP.n222 VINP.n103 4.5005
R52049 VINP.n388 VINP.n103 4.5005
R52050 VINP.n221 VINP.n103 4.5005
R52051 VINP.n390 VINP.n103 4.5005
R52052 VINP.n220 VINP.n103 4.5005
R52053 VINP.n392 VINP.n103 4.5005
R52054 VINP.n219 VINP.n103 4.5005
R52055 VINP.n394 VINP.n103 4.5005
R52056 VINP.n218 VINP.n103 4.5005
R52057 VINP.n396 VINP.n103 4.5005
R52058 VINP.n217 VINP.n103 4.5005
R52059 VINP.n398 VINP.n103 4.5005
R52060 VINP.n216 VINP.n103 4.5005
R52061 VINP.n400 VINP.n103 4.5005
R52062 VINP.n215 VINP.n103 4.5005
R52063 VINP.n654 VINP.n103 4.5005
R52064 VINP.n656 VINP.n103 4.5005
R52065 VINP.n103 VINP.n0 4.5005
R52066 VINP.n278 VINP.n198 4.5005
R52067 VINP.n276 VINP.n198 4.5005
R52068 VINP.n280 VINP.n198 4.5005
R52069 VINP.n275 VINP.n198 4.5005
R52070 VINP.n282 VINP.n198 4.5005
R52071 VINP.n274 VINP.n198 4.5005
R52072 VINP.n284 VINP.n198 4.5005
R52073 VINP.n273 VINP.n198 4.5005
R52074 VINP.n286 VINP.n198 4.5005
R52075 VINP.n272 VINP.n198 4.5005
R52076 VINP.n288 VINP.n198 4.5005
R52077 VINP.n271 VINP.n198 4.5005
R52078 VINP.n290 VINP.n198 4.5005
R52079 VINP.n270 VINP.n198 4.5005
R52080 VINP.n292 VINP.n198 4.5005
R52081 VINP.n269 VINP.n198 4.5005
R52082 VINP.n294 VINP.n198 4.5005
R52083 VINP.n268 VINP.n198 4.5005
R52084 VINP.n296 VINP.n198 4.5005
R52085 VINP.n267 VINP.n198 4.5005
R52086 VINP.n298 VINP.n198 4.5005
R52087 VINP.n266 VINP.n198 4.5005
R52088 VINP.n300 VINP.n198 4.5005
R52089 VINP.n265 VINP.n198 4.5005
R52090 VINP.n302 VINP.n198 4.5005
R52091 VINP.n264 VINP.n198 4.5005
R52092 VINP.n304 VINP.n198 4.5005
R52093 VINP.n263 VINP.n198 4.5005
R52094 VINP.n306 VINP.n198 4.5005
R52095 VINP.n262 VINP.n198 4.5005
R52096 VINP.n308 VINP.n198 4.5005
R52097 VINP.n261 VINP.n198 4.5005
R52098 VINP.n310 VINP.n198 4.5005
R52099 VINP.n260 VINP.n198 4.5005
R52100 VINP.n312 VINP.n198 4.5005
R52101 VINP.n259 VINP.n198 4.5005
R52102 VINP.n314 VINP.n198 4.5005
R52103 VINP.n258 VINP.n198 4.5005
R52104 VINP.n316 VINP.n198 4.5005
R52105 VINP.n257 VINP.n198 4.5005
R52106 VINP.n318 VINP.n198 4.5005
R52107 VINP.n256 VINP.n198 4.5005
R52108 VINP.n320 VINP.n198 4.5005
R52109 VINP.n255 VINP.n198 4.5005
R52110 VINP.n322 VINP.n198 4.5005
R52111 VINP.n254 VINP.n198 4.5005
R52112 VINP.n324 VINP.n198 4.5005
R52113 VINP.n253 VINP.n198 4.5005
R52114 VINP.n326 VINP.n198 4.5005
R52115 VINP.n252 VINP.n198 4.5005
R52116 VINP.n328 VINP.n198 4.5005
R52117 VINP.n251 VINP.n198 4.5005
R52118 VINP.n330 VINP.n198 4.5005
R52119 VINP.n250 VINP.n198 4.5005
R52120 VINP.n332 VINP.n198 4.5005
R52121 VINP.n249 VINP.n198 4.5005
R52122 VINP.n334 VINP.n198 4.5005
R52123 VINP.n248 VINP.n198 4.5005
R52124 VINP.n336 VINP.n198 4.5005
R52125 VINP.n247 VINP.n198 4.5005
R52126 VINP.n338 VINP.n198 4.5005
R52127 VINP.n246 VINP.n198 4.5005
R52128 VINP.n340 VINP.n198 4.5005
R52129 VINP.n245 VINP.n198 4.5005
R52130 VINP.n342 VINP.n198 4.5005
R52131 VINP.n244 VINP.n198 4.5005
R52132 VINP.n344 VINP.n198 4.5005
R52133 VINP.n243 VINP.n198 4.5005
R52134 VINP.n346 VINP.n198 4.5005
R52135 VINP.n242 VINP.n198 4.5005
R52136 VINP.n348 VINP.n198 4.5005
R52137 VINP.n241 VINP.n198 4.5005
R52138 VINP.n350 VINP.n198 4.5005
R52139 VINP.n240 VINP.n198 4.5005
R52140 VINP.n352 VINP.n198 4.5005
R52141 VINP.n239 VINP.n198 4.5005
R52142 VINP.n354 VINP.n198 4.5005
R52143 VINP.n238 VINP.n198 4.5005
R52144 VINP.n356 VINP.n198 4.5005
R52145 VINP.n237 VINP.n198 4.5005
R52146 VINP.n358 VINP.n198 4.5005
R52147 VINP.n236 VINP.n198 4.5005
R52148 VINP.n360 VINP.n198 4.5005
R52149 VINP.n235 VINP.n198 4.5005
R52150 VINP.n362 VINP.n198 4.5005
R52151 VINP.n234 VINP.n198 4.5005
R52152 VINP.n364 VINP.n198 4.5005
R52153 VINP.n233 VINP.n198 4.5005
R52154 VINP.n366 VINP.n198 4.5005
R52155 VINP.n232 VINP.n198 4.5005
R52156 VINP.n368 VINP.n198 4.5005
R52157 VINP.n231 VINP.n198 4.5005
R52158 VINP.n370 VINP.n198 4.5005
R52159 VINP.n230 VINP.n198 4.5005
R52160 VINP.n372 VINP.n198 4.5005
R52161 VINP.n229 VINP.n198 4.5005
R52162 VINP.n374 VINP.n198 4.5005
R52163 VINP.n228 VINP.n198 4.5005
R52164 VINP.n376 VINP.n198 4.5005
R52165 VINP.n227 VINP.n198 4.5005
R52166 VINP.n378 VINP.n198 4.5005
R52167 VINP.n226 VINP.n198 4.5005
R52168 VINP.n380 VINP.n198 4.5005
R52169 VINP.n225 VINP.n198 4.5005
R52170 VINP.n382 VINP.n198 4.5005
R52171 VINP.n224 VINP.n198 4.5005
R52172 VINP.n384 VINP.n198 4.5005
R52173 VINP.n223 VINP.n198 4.5005
R52174 VINP.n386 VINP.n198 4.5005
R52175 VINP.n222 VINP.n198 4.5005
R52176 VINP.n388 VINP.n198 4.5005
R52177 VINP.n221 VINP.n198 4.5005
R52178 VINP.n390 VINP.n198 4.5005
R52179 VINP.n220 VINP.n198 4.5005
R52180 VINP.n392 VINP.n198 4.5005
R52181 VINP.n219 VINP.n198 4.5005
R52182 VINP.n394 VINP.n198 4.5005
R52183 VINP.n218 VINP.n198 4.5005
R52184 VINP.n396 VINP.n198 4.5005
R52185 VINP.n217 VINP.n198 4.5005
R52186 VINP.n398 VINP.n198 4.5005
R52187 VINP.n216 VINP.n198 4.5005
R52188 VINP.n400 VINP.n198 4.5005
R52189 VINP.n215 VINP.n198 4.5005
R52190 VINP.n654 VINP.n198 4.5005
R52191 VINP.n656 VINP.n198 4.5005
R52192 VINP.n198 VINP.n0 4.5005
R52193 VINP.n278 VINP.n102 4.5005
R52194 VINP.n276 VINP.n102 4.5005
R52195 VINP.n280 VINP.n102 4.5005
R52196 VINP.n275 VINP.n102 4.5005
R52197 VINP.n282 VINP.n102 4.5005
R52198 VINP.n274 VINP.n102 4.5005
R52199 VINP.n284 VINP.n102 4.5005
R52200 VINP.n273 VINP.n102 4.5005
R52201 VINP.n286 VINP.n102 4.5005
R52202 VINP.n272 VINP.n102 4.5005
R52203 VINP.n288 VINP.n102 4.5005
R52204 VINP.n271 VINP.n102 4.5005
R52205 VINP.n290 VINP.n102 4.5005
R52206 VINP.n270 VINP.n102 4.5005
R52207 VINP.n292 VINP.n102 4.5005
R52208 VINP.n269 VINP.n102 4.5005
R52209 VINP.n294 VINP.n102 4.5005
R52210 VINP.n268 VINP.n102 4.5005
R52211 VINP.n296 VINP.n102 4.5005
R52212 VINP.n267 VINP.n102 4.5005
R52213 VINP.n298 VINP.n102 4.5005
R52214 VINP.n266 VINP.n102 4.5005
R52215 VINP.n300 VINP.n102 4.5005
R52216 VINP.n265 VINP.n102 4.5005
R52217 VINP.n302 VINP.n102 4.5005
R52218 VINP.n264 VINP.n102 4.5005
R52219 VINP.n304 VINP.n102 4.5005
R52220 VINP.n263 VINP.n102 4.5005
R52221 VINP.n306 VINP.n102 4.5005
R52222 VINP.n262 VINP.n102 4.5005
R52223 VINP.n308 VINP.n102 4.5005
R52224 VINP.n261 VINP.n102 4.5005
R52225 VINP.n310 VINP.n102 4.5005
R52226 VINP.n260 VINP.n102 4.5005
R52227 VINP.n312 VINP.n102 4.5005
R52228 VINP.n259 VINP.n102 4.5005
R52229 VINP.n314 VINP.n102 4.5005
R52230 VINP.n258 VINP.n102 4.5005
R52231 VINP.n316 VINP.n102 4.5005
R52232 VINP.n257 VINP.n102 4.5005
R52233 VINP.n318 VINP.n102 4.5005
R52234 VINP.n256 VINP.n102 4.5005
R52235 VINP.n320 VINP.n102 4.5005
R52236 VINP.n255 VINP.n102 4.5005
R52237 VINP.n322 VINP.n102 4.5005
R52238 VINP.n254 VINP.n102 4.5005
R52239 VINP.n324 VINP.n102 4.5005
R52240 VINP.n253 VINP.n102 4.5005
R52241 VINP.n326 VINP.n102 4.5005
R52242 VINP.n252 VINP.n102 4.5005
R52243 VINP.n328 VINP.n102 4.5005
R52244 VINP.n251 VINP.n102 4.5005
R52245 VINP.n330 VINP.n102 4.5005
R52246 VINP.n250 VINP.n102 4.5005
R52247 VINP.n332 VINP.n102 4.5005
R52248 VINP.n249 VINP.n102 4.5005
R52249 VINP.n334 VINP.n102 4.5005
R52250 VINP.n248 VINP.n102 4.5005
R52251 VINP.n336 VINP.n102 4.5005
R52252 VINP.n247 VINP.n102 4.5005
R52253 VINP.n338 VINP.n102 4.5005
R52254 VINP.n246 VINP.n102 4.5005
R52255 VINP.n340 VINP.n102 4.5005
R52256 VINP.n245 VINP.n102 4.5005
R52257 VINP.n342 VINP.n102 4.5005
R52258 VINP.n244 VINP.n102 4.5005
R52259 VINP.n344 VINP.n102 4.5005
R52260 VINP.n243 VINP.n102 4.5005
R52261 VINP.n346 VINP.n102 4.5005
R52262 VINP.n242 VINP.n102 4.5005
R52263 VINP.n348 VINP.n102 4.5005
R52264 VINP.n241 VINP.n102 4.5005
R52265 VINP.n350 VINP.n102 4.5005
R52266 VINP.n240 VINP.n102 4.5005
R52267 VINP.n352 VINP.n102 4.5005
R52268 VINP.n239 VINP.n102 4.5005
R52269 VINP.n354 VINP.n102 4.5005
R52270 VINP.n238 VINP.n102 4.5005
R52271 VINP.n356 VINP.n102 4.5005
R52272 VINP.n237 VINP.n102 4.5005
R52273 VINP.n358 VINP.n102 4.5005
R52274 VINP.n236 VINP.n102 4.5005
R52275 VINP.n360 VINP.n102 4.5005
R52276 VINP.n235 VINP.n102 4.5005
R52277 VINP.n362 VINP.n102 4.5005
R52278 VINP.n234 VINP.n102 4.5005
R52279 VINP.n364 VINP.n102 4.5005
R52280 VINP.n233 VINP.n102 4.5005
R52281 VINP.n366 VINP.n102 4.5005
R52282 VINP.n232 VINP.n102 4.5005
R52283 VINP.n368 VINP.n102 4.5005
R52284 VINP.n231 VINP.n102 4.5005
R52285 VINP.n370 VINP.n102 4.5005
R52286 VINP.n230 VINP.n102 4.5005
R52287 VINP.n372 VINP.n102 4.5005
R52288 VINP.n229 VINP.n102 4.5005
R52289 VINP.n374 VINP.n102 4.5005
R52290 VINP.n228 VINP.n102 4.5005
R52291 VINP.n376 VINP.n102 4.5005
R52292 VINP.n227 VINP.n102 4.5005
R52293 VINP.n378 VINP.n102 4.5005
R52294 VINP.n226 VINP.n102 4.5005
R52295 VINP.n380 VINP.n102 4.5005
R52296 VINP.n225 VINP.n102 4.5005
R52297 VINP.n382 VINP.n102 4.5005
R52298 VINP.n224 VINP.n102 4.5005
R52299 VINP.n384 VINP.n102 4.5005
R52300 VINP.n223 VINP.n102 4.5005
R52301 VINP.n386 VINP.n102 4.5005
R52302 VINP.n222 VINP.n102 4.5005
R52303 VINP.n388 VINP.n102 4.5005
R52304 VINP.n221 VINP.n102 4.5005
R52305 VINP.n390 VINP.n102 4.5005
R52306 VINP.n220 VINP.n102 4.5005
R52307 VINP.n392 VINP.n102 4.5005
R52308 VINP.n219 VINP.n102 4.5005
R52309 VINP.n394 VINP.n102 4.5005
R52310 VINP.n218 VINP.n102 4.5005
R52311 VINP.n396 VINP.n102 4.5005
R52312 VINP.n217 VINP.n102 4.5005
R52313 VINP.n398 VINP.n102 4.5005
R52314 VINP.n216 VINP.n102 4.5005
R52315 VINP.n400 VINP.n102 4.5005
R52316 VINP.n215 VINP.n102 4.5005
R52317 VINP.n654 VINP.n102 4.5005
R52318 VINP.n656 VINP.n102 4.5005
R52319 VINP.n102 VINP.n0 4.5005
R52320 VINP.n278 VINP.n199 4.5005
R52321 VINP.n276 VINP.n199 4.5005
R52322 VINP.n280 VINP.n199 4.5005
R52323 VINP.n275 VINP.n199 4.5005
R52324 VINP.n282 VINP.n199 4.5005
R52325 VINP.n274 VINP.n199 4.5005
R52326 VINP.n284 VINP.n199 4.5005
R52327 VINP.n273 VINP.n199 4.5005
R52328 VINP.n286 VINP.n199 4.5005
R52329 VINP.n272 VINP.n199 4.5005
R52330 VINP.n288 VINP.n199 4.5005
R52331 VINP.n271 VINP.n199 4.5005
R52332 VINP.n290 VINP.n199 4.5005
R52333 VINP.n270 VINP.n199 4.5005
R52334 VINP.n292 VINP.n199 4.5005
R52335 VINP.n269 VINP.n199 4.5005
R52336 VINP.n294 VINP.n199 4.5005
R52337 VINP.n268 VINP.n199 4.5005
R52338 VINP.n296 VINP.n199 4.5005
R52339 VINP.n267 VINP.n199 4.5005
R52340 VINP.n298 VINP.n199 4.5005
R52341 VINP.n266 VINP.n199 4.5005
R52342 VINP.n300 VINP.n199 4.5005
R52343 VINP.n265 VINP.n199 4.5005
R52344 VINP.n302 VINP.n199 4.5005
R52345 VINP.n264 VINP.n199 4.5005
R52346 VINP.n304 VINP.n199 4.5005
R52347 VINP.n263 VINP.n199 4.5005
R52348 VINP.n306 VINP.n199 4.5005
R52349 VINP.n262 VINP.n199 4.5005
R52350 VINP.n308 VINP.n199 4.5005
R52351 VINP.n261 VINP.n199 4.5005
R52352 VINP.n310 VINP.n199 4.5005
R52353 VINP.n260 VINP.n199 4.5005
R52354 VINP.n312 VINP.n199 4.5005
R52355 VINP.n259 VINP.n199 4.5005
R52356 VINP.n314 VINP.n199 4.5005
R52357 VINP.n258 VINP.n199 4.5005
R52358 VINP.n316 VINP.n199 4.5005
R52359 VINP.n257 VINP.n199 4.5005
R52360 VINP.n318 VINP.n199 4.5005
R52361 VINP.n256 VINP.n199 4.5005
R52362 VINP.n320 VINP.n199 4.5005
R52363 VINP.n255 VINP.n199 4.5005
R52364 VINP.n322 VINP.n199 4.5005
R52365 VINP.n254 VINP.n199 4.5005
R52366 VINP.n324 VINP.n199 4.5005
R52367 VINP.n253 VINP.n199 4.5005
R52368 VINP.n326 VINP.n199 4.5005
R52369 VINP.n252 VINP.n199 4.5005
R52370 VINP.n328 VINP.n199 4.5005
R52371 VINP.n251 VINP.n199 4.5005
R52372 VINP.n330 VINP.n199 4.5005
R52373 VINP.n250 VINP.n199 4.5005
R52374 VINP.n332 VINP.n199 4.5005
R52375 VINP.n249 VINP.n199 4.5005
R52376 VINP.n334 VINP.n199 4.5005
R52377 VINP.n248 VINP.n199 4.5005
R52378 VINP.n336 VINP.n199 4.5005
R52379 VINP.n247 VINP.n199 4.5005
R52380 VINP.n338 VINP.n199 4.5005
R52381 VINP.n246 VINP.n199 4.5005
R52382 VINP.n340 VINP.n199 4.5005
R52383 VINP.n245 VINP.n199 4.5005
R52384 VINP.n342 VINP.n199 4.5005
R52385 VINP.n244 VINP.n199 4.5005
R52386 VINP.n344 VINP.n199 4.5005
R52387 VINP.n243 VINP.n199 4.5005
R52388 VINP.n346 VINP.n199 4.5005
R52389 VINP.n242 VINP.n199 4.5005
R52390 VINP.n348 VINP.n199 4.5005
R52391 VINP.n241 VINP.n199 4.5005
R52392 VINP.n350 VINP.n199 4.5005
R52393 VINP.n240 VINP.n199 4.5005
R52394 VINP.n352 VINP.n199 4.5005
R52395 VINP.n239 VINP.n199 4.5005
R52396 VINP.n354 VINP.n199 4.5005
R52397 VINP.n238 VINP.n199 4.5005
R52398 VINP.n356 VINP.n199 4.5005
R52399 VINP.n237 VINP.n199 4.5005
R52400 VINP.n358 VINP.n199 4.5005
R52401 VINP.n236 VINP.n199 4.5005
R52402 VINP.n360 VINP.n199 4.5005
R52403 VINP.n235 VINP.n199 4.5005
R52404 VINP.n362 VINP.n199 4.5005
R52405 VINP.n234 VINP.n199 4.5005
R52406 VINP.n364 VINP.n199 4.5005
R52407 VINP.n233 VINP.n199 4.5005
R52408 VINP.n366 VINP.n199 4.5005
R52409 VINP.n232 VINP.n199 4.5005
R52410 VINP.n368 VINP.n199 4.5005
R52411 VINP.n231 VINP.n199 4.5005
R52412 VINP.n370 VINP.n199 4.5005
R52413 VINP.n230 VINP.n199 4.5005
R52414 VINP.n372 VINP.n199 4.5005
R52415 VINP.n229 VINP.n199 4.5005
R52416 VINP.n374 VINP.n199 4.5005
R52417 VINP.n228 VINP.n199 4.5005
R52418 VINP.n376 VINP.n199 4.5005
R52419 VINP.n227 VINP.n199 4.5005
R52420 VINP.n378 VINP.n199 4.5005
R52421 VINP.n226 VINP.n199 4.5005
R52422 VINP.n380 VINP.n199 4.5005
R52423 VINP.n225 VINP.n199 4.5005
R52424 VINP.n382 VINP.n199 4.5005
R52425 VINP.n224 VINP.n199 4.5005
R52426 VINP.n384 VINP.n199 4.5005
R52427 VINP.n223 VINP.n199 4.5005
R52428 VINP.n386 VINP.n199 4.5005
R52429 VINP.n222 VINP.n199 4.5005
R52430 VINP.n388 VINP.n199 4.5005
R52431 VINP.n221 VINP.n199 4.5005
R52432 VINP.n390 VINP.n199 4.5005
R52433 VINP.n220 VINP.n199 4.5005
R52434 VINP.n392 VINP.n199 4.5005
R52435 VINP.n219 VINP.n199 4.5005
R52436 VINP.n394 VINP.n199 4.5005
R52437 VINP.n218 VINP.n199 4.5005
R52438 VINP.n396 VINP.n199 4.5005
R52439 VINP.n217 VINP.n199 4.5005
R52440 VINP.n398 VINP.n199 4.5005
R52441 VINP.n216 VINP.n199 4.5005
R52442 VINP.n400 VINP.n199 4.5005
R52443 VINP.n215 VINP.n199 4.5005
R52444 VINP.n654 VINP.n199 4.5005
R52445 VINP.n656 VINP.n199 4.5005
R52446 VINP.n199 VINP.n0 4.5005
R52447 VINP.n278 VINP.n101 4.5005
R52448 VINP.n276 VINP.n101 4.5005
R52449 VINP.n280 VINP.n101 4.5005
R52450 VINP.n275 VINP.n101 4.5005
R52451 VINP.n282 VINP.n101 4.5005
R52452 VINP.n274 VINP.n101 4.5005
R52453 VINP.n284 VINP.n101 4.5005
R52454 VINP.n273 VINP.n101 4.5005
R52455 VINP.n286 VINP.n101 4.5005
R52456 VINP.n272 VINP.n101 4.5005
R52457 VINP.n288 VINP.n101 4.5005
R52458 VINP.n271 VINP.n101 4.5005
R52459 VINP.n290 VINP.n101 4.5005
R52460 VINP.n270 VINP.n101 4.5005
R52461 VINP.n292 VINP.n101 4.5005
R52462 VINP.n269 VINP.n101 4.5005
R52463 VINP.n294 VINP.n101 4.5005
R52464 VINP.n268 VINP.n101 4.5005
R52465 VINP.n296 VINP.n101 4.5005
R52466 VINP.n267 VINP.n101 4.5005
R52467 VINP.n298 VINP.n101 4.5005
R52468 VINP.n266 VINP.n101 4.5005
R52469 VINP.n300 VINP.n101 4.5005
R52470 VINP.n265 VINP.n101 4.5005
R52471 VINP.n302 VINP.n101 4.5005
R52472 VINP.n264 VINP.n101 4.5005
R52473 VINP.n304 VINP.n101 4.5005
R52474 VINP.n263 VINP.n101 4.5005
R52475 VINP.n306 VINP.n101 4.5005
R52476 VINP.n262 VINP.n101 4.5005
R52477 VINP.n308 VINP.n101 4.5005
R52478 VINP.n261 VINP.n101 4.5005
R52479 VINP.n310 VINP.n101 4.5005
R52480 VINP.n260 VINP.n101 4.5005
R52481 VINP.n312 VINP.n101 4.5005
R52482 VINP.n259 VINP.n101 4.5005
R52483 VINP.n314 VINP.n101 4.5005
R52484 VINP.n258 VINP.n101 4.5005
R52485 VINP.n316 VINP.n101 4.5005
R52486 VINP.n257 VINP.n101 4.5005
R52487 VINP.n318 VINP.n101 4.5005
R52488 VINP.n256 VINP.n101 4.5005
R52489 VINP.n320 VINP.n101 4.5005
R52490 VINP.n255 VINP.n101 4.5005
R52491 VINP.n322 VINP.n101 4.5005
R52492 VINP.n254 VINP.n101 4.5005
R52493 VINP.n324 VINP.n101 4.5005
R52494 VINP.n253 VINP.n101 4.5005
R52495 VINP.n326 VINP.n101 4.5005
R52496 VINP.n252 VINP.n101 4.5005
R52497 VINP.n328 VINP.n101 4.5005
R52498 VINP.n251 VINP.n101 4.5005
R52499 VINP.n330 VINP.n101 4.5005
R52500 VINP.n250 VINP.n101 4.5005
R52501 VINP.n332 VINP.n101 4.5005
R52502 VINP.n249 VINP.n101 4.5005
R52503 VINP.n334 VINP.n101 4.5005
R52504 VINP.n248 VINP.n101 4.5005
R52505 VINP.n336 VINP.n101 4.5005
R52506 VINP.n247 VINP.n101 4.5005
R52507 VINP.n338 VINP.n101 4.5005
R52508 VINP.n246 VINP.n101 4.5005
R52509 VINP.n340 VINP.n101 4.5005
R52510 VINP.n245 VINP.n101 4.5005
R52511 VINP.n342 VINP.n101 4.5005
R52512 VINP.n244 VINP.n101 4.5005
R52513 VINP.n344 VINP.n101 4.5005
R52514 VINP.n243 VINP.n101 4.5005
R52515 VINP.n346 VINP.n101 4.5005
R52516 VINP.n242 VINP.n101 4.5005
R52517 VINP.n348 VINP.n101 4.5005
R52518 VINP.n241 VINP.n101 4.5005
R52519 VINP.n350 VINP.n101 4.5005
R52520 VINP.n240 VINP.n101 4.5005
R52521 VINP.n352 VINP.n101 4.5005
R52522 VINP.n239 VINP.n101 4.5005
R52523 VINP.n354 VINP.n101 4.5005
R52524 VINP.n238 VINP.n101 4.5005
R52525 VINP.n356 VINP.n101 4.5005
R52526 VINP.n237 VINP.n101 4.5005
R52527 VINP.n358 VINP.n101 4.5005
R52528 VINP.n236 VINP.n101 4.5005
R52529 VINP.n360 VINP.n101 4.5005
R52530 VINP.n235 VINP.n101 4.5005
R52531 VINP.n362 VINP.n101 4.5005
R52532 VINP.n234 VINP.n101 4.5005
R52533 VINP.n364 VINP.n101 4.5005
R52534 VINP.n233 VINP.n101 4.5005
R52535 VINP.n366 VINP.n101 4.5005
R52536 VINP.n232 VINP.n101 4.5005
R52537 VINP.n368 VINP.n101 4.5005
R52538 VINP.n231 VINP.n101 4.5005
R52539 VINP.n370 VINP.n101 4.5005
R52540 VINP.n230 VINP.n101 4.5005
R52541 VINP.n372 VINP.n101 4.5005
R52542 VINP.n229 VINP.n101 4.5005
R52543 VINP.n374 VINP.n101 4.5005
R52544 VINP.n228 VINP.n101 4.5005
R52545 VINP.n376 VINP.n101 4.5005
R52546 VINP.n227 VINP.n101 4.5005
R52547 VINP.n378 VINP.n101 4.5005
R52548 VINP.n226 VINP.n101 4.5005
R52549 VINP.n380 VINP.n101 4.5005
R52550 VINP.n225 VINP.n101 4.5005
R52551 VINP.n382 VINP.n101 4.5005
R52552 VINP.n224 VINP.n101 4.5005
R52553 VINP.n384 VINP.n101 4.5005
R52554 VINP.n223 VINP.n101 4.5005
R52555 VINP.n386 VINP.n101 4.5005
R52556 VINP.n222 VINP.n101 4.5005
R52557 VINP.n388 VINP.n101 4.5005
R52558 VINP.n221 VINP.n101 4.5005
R52559 VINP.n390 VINP.n101 4.5005
R52560 VINP.n220 VINP.n101 4.5005
R52561 VINP.n392 VINP.n101 4.5005
R52562 VINP.n219 VINP.n101 4.5005
R52563 VINP.n394 VINP.n101 4.5005
R52564 VINP.n218 VINP.n101 4.5005
R52565 VINP.n396 VINP.n101 4.5005
R52566 VINP.n217 VINP.n101 4.5005
R52567 VINP.n398 VINP.n101 4.5005
R52568 VINP.n216 VINP.n101 4.5005
R52569 VINP.n400 VINP.n101 4.5005
R52570 VINP.n215 VINP.n101 4.5005
R52571 VINP.n654 VINP.n101 4.5005
R52572 VINP.n656 VINP.n101 4.5005
R52573 VINP.n101 VINP.n0 4.5005
R52574 VINP.n278 VINP.n200 4.5005
R52575 VINP.n276 VINP.n200 4.5005
R52576 VINP.n280 VINP.n200 4.5005
R52577 VINP.n275 VINP.n200 4.5005
R52578 VINP.n282 VINP.n200 4.5005
R52579 VINP.n274 VINP.n200 4.5005
R52580 VINP.n284 VINP.n200 4.5005
R52581 VINP.n273 VINP.n200 4.5005
R52582 VINP.n286 VINP.n200 4.5005
R52583 VINP.n272 VINP.n200 4.5005
R52584 VINP.n288 VINP.n200 4.5005
R52585 VINP.n271 VINP.n200 4.5005
R52586 VINP.n290 VINP.n200 4.5005
R52587 VINP.n270 VINP.n200 4.5005
R52588 VINP.n292 VINP.n200 4.5005
R52589 VINP.n269 VINP.n200 4.5005
R52590 VINP.n294 VINP.n200 4.5005
R52591 VINP.n268 VINP.n200 4.5005
R52592 VINP.n296 VINP.n200 4.5005
R52593 VINP.n267 VINP.n200 4.5005
R52594 VINP.n298 VINP.n200 4.5005
R52595 VINP.n266 VINP.n200 4.5005
R52596 VINP.n300 VINP.n200 4.5005
R52597 VINP.n265 VINP.n200 4.5005
R52598 VINP.n302 VINP.n200 4.5005
R52599 VINP.n264 VINP.n200 4.5005
R52600 VINP.n304 VINP.n200 4.5005
R52601 VINP.n263 VINP.n200 4.5005
R52602 VINP.n306 VINP.n200 4.5005
R52603 VINP.n262 VINP.n200 4.5005
R52604 VINP.n308 VINP.n200 4.5005
R52605 VINP.n261 VINP.n200 4.5005
R52606 VINP.n310 VINP.n200 4.5005
R52607 VINP.n260 VINP.n200 4.5005
R52608 VINP.n312 VINP.n200 4.5005
R52609 VINP.n259 VINP.n200 4.5005
R52610 VINP.n314 VINP.n200 4.5005
R52611 VINP.n258 VINP.n200 4.5005
R52612 VINP.n316 VINP.n200 4.5005
R52613 VINP.n257 VINP.n200 4.5005
R52614 VINP.n318 VINP.n200 4.5005
R52615 VINP.n256 VINP.n200 4.5005
R52616 VINP.n320 VINP.n200 4.5005
R52617 VINP.n255 VINP.n200 4.5005
R52618 VINP.n322 VINP.n200 4.5005
R52619 VINP.n254 VINP.n200 4.5005
R52620 VINP.n324 VINP.n200 4.5005
R52621 VINP.n253 VINP.n200 4.5005
R52622 VINP.n326 VINP.n200 4.5005
R52623 VINP.n252 VINP.n200 4.5005
R52624 VINP.n328 VINP.n200 4.5005
R52625 VINP.n251 VINP.n200 4.5005
R52626 VINP.n330 VINP.n200 4.5005
R52627 VINP.n250 VINP.n200 4.5005
R52628 VINP.n332 VINP.n200 4.5005
R52629 VINP.n249 VINP.n200 4.5005
R52630 VINP.n334 VINP.n200 4.5005
R52631 VINP.n248 VINP.n200 4.5005
R52632 VINP.n336 VINP.n200 4.5005
R52633 VINP.n247 VINP.n200 4.5005
R52634 VINP.n338 VINP.n200 4.5005
R52635 VINP.n246 VINP.n200 4.5005
R52636 VINP.n340 VINP.n200 4.5005
R52637 VINP.n245 VINP.n200 4.5005
R52638 VINP.n342 VINP.n200 4.5005
R52639 VINP.n244 VINP.n200 4.5005
R52640 VINP.n344 VINP.n200 4.5005
R52641 VINP.n243 VINP.n200 4.5005
R52642 VINP.n346 VINP.n200 4.5005
R52643 VINP.n242 VINP.n200 4.5005
R52644 VINP.n348 VINP.n200 4.5005
R52645 VINP.n241 VINP.n200 4.5005
R52646 VINP.n350 VINP.n200 4.5005
R52647 VINP.n240 VINP.n200 4.5005
R52648 VINP.n352 VINP.n200 4.5005
R52649 VINP.n239 VINP.n200 4.5005
R52650 VINP.n354 VINP.n200 4.5005
R52651 VINP.n238 VINP.n200 4.5005
R52652 VINP.n356 VINP.n200 4.5005
R52653 VINP.n237 VINP.n200 4.5005
R52654 VINP.n358 VINP.n200 4.5005
R52655 VINP.n236 VINP.n200 4.5005
R52656 VINP.n360 VINP.n200 4.5005
R52657 VINP.n235 VINP.n200 4.5005
R52658 VINP.n362 VINP.n200 4.5005
R52659 VINP.n234 VINP.n200 4.5005
R52660 VINP.n364 VINP.n200 4.5005
R52661 VINP.n233 VINP.n200 4.5005
R52662 VINP.n366 VINP.n200 4.5005
R52663 VINP.n232 VINP.n200 4.5005
R52664 VINP.n368 VINP.n200 4.5005
R52665 VINP.n231 VINP.n200 4.5005
R52666 VINP.n370 VINP.n200 4.5005
R52667 VINP.n230 VINP.n200 4.5005
R52668 VINP.n372 VINP.n200 4.5005
R52669 VINP.n229 VINP.n200 4.5005
R52670 VINP.n374 VINP.n200 4.5005
R52671 VINP.n228 VINP.n200 4.5005
R52672 VINP.n376 VINP.n200 4.5005
R52673 VINP.n227 VINP.n200 4.5005
R52674 VINP.n378 VINP.n200 4.5005
R52675 VINP.n226 VINP.n200 4.5005
R52676 VINP.n380 VINP.n200 4.5005
R52677 VINP.n225 VINP.n200 4.5005
R52678 VINP.n382 VINP.n200 4.5005
R52679 VINP.n224 VINP.n200 4.5005
R52680 VINP.n384 VINP.n200 4.5005
R52681 VINP.n223 VINP.n200 4.5005
R52682 VINP.n386 VINP.n200 4.5005
R52683 VINP.n222 VINP.n200 4.5005
R52684 VINP.n388 VINP.n200 4.5005
R52685 VINP.n221 VINP.n200 4.5005
R52686 VINP.n390 VINP.n200 4.5005
R52687 VINP.n220 VINP.n200 4.5005
R52688 VINP.n392 VINP.n200 4.5005
R52689 VINP.n219 VINP.n200 4.5005
R52690 VINP.n394 VINP.n200 4.5005
R52691 VINP.n218 VINP.n200 4.5005
R52692 VINP.n396 VINP.n200 4.5005
R52693 VINP.n217 VINP.n200 4.5005
R52694 VINP.n398 VINP.n200 4.5005
R52695 VINP.n216 VINP.n200 4.5005
R52696 VINP.n400 VINP.n200 4.5005
R52697 VINP.n215 VINP.n200 4.5005
R52698 VINP.n654 VINP.n200 4.5005
R52699 VINP.n656 VINP.n200 4.5005
R52700 VINP.n200 VINP.n0 4.5005
R52701 VINP.n278 VINP.n100 4.5005
R52702 VINP.n276 VINP.n100 4.5005
R52703 VINP.n280 VINP.n100 4.5005
R52704 VINP.n275 VINP.n100 4.5005
R52705 VINP.n282 VINP.n100 4.5005
R52706 VINP.n274 VINP.n100 4.5005
R52707 VINP.n284 VINP.n100 4.5005
R52708 VINP.n273 VINP.n100 4.5005
R52709 VINP.n286 VINP.n100 4.5005
R52710 VINP.n272 VINP.n100 4.5005
R52711 VINP.n288 VINP.n100 4.5005
R52712 VINP.n271 VINP.n100 4.5005
R52713 VINP.n290 VINP.n100 4.5005
R52714 VINP.n270 VINP.n100 4.5005
R52715 VINP.n292 VINP.n100 4.5005
R52716 VINP.n269 VINP.n100 4.5005
R52717 VINP.n294 VINP.n100 4.5005
R52718 VINP.n268 VINP.n100 4.5005
R52719 VINP.n296 VINP.n100 4.5005
R52720 VINP.n267 VINP.n100 4.5005
R52721 VINP.n298 VINP.n100 4.5005
R52722 VINP.n266 VINP.n100 4.5005
R52723 VINP.n300 VINP.n100 4.5005
R52724 VINP.n265 VINP.n100 4.5005
R52725 VINP.n302 VINP.n100 4.5005
R52726 VINP.n264 VINP.n100 4.5005
R52727 VINP.n304 VINP.n100 4.5005
R52728 VINP.n263 VINP.n100 4.5005
R52729 VINP.n306 VINP.n100 4.5005
R52730 VINP.n262 VINP.n100 4.5005
R52731 VINP.n308 VINP.n100 4.5005
R52732 VINP.n261 VINP.n100 4.5005
R52733 VINP.n310 VINP.n100 4.5005
R52734 VINP.n260 VINP.n100 4.5005
R52735 VINP.n312 VINP.n100 4.5005
R52736 VINP.n259 VINP.n100 4.5005
R52737 VINP.n314 VINP.n100 4.5005
R52738 VINP.n258 VINP.n100 4.5005
R52739 VINP.n316 VINP.n100 4.5005
R52740 VINP.n257 VINP.n100 4.5005
R52741 VINP.n318 VINP.n100 4.5005
R52742 VINP.n256 VINP.n100 4.5005
R52743 VINP.n320 VINP.n100 4.5005
R52744 VINP.n255 VINP.n100 4.5005
R52745 VINP.n322 VINP.n100 4.5005
R52746 VINP.n254 VINP.n100 4.5005
R52747 VINP.n324 VINP.n100 4.5005
R52748 VINP.n253 VINP.n100 4.5005
R52749 VINP.n326 VINP.n100 4.5005
R52750 VINP.n252 VINP.n100 4.5005
R52751 VINP.n328 VINP.n100 4.5005
R52752 VINP.n251 VINP.n100 4.5005
R52753 VINP.n330 VINP.n100 4.5005
R52754 VINP.n250 VINP.n100 4.5005
R52755 VINP.n332 VINP.n100 4.5005
R52756 VINP.n249 VINP.n100 4.5005
R52757 VINP.n334 VINP.n100 4.5005
R52758 VINP.n248 VINP.n100 4.5005
R52759 VINP.n336 VINP.n100 4.5005
R52760 VINP.n247 VINP.n100 4.5005
R52761 VINP.n338 VINP.n100 4.5005
R52762 VINP.n246 VINP.n100 4.5005
R52763 VINP.n340 VINP.n100 4.5005
R52764 VINP.n245 VINP.n100 4.5005
R52765 VINP.n342 VINP.n100 4.5005
R52766 VINP.n244 VINP.n100 4.5005
R52767 VINP.n344 VINP.n100 4.5005
R52768 VINP.n243 VINP.n100 4.5005
R52769 VINP.n346 VINP.n100 4.5005
R52770 VINP.n242 VINP.n100 4.5005
R52771 VINP.n348 VINP.n100 4.5005
R52772 VINP.n241 VINP.n100 4.5005
R52773 VINP.n350 VINP.n100 4.5005
R52774 VINP.n240 VINP.n100 4.5005
R52775 VINP.n352 VINP.n100 4.5005
R52776 VINP.n239 VINP.n100 4.5005
R52777 VINP.n354 VINP.n100 4.5005
R52778 VINP.n238 VINP.n100 4.5005
R52779 VINP.n356 VINP.n100 4.5005
R52780 VINP.n237 VINP.n100 4.5005
R52781 VINP.n358 VINP.n100 4.5005
R52782 VINP.n236 VINP.n100 4.5005
R52783 VINP.n360 VINP.n100 4.5005
R52784 VINP.n235 VINP.n100 4.5005
R52785 VINP.n362 VINP.n100 4.5005
R52786 VINP.n234 VINP.n100 4.5005
R52787 VINP.n364 VINP.n100 4.5005
R52788 VINP.n233 VINP.n100 4.5005
R52789 VINP.n366 VINP.n100 4.5005
R52790 VINP.n232 VINP.n100 4.5005
R52791 VINP.n368 VINP.n100 4.5005
R52792 VINP.n231 VINP.n100 4.5005
R52793 VINP.n370 VINP.n100 4.5005
R52794 VINP.n230 VINP.n100 4.5005
R52795 VINP.n372 VINP.n100 4.5005
R52796 VINP.n229 VINP.n100 4.5005
R52797 VINP.n374 VINP.n100 4.5005
R52798 VINP.n228 VINP.n100 4.5005
R52799 VINP.n376 VINP.n100 4.5005
R52800 VINP.n227 VINP.n100 4.5005
R52801 VINP.n378 VINP.n100 4.5005
R52802 VINP.n226 VINP.n100 4.5005
R52803 VINP.n380 VINP.n100 4.5005
R52804 VINP.n225 VINP.n100 4.5005
R52805 VINP.n382 VINP.n100 4.5005
R52806 VINP.n224 VINP.n100 4.5005
R52807 VINP.n384 VINP.n100 4.5005
R52808 VINP.n223 VINP.n100 4.5005
R52809 VINP.n386 VINP.n100 4.5005
R52810 VINP.n222 VINP.n100 4.5005
R52811 VINP.n388 VINP.n100 4.5005
R52812 VINP.n221 VINP.n100 4.5005
R52813 VINP.n390 VINP.n100 4.5005
R52814 VINP.n220 VINP.n100 4.5005
R52815 VINP.n392 VINP.n100 4.5005
R52816 VINP.n219 VINP.n100 4.5005
R52817 VINP.n394 VINP.n100 4.5005
R52818 VINP.n218 VINP.n100 4.5005
R52819 VINP.n396 VINP.n100 4.5005
R52820 VINP.n217 VINP.n100 4.5005
R52821 VINP.n398 VINP.n100 4.5005
R52822 VINP.n216 VINP.n100 4.5005
R52823 VINP.n400 VINP.n100 4.5005
R52824 VINP.n215 VINP.n100 4.5005
R52825 VINP.n654 VINP.n100 4.5005
R52826 VINP.n656 VINP.n100 4.5005
R52827 VINP.n100 VINP.n0 4.5005
R52828 VINP.n278 VINP.n201 4.5005
R52829 VINP.n276 VINP.n201 4.5005
R52830 VINP.n280 VINP.n201 4.5005
R52831 VINP.n275 VINP.n201 4.5005
R52832 VINP.n282 VINP.n201 4.5005
R52833 VINP.n274 VINP.n201 4.5005
R52834 VINP.n284 VINP.n201 4.5005
R52835 VINP.n273 VINP.n201 4.5005
R52836 VINP.n286 VINP.n201 4.5005
R52837 VINP.n272 VINP.n201 4.5005
R52838 VINP.n288 VINP.n201 4.5005
R52839 VINP.n271 VINP.n201 4.5005
R52840 VINP.n290 VINP.n201 4.5005
R52841 VINP.n270 VINP.n201 4.5005
R52842 VINP.n292 VINP.n201 4.5005
R52843 VINP.n269 VINP.n201 4.5005
R52844 VINP.n294 VINP.n201 4.5005
R52845 VINP.n268 VINP.n201 4.5005
R52846 VINP.n296 VINP.n201 4.5005
R52847 VINP.n267 VINP.n201 4.5005
R52848 VINP.n298 VINP.n201 4.5005
R52849 VINP.n266 VINP.n201 4.5005
R52850 VINP.n300 VINP.n201 4.5005
R52851 VINP.n265 VINP.n201 4.5005
R52852 VINP.n302 VINP.n201 4.5005
R52853 VINP.n264 VINP.n201 4.5005
R52854 VINP.n304 VINP.n201 4.5005
R52855 VINP.n263 VINP.n201 4.5005
R52856 VINP.n306 VINP.n201 4.5005
R52857 VINP.n262 VINP.n201 4.5005
R52858 VINP.n308 VINP.n201 4.5005
R52859 VINP.n261 VINP.n201 4.5005
R52860 VINP.n310 VINP.n201 4.5005
R52861 VINP.n260 VINP.n201 4.5005
R52862 VINP.n312 VINP.n201 4.5005
R52863 VINP.n259 VINP.n201 4.5005
R52864 VINP.n314 VINP.n201 4.5005
R52865 VINP.n258 VINP.n201 4.5005
R52866 VINP.n316 VINP.n201 4.5005
R52867 VINP.n257 VINP.n201 4.5005
R52868 VINP.n318 VINP.n201 4.5005
R52869 VINP.n256 VINP.n201 4.5005
R52870 VINP.n320 VINP.n201 4.5005
R52871 VINP.n255 VINP.n201 4.5005
R52872 VINP.n322 VINP.n201 4.5005
R52873 VINP.n254 VINP.n201 4.5005
R52874 VINP.n324 VINP.n201 4.5005
R52875 VINP.n253 VINP.n201 4.5005
R52876 VINP.n326 VINP.n201 4.5005
R52877 VINP.n252 VINP.n201 4.5005
R52878 VINP.n328 VINP.n201 4.5005
R52879 VINP.n251 VINP.n201 4.5005
R52880 VINP.n330 VINP.n201 4.5005
R52881 VINP.n250 VINP.n201 4.5005
R52882 VINP.n332 VINP.n201 4.5005
R52883 VINP.n249 VINP.n201 4.5005
R52884 VINP.n334 VINP.n201 4.5005
R52885 VINP.n248 VINP.n201 4.5005
R52886 VINP.n336 VINP.n201 4.5005
R52887 VINP.n247 VINP.n201 4.5005
R52888 VINP.n338 VINP.n201 4.5005
R52889 VINP.n246 VINP.n201 4.5005
R52890 VINP.n340 VINP.n201 4.5005
R52891 VINP.n245 VINP.n201 4.5005
R52892 VINP.n342 VINP.n201 4.5005
R52893 VINP.n244 VINP.n201 4.5005
R52894 VINP.n344 VINP.n201 4.5005
R52895 VINP.n243 VINP.n201 4.5005
R52896 VINP.n346 VINP.n201 4.5005
R52897 VINP.n242 VINP.n201 4.5005
R52898 VINP.n348 VINP.n201 4.5005
R52899 VINP.n241 VINP.n201 4.5005
R52900 VINP.n350 VINP.n201 4.5005
R52901 VINP.n240 VINP.n201 4.5005
R52902 VINP.n352 VINP.n201 4.5005
R52903 VINP.n239 VINP.n201 4.5005
R52904 VINP.n354 VINP.n201 4.5005
R52905 VINP.n238 VINP.n201 4.5005
R52906 VINP.n356 VINP.n201 4.5005
R52907 VINP.n237 VINP.n201 4.5005
R52908 VINP.n358 VINP.n201 4.5005
R52909 VINP.n236 VINP.n201 4.5005
R52910 VINP.n360 VINP.n201 4.5005
R52911 VINP.n235 VINP.n201 4.5005
R52912 VINP.n362 VINP.n201 4.5005
R52913 VINP.n234 VINP.n201 4.5005
R52914 VINP.n364 VINP.n201 4.5005
R52915 VINP.n233 VINP.n201 4.5005
R52916 VINP.n366 VINP.n201 4.5005
R52917 VINP.n232 VINP.n201 4.5005
R52918 VINP.n368 VINP.n201 4.5005
R52919 VINP.n231 VINP.n201 4.5005
R52920 VINP.n370 VINP.n201 4.5005
R52921 VINP.n230 VINP.n201 4.5005
R52922 VINP.n372 VINP.n201 4.5005
R52923 VINP.n229 VINP.n201 4.5005
R52924 VINP.n374 VINP.n201 4.5005
R52925 VINP.n228 VINP.n201 4.5005
R52926 VINP.n376 VINP.n201 4.5005
R52927 VINP.n227 VINP.n201 4.5005
R52928 VINP.n378 VINP.n201 4.5005
R52929 VINP.n226 VINP.n201 4.5005
R52930 VINP.n380 VINP.n201 4.5005
R52931 VINP.n225 VINP.n201 4.5005
R52932 VINP.n382 VINP.n201 4.5005
R52933 VINP.n224 VINP.n201 4.5005
R52934 VINP.n384 VINP.n201 4.5005
R52935 VINP.n223 VINP.n201 4.5005
R52936 VINP.n386 VINP.n201 4.5005
R52937 VINP.n222 VINP.n201 4.5005
R52938 VINP.n388 VINP.n201 4.5005
R52939 VINP.n221 VINP.n201 4.5005
R52940 VINP.n390 VINP.n201 4.5005
R52941 VINP.n220 VINP.n201 4.5005
R52942 VINP.n392 VINP.n201 4.5005
R52943 VINP.n219 VINP.n201 4.5005
R52944 VINP.n394 VINP.n201 4.5005
R52945 VINP.n218 VINP.n201 4.5005
R52946 VINP.n396 VINP.n201 4.5005
R52947 VINP.n217 VINP.n201 4.5005
R52948 VINP.n398 VINP.n201 4.5005
R52949 VINP.n216 VINP.n201 4.5005
R52950 VINP.n400 VINP.n201 4.5005
R52951 VINP.n215 VINP.n201 4.5005
R52952 VINP.n654 VINP.n201 4.5005
R52953 VINP.n656 VINP.n201 4.5005
R52954 VINP.n201 VINP.n0 4.5005
R52955 VINP.n278 VINP.n99 4.5005
R52956 VINP.n276 VINP.n99 4.5005
R52957 VINP.n280 VINP.n99 4.5005
R52958 VINP.n275 VINP.n99 4.5005
R52959 VINP.n282 VINP.n99 4.5005
R52960 VINP.n274 VINP.n99 4.5005
R52961 VINP.n284 VINP.n99 4.5005
R52962 VINP.n273 VINP.n99 4.5005
R52963 VINP.n286 VINP.n99 4.5005
R52964 VINP.n272 VINP.n99 4.5005
R52965 VINP.n288 VINP.n99 4.5005
R52966 VINP.n271 VINP.n99 4.5005
R52967 VINP.n290 VINP.n99 4.5005
R52968 VINP.n270 VINP.n99 4.5005
R52969 VINP.n292 VINP.n99 4.5005
R52970 VINP.n269 VINP.n99 4.5005
R52971 VINP.n294 VINP.n99 4.5005
R52972 VINP.n268 VINP.n99 4.5005
R52973 VINP.n296 VINP.n99 4.5005
R52974 VINP.n267 VINP.n99 4.5005
R52975 VINP.n298 VINP.n99 4.5005
R52976 VINP.n266 VINP.n99 4.5005
R52977 VINP.n300 VINP.n99 4.5005
R52978 VINP.n265 VINP.n99 4.5005
R52979 VINP.n302 VINP.n99 4.5005
R52980 VINP.n264 VINP.n99 4.5005
R52981 VINP.n304 VINP.n99 4.5005
R52982 VINP.n263 VINP.n99 4.5005
R52983 VINP.n306 VINP.n99 4.5005
R52984 VINP.n262 VINP.n99 4.5005
R52985 VINP.n308 VINP.n99 4.5005
R52986 VINP.n261 VINP.n99 4.5005
R52987 VINP.n310 VINP.n99 4.5005
R52988 VINP.n260 VINP.n99 4.5005
R52989 VINP.n312 VINP.n99 4.5005
R52990 VINP.n259 VINP.n99 4.5005
R52991 VINP.n314 VINP.n99 4.5005
R52992 VINP.n258 VINP.n99 4.5005
R52993 VINP.n316 VINP.n99 4.5005
R52994 VINP.n257 VINP.n99 4.5005
R52995 VINP.n318 VINP.n99 4.5005
R52996 VINP.n256 VINP.n99 4.5005
R52997 VINP.n320 VINP.n99 4.5005
R52998 VINP.n255 VINP.n99 4.5005
R52999 VINP.n322 VINP.n99 4.5005
R53000 VINP.n254 VINP.n99 4.5005
R53001 VINP.n324 VINP.n99 4.5005
R53002 VINP.n253 VINP.n99 4.5005
R53003 VINP.n326 VINP.n99 4.5005
R53004 VINP.n252 VINP.n99 4.5005
R53005 VINP.n328 VINP.n99 4.5005
R53006 VINP.n251 VINP.n99 4.5005
R53007 VINP.n330 VINP.n99 4.5005
R53008 VINP.n250 VINP.n99 4.5005
R53009 VINP.n332 VINP.n99 4.5005
R53010 VINP.n249 VINP.n99 4.5005
R53011 VINP.n334 VINP.n99 4.5005
R53012 VINP.n248 VINP.n99 4.5005
R53013 VINP.n336 VINP.n99 4.5005
R53014 VINP.n247 VINP.n99 4.5005
R53015 VINP.n338 VINP.n99 4.5005
R53016 VINP.n246 VINP.n99 4.5005
R53017 VINP.n340 VINP.n99 4.5005
R53018 VINP.n245 VINP.n99 4.5005
R53019 VINP.n342 VINP.n99 4.5005
R53020 VINP.n244 VINP.n99 4.5005
R53021 VINP.n344 VINP.n99 4.5005
R53022 VINP.n243 VINP.n99 4.5005
R53023 VINP.n346 VINP.n99 4.5005
R53024 VINP.n242 VINP.n99 4.5005
R53025 VINP.n348 VINP.n99 4.5005
R53026 VINP.n241 VINP.n99 4.5005
R53027 VINP.n350 VINP.n99 4.5005
R53028 VINP.n240 VINP.n99 4.5005
R53029 VINP.n352 VINP.n99 4.5005
R53030 VINP.n239 VINP.n99 4.5005
R53031 VINP.n354 VINP.n99 4.5005
R53032 VINP.n238 VINP.n99 4.5005
R53033 VINP.n356 VINP.n99 4.5005
R53034 VINP.n237 VINP.n99 4.5005
R53035 VINP.n358 VINP.n99 4.5005
R53036 VINP.n236 VINP.n99 4.5005
R53037 VINP.n360 VINP.n99 4.5005
R53038 VINP.n235 VINP.n99 4.5005
R53039 VINP.n362 VINP.n99 4.5005
R53040 VINP.n234 VINP.n99 4.5005
R53041 VINP.n364 VINP.n99 4.5005
R53042 VINP.n233 VINP.n99 4.5005
R53043 VINP.n366 VINP.n99 4.5005
R53044 VINP.n232 VINP.n99 4.5005
R53045 VINP.n368 VINP.n99 4.5005
R53046 VINP.n231 VINP.n99 4.5005
R53047 VINP.n370 VINP.n99 4.5005
R53048 VINP.n230 VINP.n99 4.5005
R53049 VINP.n372 VINP.n99 4.5005
R53050 VINP.n229 VINP.n99 4.5005
R53051 VINP.n374 VINP.n99 4.5005
R53052 VINP.n228 VINP.n99 4.5005
R53053 VINP.n376 VINP.n99 4.5005
R53054 VINP.n227 VINP.n99 4.5005
R53055 VINP.n378 VINP.n99 4.5005
R53056 VINP.n226 VINP.n99 4.5005
R53057 VINP.n380 VINP.n99 4.5005
R53058 VINP.n225 VINP.n99 4.5005
R53059 VINP.n382 VINP.n99 4.5005
R53060 VINP.n224 VINP.n99 4.5005
R53061 VINP.n384 VINP.n99 4.5005
R53062 VINP.n223 VINP.n99 4.5005
R53063 VINP.n386 VINP.n99 4.5005
R53064 VINP.n222 VINP.n99 4.5005
R53065 VINP.n388 VINP.n99 4.5005
R53066 VINP.n221 VINP.n99 4.5005
R53067 VINP.n390 VINP.n99 4.5005
R53068 VINP.n220 VINP.n99 4.5005
R53069 VINP.n392 VINP.n99 4.5005
R53070 VINP.n219 VINP.n99 4.5005
R53071 VINP.n394 VINP.n99 4.5005
R53072 VINP.n218 VINP.n99 4.5005
R53073 VINP.n396 VINP.n99 4.5005
R53074 VINP.n217 VINP.n99 4.5005
R53075 VINP.n398 VINP.n99 4.5005
R53076 VINP.n216 VINP.n99 4.5005
R53077 VINP.n400 VINP.n99 4.5005
R53078 VINP.n215 VINP.n99 4.5005
R53079 VINP.n654 VINP.n99 4.5005
R53080 VINP.n656 VINP.n99 4.5005
R53081 VINP.n99 VINP.n0 4.5005
R53082 VINP.n278 VINP.n202 4.5005
R53083 VINP.n276 VINP.n202 4.5005
R53084 VINP.n280 VINP.n202 4.5005
R53085 VINP.n275 VINP.n202 4.5005
R53086 VINP.n282 VINP.n202 4.5005
R53087 VINP.n274 VINP.n202 4.5005
R53088 VINP.n284 VINP.n202 4.5005
R53089 VINP.n273 VINP.n202 4.5005
R53090 VINP.n286 VINP.n202 4.5005
R53091 VINP.n272 VINP.n202 4.5005
R53092 VINP.n288 VINP.n202 4.5005
R53093 VINP.n271 VINP.n202 4.5005
R53094 VINP.n290 VINP.n202 4.5005
R53095 VINP.n270 VINP.n202 4.5005
R53096 VINP.n292 VINP.n202 4.5005
R53097 VINP.n269 VINP.n202 4.5005
R53098 VINP.n294 VINP.n202 4.5005
R53099 VINP.n268 VINP.n202 4.5005
R53100 VINP.n296 VINP.n202 4.5005
R53101 VINP.n267 VINP.n202 4.5005
R53102 VINP.n298 VINP.n202 4.5005
R53103 VINP.n266 VINP.n202 4.5005
R53104 VINP.n300 VINP.n202 4.5005
R53105 VINP.n265 VINP.n202 4.5005
R53106 VINP.n302 VINP.n202 4.5005
R53107 VINP.n264 VINP.n202 4.5005
R53108 VINP.n304 VINP.n202 4.5005
R53109 VINP.n263 VINP.n202 4.5005
R53110 VINP.n306 VINP.n202 4.5005
R53111 VINP.n262 VINP.n202 4.5005
R53112 VINP.n308 VINP.n202 4.5005
R53113 VINP.n261 VINP.n202 4.5005
R53114 VINP.n310 VINP.n202 4.5005
R53115 VINP.n260 VINP.n202 4.5005
R53116 VINP.n312 VINP.n202 4.5005
R53117 VINP.n259 VINP.n202 4.5005
R53118 VINP.n314 VINP.n202 4.5005
R53119 VINP.n258 VINP.n202 4.5005
R53120 VINP.n316 VINP.n202 4.5005
R53121 VINP.n257 VINP.n202 4.5005
R53122 VINP.n318 VINP.n202 4.5005
R53123 VINP.n256 VINP.n202 4.5005
R53124 VINP.n320 VINP.n202 4.5005
R53125 VINP.n255 VINP.n202 4.5005
R53126 VINP.n322 VINP.n202 4.5005
R53127 VINP.n254 VINP.n202 4.5005
R53128 VINP.n324 VINP.n202 4.5005
R53129 VINP.n253 VINP.n202 4.5005
R53130 VINP.n326 VINP.n202 4.5005
R53131 VINP.n252 VINP.n202 4.5005
R53132 VINP.n328 VINP.n202 4.5005
R53133 VINP.n251 VINP.n202 4.5005
R53134 VINP.n330 VINP.n202 4.5005
R53135 VINP.n250 VINP.n202 4.5005
R53136 VINP.n332 VINP.n202 4.5005
R53137 VINP.n249 VINP.n202 4.5005
R53138 VINP.n334 VINP.n202 4.5005
R53139 VINP.n248 VINP.n202 4.5005
R53140 VINP.n336 VINP.n202 4.5005
R53141 VINP.n247 VINP.n202 4.5005
R53142 VINP.n338 VINP.n202 4.5005
R53143 VINP.n246 VINP.n202 4.5005
R53144 VINP.n340 VINP.n202 4.5005
R53145 VINP.n245 VINP.n202 4.5005
R53146 VINP.n342 VINP.n202 4.5005
R53147 VINP.n244 VINP.n202 4.5005
R53148 VINP.n344 VINP.n202 4.5005
R53149 VINP.n243 VINP.n202 4.5005
R53150 VINP.n346 VINP.n202 4.5005
R53151 VINP.n242 VINP.n202 4.5005
R53152 VINP.n348 VINP.n202 4.5005
R53153 VINP.n241 VINP.n202 4.5005
R53154 VINP.n350 VINP.n202 4.5005
R53155 VINP.n240 VINP.n202 4.5005
R53156 VINP.n352 VINP.n202 4.5005
R53157 VINP.n239 VINP.n202 4.5005
R53158 VINP.n354 VINP.n202 4.5005
R53159 VINP.n238 VINP.n202 4.5005
R53160 VINP.n356 VINP.n202 4.5005
R53161 VINP.n237 VINP.n202 4.5005
R53162 VINP.n358 VINP.n202 4.5005
R53163 VINP.n236 VINP.n202 4.5005
R53164 VINP.n360 VINP.n202 4.5005
R53165 VINP.n235 VINP.n202 4.5005
R53166 VINP.n362 VINP.n202 4.5005
R53167 VINP.n234 VINP.n202 4.5005
R53168 VINP.n364 VINP.n202 4.5005
R53169 VINP.n233 VINP.n202 4.5005
R53170 VINP.n366 VINP.n202 4.5005
R53171 VINP.n232 VINP.n202 4.5005
R53172 VINP.n368 VINP.n202 4.5005
R53173 VINP.n231 VINP.n202 4.5005
R53174 VINP.n370 VINP.n202 4.5005
R53175 VINP.n230 VINP.n202 4.5005
R53176 VINP.n372 VINP.n202 4.5005
R53177 VINP.n229 VINP.n202 4.5005
R53178 VINP.n374 VINP.n202 4.5005
R53179 VINP.n228 VINP.n202 4.5005
R53180 VINP.n376 VINP.n202 4.5005
R53181 VINP.n227 VINP.n202 4.5005
R53182 VINP.n378 VINP.n202 4.5005
R53183 VINP.n226 VINP.n202 4.5005
R53184 VINP.n380 VINP.n202 4.5005
R53185 VINP.n225 VINP.n202 4.5005
R53186 VINP.n382 VINP.n202 4.5005
R53187 VINP.n224 VINP.n202 4.5005
R53188 VINP.n384 VINP.n202 4.5005
R53189 VINP.n223 VINP.n202 4.5005
R53190 VINP.n386 VINP.n202 4.5005
R53191 VINP.n222 VINP.n202 4.5005
R53192 VINP.n388 VINP.n202 4.5005
R53193 VINP.n221 VINP.n202 4.5005
R53194 VINP.n390 VINP.n202 4.5005
R53195 VINP.n220 VINP.n202 4.5005
R53196 VINP.n392 VINP.n202 4.5005
R53197 VINP.n219 VINP.n202 4.5005
R53198 VINP.n394 VINP.n202 4.5005
R53199 VINP.n218 VINP.n202 4.5005
R53200 VINP.n396 VINP.n202 4.5005
R53201 VINP.n217 VINP.n202 4.5005
R53202 VINP.n398 VINP.n202 4.5005
R53203 VINP.n216 VINP.n202 4.5005
R53204 VINP.n400 VINP.n202 4.5005
R53205 VINP.n215 VINP.n202 4.5005
R53206 VINP.n654 VINP.n202 4.5005
R53207 VINP.n656 VINP.n202 4.5005
R53208 VINP.n202 VINP.n0 4.5005
R53209 VINP.n278 VINP.n98 4.5005
R53210 VINP.n276 VINP.n98 4.5005
R53211 VINP.n280 VINP.n98 4.5005
R53212 VINP.n275 VINP.n98 4.5005
R53213 VINP.n282 VINP.n98 4.5005
R53214 VINP.n274 VINP.n98 4.5005
R53215 VINP.n284 VINP.n98 4.5005
R53216 VINP.n273 VINP.n98 4.5005
R53217 VINP.n286 VINP.n98 4.5005
R53218 VINP.n272 VINP.n98 4.5005
R53219 VINP.n288 VINP.n98 4.5005
R53220 VINP.n271 VINP.n98 4.5005
R53221 VINP.n290 VINP.n98 4.5005
R53222 VINP.n270 VINP.n98 4.5005
R53223 VINP.n292 VINP.n98 4.5005
R53224 VINP.n269 VINP.n98 4.5005
R53225 VINP.n294 VINP.n98 4.5005
R53226 VINP.n268 VINP.n98 4.5005
R53227 VINP.n296 VINP.n98 4.5005
R53228 VINP.n267 VINP.n98 4.5005
R53229 VINP.n298 VINP.n98 4.5005
R53230 VINP.n266 VINP.n98 4.5005
R53231 VINP.n300 VINP.n98 4.5005
R53232 VINP.n265 VINP.n98 4.5005
R53233 VINP.n302 VINP.n98 4.5005
R53234 VINP.n264 VINP.n98 4.5005
R53235 VINP.n304 VINP.n98 4.5005
R53236 VINP.n263 VINP.n98 4.5005
R53237 VINP.n306 VINP.n98 4.5005
R53238 VINP.n262 VINP.n98 4.5005
R53239 VINP.n308 VINP.n98 4.5005
R53240 VINP.n261 VINP.n98 4.5005
R53241 VINP.n310 VINP.n98 4.5005
R53242 VINP.n260 VINP.n98 4.5005
R53243 VINP.n312 VINP.n98 4.5005
R53244 VINP.n259 VINP.n98 4.5005
R53245 VINP.n314 VINP.n98 4.5005
R53246 VINP.n258 VINP.n98 4.5005
R53247 VINP.n316 VINP.n98 4.5005
R53248 VINP.n257 VINP.n98 4.5005
R53249 VINP.n318 VINP.n98 4.5005
R53250 VINP.n256 VINP.n98 4.5005
R53251 VINP.n320 VINP.n98 4.5005
R53252 VINP.n255 VINP.n98 4.5005
R53253 VINP.n322 VINP.n98 4.5005
R53254 VINP.n254 VINP.n98 4.5005
R53255 VINP.n324 VINP.n98 4.5005
R53256 VINP.n253 VINP.n98 4.5005
R53257 VINP.n326 VINP.n98 4.5005
R53258 VINP.n252 VINP.n98 4.5005
R53259 VINP.n328 VINP.n98 4.5005
R53260 VINP.n251 VINP.n98 4.5005
R53261 VINP.n330 VINP.n98 4.5005
R53262 VINP.n250 VINP.n98 4.5005
R53263 VINP.n332 VINP.n98 4.5005
R53264 VINP.n249 VINP.n98 4.5005
R53265 VINP.n334 VINP.n98 4.5005
R53266 VINP.n248 VINP.n98 4.5005
R53267 VINP.n336 VINP.n98 4.5005
R53268 VINP.n247 VINP.n98 4.5005
R53269 VINP.n338 VINP.n98 4.5005
R53270 VINP.n246 VINP.n98 4.5005
R53271 VINP.n340 VINP.n98 4.5005
R53272 VINP.n245 VINP.n98 4.5005
R53273 VINP.n342 VINP.n98 4.5005
R53274 VINP.n244 VINP.n98 4.5005
R53275 VINP.n344 VINP.n98 4.5005
R53276 VINP.n243 VINP.n98 4.5005
R53277 VINP.n346 VINP.n98 4.5005
R53278 VINP.n242 VINP.n98 4.5005
R53279 VINP.n348 VINP.n98 4.5005
R53280 VINP.n241 VINP.n98 4.5005
R53281 VINP.n350 VINP.n98 4.5005
R53282 VINP.n240 VINP.n98 4.5005
R53283 VINP.n352 VINP.n98 4.5005
R53284 VINP.n239 VINP.n98 4.5005
R53285 VINP.n354 VINP.n98 4.5005
R53286 VINP.n238 VINP.n98 4.5005
R53287 VINP.n356 VINP.n98 4.5005
R53288 VINP.n237 VINP.n98 4.5005
R53289 VINP.n358 VINP.n98 4.5005
R53290 VINP.n236 VINP.n98 4.5005
R53291 VINP.n360 VINP.n98 4.5005
R53292 VINP.n235 VINP.n98 4.5005
R53293 VINP.n362 VINP.n98 4.5005
R53294 VINP.n234 VINP.n98 4.5005
R53295 VINP.n364 VINP.n98 4.5005
R53296 VINP.n233 VINP.n98 4.5005
R53297 VINP.n366 VINP.n98 4.5005
R53298 VINP.n232 VINP.n98 4.5005
R53299 VINP.n368 VINP.n98 4.5005
R53300 VINP.n231 VINP.n98 4.5005
R53301 VINP.n370 VINP.n98 4.5005
R53302 VINP.n230 VINP.n98 4.5005
R53303 VINP.n372 VINP.n98 4.5005
R53304 VINP.n229 VINP.n98 4.5005
R53305 VINP.n374 VINP.n98 4.5005
R53306 VINP.n228 VINP.n98 4.5005
R53307 VINP.n376 VINP.n98 4.5005
R53308 VINP.n227 VINP.n98 4.5005
R53309 VINP.n378 VINP.n98 4.5005
R53310 VINP.n226 VINP.n98 4.5005
R53311 VINP.n380 VINP.n98 4.5005
R53312 VINP.n225 VINP.n98 4.5005
R53313 VINP.n382 VINP.n98 4.5005
R53314 VINP.n224 VINP.n98 4.5005
R53315 VINP.n384 VINP.n98 4.5005
R53316 VINP.n223 VINP.n98 4.5005
R53317 VINP.n386 VINP.n98 4.5005
R53318 VINP.n222 VINP.n98 4.5005
R53319 VINP.n388 VINP.n98 4.5005
R53320 VINP.n221 VINP.n98 4.5005
R53321 VINP.n390 VINP.n98 4.5005
R53322 VINP.n220 VINP.n98 4.5005
R53323 VINP.n392 VINP.n98 4.5005
R53324 VINP.n219 VINP.n98 4.5005
R53325 VINP.n394 VINP.n98 4.5005
R53326 VINP.n218 VINP.n98 4.5005
R53327 VINP.n396 VINP.n98 4.5005
R53328 VINP.n217 VINP.n98 4.5005
R53329 VINP.n398 VINP.n98 4.5005
R53330 VINP.n216 VINP.n98 4.5005
R53331 VINP.n400 VINP.n98 4.5005
R53332 VINP.n215 VINP.n98 4.5005
R53333 VINP.n654 VINP.n98 4.5005
R53334 VINP.n656 VINP.n98 4.5005
R53335 VINP.n98 VINP.n0 4.5005
R53336 VINP.n278 VINP.n203 4.5005
R53337 VINP.n276 VINP.n203 4.5005
R53338 VINP.n280 VINP.n203 4.5005
R53339 VINP.n275 VINP.n203 4.5005
R53340 VINP.n282 VINP.n203 4.5005
R53341 VINP.n274 VINP.n203 4.5005
R53342 VINP.n284 VINP.n203 4.5005
R53343 VINP.n273 VINP.n203 4.5005
R53344 VINP.n286 VINP.n203 4.5005
R53345 VINP.n272 VINP.n203 4.5005
R53346 VINP.n288 VINP.n203 4.5005
R53347 VINP.n271 VINP.n203 4.5005
R53348 VINP.n290 VINP.n203 4.5005
R53349 VINP.n270 VINP.n203 4.5005
R53350 VINP.n292 VINP.n203 4.5005
R53351 VINP.n269 VINP.n203 4.5005
R53352 VINP.n294 VINP.n203 4.5005
R53353 VINP.n268 VINP.n203 4.5005
R53354 VINP.n296 VINP.n203 4.5005
R53355 VINP.n267 VINP.n203 4.5005
R53356 VINP.n298 VINP.n203 4.5005
R53357 VINP.n266 VINP.n203 4.5005
R53358 VINP.n300 VINP.n203 4.5005
R53359 VINP.n265 VINP.n203 4.5005
R53360 VINP.n302 VINP.n203 4.5005
R53361 VINP.n264 VINP.n203 4.5005
R53362 VINP.n304 VINP.n203 4.5005
R53363 VINP.n263 VINP.n203 4.5005
R53364 VINP.n306 VINP.n203 4.5005
R53365 VINP.n262 VINP.n203 4.5005
R53366 VINP.n308 VINP.n203 4.5005
R53367 VINP.n261 VINP.n203 4.5005
R53368 VINP.n310 VINP.n203 4.5005
R53369 VINP.n260 VINP.n203 4.5005
R53370 VINP.n312 VINP.n203 4.5005
R53371 VINP.n259 VINP.n203 4.5005
R53372 VINP.n314 VINP.n203 4.5005
R53373 VINP.n258 VINP.n203 4.5005
R53374 VINP.n316 VINP.n203 4.5005
R53375 VINP.n257 VINP.n203 4.5005
R53376 VINP.n318 VINP.n203 4.5005
R53377 VINP.n256 VINP.n203 4.5005
R53378 VINP.n320 VINP.n203 4.5005
R53379 VINP.n255 VINP.n203 4.5005
R53380 VINP.n322 VINP.n203 4.5005
R53381 VINP.n254 VINP.n203 4.5005
R53382 VINP.n324 VINP.n203 4.5005
R53383 VINP.n253 VINP.n203 4.5005
R53384 VINP.n326 VINP.n203 4.5005
R53385 VINP.n252 VINP.n203 4.5005
R53386 VINP.n328 VINP.n203 4.5005
R53387 VINP.n251 VINP.n203 4.5005
R53388 VINP.n330 VINP.n203 4.5005
R53389 VINP.n250 VINP.n203 4.5005
R53390 VINP.n332 VINP.n203 4.5005
R53391 VINP.n249 VINP.n203 4.5005
R53392 VINP.n334 VINP.n203 4.5005
R53393 VINP.n248 VINP.n203 4.5005
R53394 VINP.n336 VINP.n203 4.5005
R53395 VINP.n247 VINP.n203 4.5005
R53396 VINP.n338 VINP.n203 4.5005
R53397 VINP.n246 VINP.n203 4.5005
R53398 VINP.n340 VINP.n203 4.5005
R53399 VINP.n245 VINP.n203 4.5005
R53400 VINP.n342 VINP.n203 4.5005
R53401 VINP.n244 VINP.n203 4.5005
R53402 VINP.n344 VINP.n203 4.5005
R53403 VINP.n243 VINP.n203 4.5005
R53404 VINP.n346 VINP.n203 4.5005
R53405 VINP.n242 VINP.n203 4.5005
R53406 VINP.n348 VINP.n203 4.5005
R53407 VINP.n241 VINP.n203 4.5005
R53408 VINP.n350 VINP.n203 4.5005
R53409 VINP.n240 VINP.n203 4.5005
R53410 VINP.n352 VINP.n203 4.5005
R53411 VINP.n239 VINP.n203 4.5005
R53412 VINP.n354 VINP.n203 4.5005
R53413 VINP.n238 VINP.n203 4.5005
R53414 VINP.n356 VINP.n203 4.5005
R53415 VINP.n237 VINP.n203 4.5005
R53416 VINP.n358 VINP.n203 4.5005
R53417 VINP.n236 VINP.n203 4.5005
R53418 VINP.n360 VINP.n203 4.5005
R53419 VINP.n235 VINP.n203 4.5005
R53420 VINP.n362 VINP.n203 4.5005
R53421 VINP.n234 VINP.n203 4.5005
R53422 VINP.n364 VINP.n203 4.5005
R53423 VINP.n233 VINP.n203 4.5005
R53424 VINP.n366 VINP.n203 4.5005
R53425 VINP.n232 VINP.n203 4.5005
R53426 VINP.n368 VINP.n203 4.5005
R53427 VINP.n231 VINP.n203 4.5005
R53428 VINP.n370 VINP.n203 4.5005
R53429 VINP.n230 VINP.n203 4.5005
R53430 VINP.n372 VINP.n203 4.5005
R53431 VINP.n229 VINP.n203 4.5005
R53432 VINP.n374 VINP.n203 4.5005
R53433 VINP.n228 VINP.n203 4.5005
R53434 VINP.n376 VINP.n203 4.5005
R53435 VINP.n227 VINP.n203 4.5005
R53436 VINP.n378 VINP.n203 4.5005
R53437 VINP.n226 VINP.n203 4.5005
R53438 VINP.n380 VINP.n203 4.5005
R53439 VINP.n225 VINP.n203 4.5005
R53440 VINP.n382 VINP.n203 4.5005
R53441 VINP.n224 VINP.n203 4.5005
R53442 VINP.n384 VINP.n203 4.5005
R53443 VINP.n223 VINP.n203 4.5005
R53444 VINP.n386 VINP.n203 4.5005
R53445 VINP.n222 VINP.n203 4.5005
R53446 VINP.n388 VINP.n203 4.5005
R53447 VINP.n221 VINP.n203 4.5005
R53448 VINP.n390 VINP.n203 4.5005
R53449 VINP.n220 VINP.n203 4.5005
R53450 VINP.n392 VINP.n203 4.5005
R53451 VINP.n219 VINP.n203 4.5005
R53452 VINP.n394 VINP.n203 4.5005
R53453 VINP.n218 VINP.n203 4.5005
R53454 VINP.n396 VINP.n203 4.5005
R53455 VINP.n217 VINP.n203 4.5005
R53456 VINP.n398 VINP.n203 4.5005
R53457 VINP.n216 VINP.n203 4.5005
R53458 VINP.n400 VINP.n203 4.5005
R53459 VINP.n215 VINP.n203 4.5005
R53460 VINP.n654 VINP.n203 4.5005
R53461 VINP.n656 VINP.n203 4.5005
R53462 VINP.n203 VINP.n0 4.5005
R53463 VINP.n278 VINP.n97 4.5005
R53464 VINP.n276 VINP.n97 4.5005
R53465 VINP.n280 VINP.n97 4.5005
R53466 VINP.n275 VINP.n97 4.5005
R53467 VINP.n282 VINP.n97 4.5005
R53468 VINP.n274 VINP.n97 4.5005
R53469 VINP.n284 VINP.n97 4.5005
R53470 VINP.n273 VINP.n97 4.5005
R53471 VINP.n286 VINP.n97 4.5005
R53472 VINP.n272 VINP.n97 4.5005
R53473 VINP.n288 VINP.n97 4.5005
R53474 VINP.n271 VINP.n97 4.5005
R53475 VINP.n290 VINP.n97 4.5005
R53476 VINP.n270 VINP.n97 4.5005
R53477 VINP.n292 VINP.n97 4.5005
R53478 VINP.n269 VINP.n97 4.5005
R53479 VINP.n294 VINP.n97 4.5005
R53480 VINP.n268 VINP.n97 4.5005
R53481 VINP.n296 VINP.n97 4.5005
R53482 VINP.n267 VINP.n97 4.5005
R53483 VINP.n298 VINP.n97 4.5005
R53484 VINP.n266 VINP.n97 4.5005
R53485 VINP.n300 VINP.n97 4.5005
R53486 VINP.n265 VINP.n97 4.5005
R53487 VINP.n302 VINP.n97 4.5005
R53488 VINP.n264 VINP.n97 4.5005
R53489 VINP.n304 VINP.n97 4.5005
R53490 VINP.n263 VINP.n97 4.5005
R53491 VINP.n306 VINP.n97 4.5005
R53492 VINP.n262 VINP.n97 4.5005
R53493 VINP.n308 VINP.n97 4.5005
R53494 VINP.n261 VINP.n97 4.5005
R53495 VINP.n310 VINP.n97 4.5005
R53496 VINP.n260 VINP.n97 4.5005
R53497 VINP.n312 VINP.n97 4.5005
R53498 VINP.n259 VINP.n97 4.5005
R53499 VINP.n314 VINP.n97 4.5005
R53500 VINP.n258 VINP.n97 4.5005
R53501 VINP.n316 VINP.n97 4.5005
R53502 VINP.n257 VINP.n97 4.5005
R53503 VINP.n318 VINP.n97 4.5005
R53504 VINP.n256 VINP.n97 4.5005
R53505 VINP.n320 VINP.n97 4.5005
R53506 VINP.n255 VINP.n97 4.5005
R53507 VINP.n322 VINP.n97 4.5005
R53508 VINP.n254 VINP.n97 4.5005
R53509 VINP.n324 VINP.n97 4.5005
R53510 VINP.n253 VINP.n97 4.5005
R53511 VINP.n326 VINP.n97 4.5005
R53512 VINP.n252 VINP.n97 4.5005
R53513 VINP.n328 VINP.n97 4.5005
R53514 VINP.n251 VINP.n97 4.5005
R53515 VINP.n330 VINP.n97 4.5005
R53516 VINP.n250 VINP.n97 4.5005
R53517 VINP.n332 VINP.n97 4.5005
R53518 VINP.n249 VINP.n97 4.5005
R53519 VINP.n334 VINP.n97 4.5005
R53520 VINP.n248 VINP.n97 4.5005
R53521 VINP.n336 VINP.n97 4.5005
R53522 VINP.n247 VINP.n97 4.5005
R53523 VINP.n338 VINP.n97 4.5005
R53524 VINP.n246 VINP.n97 4.5005
R53525 VINP.n340 VINP.n97 4.5005
R53526 VINP.n245 VINP.n97 4.5005
R53527 VINP.n342 VINP.n97 4.5005
R53528 VINP.n244 VINP.n97 4.5005
R53529 VINP.n344 VINP.n97 4.5005
R53530 VINP.n243 VINP.n97 4.5005
R53531 VINP.n346 VINP.n97 4.5005
R53532 VINP.n242 VINP.n97 4.5005
R53533 VINP.n348 VINP.n97 4.5005
R53534 VINP.n241 VINP.n97 4.5005
R53535 VINP.n350 VINP.n97 4.5005
R53536 VINP.n240 VINP.n97 4.5005
R53537 VINP.n352 VINP.n97 4.5005
R53538 VINP.n239 VINP.n97 4.5005
R53539 VINP.n354 VINP.n97 4.5005
R53540 VINP.n238 VINP.n97 4.5005
R53541 VINP.n356 VINP.n97 4.5005
R53542 VINP.n237 VINP.n97 4.5005
R53543 VINP.n358 VINP.n97 4.5005
R53544 VINP.n236 VINP.n97 4.5005
R53545 VINP.n360 VINP.n97 4.5005
R53546 VINP.n235 VINP.n97 4.5005
R53547 VINP.n362 VINP.n97 4.5005
R53548 VINP.n234 VINP.n97 4.5005
R53549 VINP.n364 VINP.n97 4.5005
R53550 VINP.n233 VINP.n97 4.5005
R53551 VINP.n366 VINP.n97 4.5005
R53552 VINP.n232 VINP.n97 4.5005
R53553 VINP.n368 VINP.n97 4.5005
R53554 VINP.n231 VINP.n97 4.5005
R53555 VINP.n370 VINP.n97 4.5005
R53556 VINP.n230 VINP.n97 4.5005
R53557 VINP.n372 VINP.n97 4.5005
R53558 VINP.n229 VINP.n97 4.5005
R53559 VINP.n374 VINP.n97 4.5005
R53560 VINP.n228 VINP.n97 4.5005
R53561 VINP.n376 VINP.n97 4.5005
R53562 VINP.n227 VINP.n97 4.5005
R53563 VINP.n378 VINP.n97 4.5005
R53564 VINP.n226 VINP.n97 4.5005
R53565 VINP.n380 VINP.n97 4.5005
R53566 VINP.n225 VINP.n97 4.5005
R53567 VINP.n382 VINP.n97 4.5005
R53568 VINP.n224 VINP.n97 4.5005
R53569 VINP.n384 VINP.n97 4.5005
R53570 VINP.n223 VINP.n97 4.5005
R53571 VINP.n386 VINP.n97 4.5005
R53572 VINP.n222 VINP.n97 4.5005
R53573 VINP.n388 VINP.n97 4.5005
R53574 VINP.n221 VINP.n97 4.5005
R53575 VINP.n390 VINP.n97 4.5005
R53576 VINP.n220 VINP.n97 4.5005
R53577 VINP.n392 VINP.n97 4.5005
R53578 VINP.n219 VINP.n97 4.5005
R53579 VINP.n394 VINP.n97 4.5005
R53580 VINP.n218 VINP.n97 4.5005
R53581 VINP.n396 VINP.n97 4.5005
R53582 VINP.n217 VINP.n97 4.5005
R53583 VINP.n398 VINP.n97 4.5005
R53584 VINP.n216 VINP.n97 4.5005
R53585 VINP.n400 VINP.n97 4.5005
R53586 VINP.n215 VINP.n97 4.5005
R53587 VINP.n654 VINP.n97 4.5005
R53588 VINP.n656 VINP.n97 4.5005
R53589 VINP.n97 VINP.n0 4.5005
R53590 VINP.n278 VINP.n204 4.5005
R53591 VINP.n276 VINP.n204 4.5005
R53592 VINP.n280 VINP.n204 4.5005
R53593 VINP.n275 VINP.n204 4.5005
R53594 VINP.n282 VINP.n204 4.5005
R53595 VINP.n274 VINP.n204 4.5005
R53596 VINP.n284 VINP.n204 4.5005
R53597 VINP.n273 VINP.n204 4.5005
R53598 VINP.n286 VINP.n204 4.5005
R53599 VINP.n272 VINP.n204 4.5005
R53600 VINP.n288 VINP.n204 4.5005
R53601 VINP.n271 VINP.n204 4.5005
R53602 VINP.n290 VINP.n204 4.5005
R53603 VINP.n270 VINP.n204 4.5005
R53604 VINP.n292 VINP.n204 4.5005
R53605 VINP.n269 VINP.n204 4.5005
R53606 VINP.n294 VINP.n204 4.5005
R53607 VINP.n268 VINP.n204 4.5005
R53608 VINP.n296 VINP.n204 4.5005
R53609 VINP.n267 VINP.n204 4.5005
R53610 VINP.n298 VINP.n204 4.5005
R53611 VINP.n266 VINP.n204 4.5005
R53612 VINP.n300 VINP.n204 4.5005
R53613 VINP.n265 VINP.n204 4.5005
R53614 VINP.n302 VINP.n204 4.5005
R53615 VINP.n264 VINP.n204 4.5005
R53616 VINP.n304 VINP.n204 4.5005
R53617 VINP.n263 VINP.n204 4.5005
R53618 VINP.n306 VINP.n204 4.5005
R53619 VINP.n262 VINP.n204 4.5005
R53620 VINP.n308 VINP.n204 4.5005
R53621 VINP.n261 VINP.n204 4.5005
R53622 VINP.n310 VINP.n204 4.5005
R53623 VINP.n260 VINP.n204 4.5005
R53624 VINP.n312 VINP.n204 4.5005
R53625 VINP.n259 VINP.n204 4.5005
R53626 VINP.n314 VINP.n204 4.5005
R53627 VINP.n258 VINP.n204 4.5005
R53628 VINP.n316 VINP.n204 4.5005
R53629 VINP.n257 VINP.n204 4.5005
R53630 VINP.n318 VINP.n204 4.5005
R53631 VINP.n256 VINP.n204 4.5005
R53632 VINP.n320 VINP.n204 4.5005
R53633 VINP.n255 VINP.n204 4.5005
R53634 VINP.n322 VINP.n204 4.5005
R53635 VINP.n254 VINP.n204 4.5005
R53636 VINP.n324 VINP.n204 4.5005
R53637 VINP.n253 VINP.n204 4.5005
R53638 VINP.n326 VINP.n204 4.5005
R53639 VINP.n252 VINP.n204 4.5005
R53640 VINP.n328 VINP.n204 4.5005
R53641 VINP.n251 VINP.n204 4.5005
R53642 VINP.n330 VINP.n204 4.5005
R53643 VINP.n250 VINP.n204 4.5005
R53644 VINP.n332 VINP.n204 4.5005
R53645 VINP.n249 VINP.n204 4.5005
R53646 VINP.n334 VINP.n204 4.5005
R53647 VINP.n248 VINP.n204 4.5005
R53648 VINP.n336 VINP.n204 4.5005
R53649 VINP.n247 VINP.n204 4.5005
R53650 VINP.n338 VINP.n204 4.5005
R53651 VINP.n246 VINP.n204 4.5005
R53652 VINP.n340 VINP.n204 4.5005
R53653 VINP.n245 VINP.n204 4.5005
R53654 VINP.n342 VINP.n204 4.5005
R53655 VINP.n244 VINP.n204 4.5005
R53656 VINP.n344 VINP.n204 4.5005
R53657 VINP.n243 VINP.n204 4.5005
R53658 VINP.n346 VINP.n204 4.5005
R53659 VINP.n242 VINP.n204 4.5005
R53660 VINP.n348 VINP.n204 4.5005
R53661 VINP.n241 VINP.n204 4.5005
R53662 VINP.n350 VINP.n204 4.5005
R53663 VINP.n240 VINP.n204 4.5005
R53664 VINP.n352 VINP.n204 4.5005
R53665 VINP.n239 VINP.n204 4.5005
R53666 VINP.n354 VINP.n204 4.5005
R53667 VINP.n238 VINP.n204 4.5005
R53668 VINP.n356 VINP.n204 4.5005
R53669 VINP.n237 VINP.n204 4.5005
R53670 VINP.n358 VINP.n204 4.5005
R53671 VINP.n236 VINP.n204 4.5005
R53672 VINP.n360 VINP.n204 4.5005
R53673 VINP.n235 VINP.n204 4.5005
R53674 VINP.n362 VINP.n204 4.5005
R53675 VINP.n234 VINP.n204 4.5005
R53676 VINP.n364 VINP.n204 4.5005
R53677 VINP.n233 VINP.n204 4.5005
R53678 VINP.n366 VINP.n204 4.5005
R53679 VINP.n232 VINP.n204 4.5005
R53680 VINP.n368 VINP.n204 4.5005
R53681 VINP.n231 VINP.n204 4.5005
R53682 VINP.n370 VINP.n204 4.5005
R53683 VINP.n230 VINP.n204 4.5005
R53684 VINP.n372 VINP.n204 4.5005
R53685 VINP.n229 VINP.n204 4.5005
R53686 VINP.n374 VINP.n204 4.5005
R53687 VINP.n228 VINP.n204 4.5005
R53688 VINP.n376 VINP.n204 4.5005
R53689 VINP.n227 VINP.n204 4.5005
R53690 VINP.n378 VINP.n204 4.5005
R53691 VINP.n226 VINP.n204 4.5005
R53692 VINP.n380 VINP.n204 4.5005
R53693 VINP.n225 VINP.n204 4.5005
R53694 VINP.n382 VINP.n204 4.5005
R53695 VINP.n224 VINP.n204 4.5005
R53696 VINP.n384 VINP.n204 4.5005
R53697 VINP.n223 VINP.n204 4.5005
R53698 VINP.n386 VINP.n204 4.5005
R53699 VINP.n222 VINP.n204 4.5005
R53700 VINP.n388 VINP.n204 4.5005
R53701 VINP.n221 VINP.n204 4.5005
R53702 VINP.n390 VINP.n204 4.5005
R53703 VINP.n220 VINP.n204 4.5005
R53704 VINP.n392 VINP.n204 4.5005
R53705 VINP.n219 VINP.n204 4.5005
R53706 VINP.n394 VINP.n204 4.5005
R53707 VINP.n218 VINP.n204 4.5005
R53708 VINP.n396 VINP.n204 4.5005
R53709 VINP.n217 VINP.n204 4.5005
R53710 VINP.n398 VINP.n204 4.5005
R53711 VINP.n216 VINP.n204 4.5005
R53712 VINP.n400 VINP.n204 4.5005
R53713 VINP.n215 VINP.n204 4.5005
R53714 VINP.n654 VINP.n204 4.5005
R53715 VINP.n656 VINP.n204 4.5005
R53716 VINP.n204 VINP.n0 4.5005
R53717 VINP.n278 VINP.n96 4.5005
R53718 VINP.n276 VINP.n96 4.5005
R53719 VINP.n280 VINP.n96 4.5005
R53720 VINP.n275 VINP.n96 4.5005
R53721 VINP.n282 VINP.n96 4.5005
R53722 VINP.n274 VINP.n96 4.5005
R53723 VINP.n284 VINP.n96 4.5005
R53724 VINP.n273 VINP.n96 4.5005
R53725 VINP.n286 VINP.n96 4.5005
R53726 VINP.n272 VINP.n96 4.5005
R53727 VINP.n288 VINP.n96 4.5005
R53728 VINP.n271 VINP.n96 4.5005
R53729 VINP.n290 VINP.n96 4.5005
R53730 VINP.n270 VINP.n96 4.5005
R53731 VINP.n292 VINP.n96 4.5005
R53732 VINP.n269 VINP.n96 4.5005
R53733 VINP.n294 VINP.n96 4.5005
R53734 VINP.n268 VINP.n96 4.5005
R53735 VINP.n296 VINP.n96 4.5005
R53736 VINP.n267 VINP.n96 4.5005
R53737 VINP.n298 VINP.n96 4.5005
R53738 VINP.n266 VINP.n96 4.5005
R53739 VINP.n300 VINP.n96 4.5005
R53740 VINP.n265 VINP.n96 4.5005
R53741 VINP.n302 VINP.n96 4.5005
R53742 VINP.n264 VINP.n96 4.5005
R53743 VINP.n304 VINP.n96 4.5005
R53744 VINP.n263 VINP.n96 4.5005
R53745 VINP.n306 VINP.n96 4.5005
R53746 VINP.n262 VINP.n96 4.5005
R53747 VINP.n308 VINP.n96 4.5005
R53748 VINP.n261 VINP.n96 4.5005
R53749 VINP.n310 VINP.n96 4.5005
R53750 VINP.n260 VINP.n96 4.5005
R53751 VINP.n312 VINP.n96 4.5005
R53752 VINP.n259 VINP.n96 4.5005
R53753 VINP.n314 VINP.n96 4.5005
R53754 VINP.n258 VINP.n96 4.5005
R53755 VINP.n316 VINP.n96 4.5005
R53756 VINP.n257 VINP.n96 4.5005
R53757 VINP.n318 VINP.n96 4.5005
R53758 VINP.n256 VINP.n96 4.5005
R53759 VINP.n320 VINP.n96 4.5005
R53760 VINP.n255 VINP.n96 4.5005
R53761 VINP.n322 VINP.n96 4.5005
R53762 VINP.n254 VINP.n96 4.5005
R53763 VINP.n324 VINP.n96 4.5005
R53764 VINP.n253 VINP.n96 4.5005
R53765 VINP.n326 VINP.n96 4.5005
R53766 VINP.n252 VINP.n96 4.5005
R53767 VINP.n328 VINP.n96 4.5005
R53768 VINP.n251 VINP.n96 4.5005
R53769 VINP.n330 VINP.n96 4.5005
R53770 VINP.n250 VINP.n96 4.5005
R53771 VINP.n332 VINP.n96 4.5005
R53772 VINP.n249 VINP.n96 4.5005
R53773 VINP.n334 VINP.n96 4.5005
R53774 VINP.n248 VINP.n96 4.5005
R53775 VINP.n336 VINP.n96 4.5005
R53776 VINP.n247 VINP.n96 4.5005
R53777 VINP.n338 VINP.n96 4.5005
R53778 VINP.n246 VINP.n96 4.5005
R53779 VINP.n340 VINP.n96 4.5005
R53780 VINP.n245 VINP.n96 4.5005
R53781 VINP.n342 VINP.n96 4.5005
R53782 VINP.n244 VINP.n96 4.5005
R53783 VINP.n344 VINP.n96 4.5005
R53784 VINP.n243 VINP.n96 4.5005
R53785 VINP.n346 VINP.n96 4.5005
R53786 VINP.n242 VINP.n96 4.5005
R53787 VINP.n348 VINP.n96 4.5005
R53788 VINP.n241 VINP.n96 4.5005
R53789 VINP.n350 VINP.n96 4.5005
R53790 VINP.n240 VINP.n96 4.5005
R53791 VINP.n352 VINP.n96 4.5005
R53792 VINP.n239 VINP.n96 4.5005
R53793 VINP.n354 VINP.n96 4.5005
R53794 VINP.n238 VINP.n96 4.5005
R53795 VINP.n356 VINP.n96 4.5005
R53796 VINP.n237 VINP.n96 4.5005
R53797 VINP.n358 VINP.n96 4.5005
R53798 VINP.n236 VINP.n96 4.5005
R53799 VINP.n360 VINP.n96 4.5005
R53800 VINP.n235 VINP.n96 4.5005
R53801 VINP.n362 VINP.n96 4.5005
R53802 VINP.n234 VINP.n96 4.5005
R53803 VINP.n364 VINP.n96 4.5005
R53804 VINP.n233 VINP.n96 4.5005
R53805 VINP.n366 VINP.n96 4.5005
R53806 VINP.n232 VINP.n96 4.5005
R53807 VINP.n368 VINP.n96 4.5005
R53808 VINP.n231 VINP.n96 4.5005
R53809 VINP.n370 VINP.n96 4.5005
R53810 VINP.n230 VINP.n96 4.5005
R53811 VINP.n372 VINP.n96 4.5005
R53812 VINP.n229 VINP.n96 4.5005
R53813 VINP.n374 VINP.n96 4.5005
R53814 VINP.n228 VINP.n96 4.5005
R53815 VINP.n376 VINP.n96 4.5005
R53816 VINP.n227 VINP.n96 4.5005
R53817 VINP.n378 VINP.n96 4.5005
R53818 VINP.n226 VINP.n96 4.5005
R53819 VINP.n380 VINP.n96 4.5005
R53820 VINP.n225 VINP.n96 4.5005
R53821 VINP.n382 VINP.n96 4.5005
R53822 VINP.n224 VINP.n96 4.5005
R53823 VINP.n384 VINP.n96 4.5005
R53824 VINP.n223 VINP.n96 4.5005
R53825 VINP.n386 VINP.n96 4.5005
R53826 VINP.n222 VINP.n96 4.5005
R53827 VINP.n388 VINP.n96 4.5005
R53828 VINP.n221 VINP.n96 4.5005
R53829 VINP.n390 VINP.n96 4.5005
R53830 VINP.n220 VINP.n96 4.5005
R53831 VINP.n392 VINP.n96 4.5005
R53832 VINP.n219 VINP.n96 4.5005
R53833 VINP.n394 VINP.n96 4.5005
R53834 VINP.n218 VINP.n96 4.5005
R53835 VINP.n396 VINP.n96 4.5005
R53836 VINP.n217 VINP.n96 4.5005
R53837 VINP.n398 VINP.n96 4.5005
R53838 VINP.n216 VINP.n96 4.5005
R53839 VINP.n400 VINP.n96 4.5005
R53840 VINP.n215 VINP.n96 4.5005
R53841 VINP.n654 VINP.n96 4.5005
R53842 VINP.n656 VINP.n96 4.5005
R53843 VINP.n96 VINP.n0 4.5005
R53844 VINP.n278 VINP.n205 4.5005
R53845 VINP.n276 VINP.n205 4.5005
R53846 VINP.n280 VINP.n205 4.5005
R53847 VINP.n275 VINP.n205 4.5005
R53848 VINP.n282 VINP.n205 4.5005
R53849 VINP.n274 VINP.n205 4.5005
R53850 VINP.n284 VINP.n205 4.5005
R53851 VINP.n273 VINP.n205 4.5005
R53852 VINP.n286 VINP.n205 4.5005
R53853 VINP.n272 VINP.n205 4.5005
R53854 VINP.n288 VINP.n205 4.5005
R53855 VINP.n271 VINP.n205 4.5005
R53856 VINP.n290 VINP.n205 4.5005
R53857 VINP.n270 VINP.n205 4.5005
R53858 VINP.n292 VINP.n205 4.5005
R53859 VINP.n269 VINP.n205 4.5005
R53860 VINP.n294 VINP.n205 4.5005
R53861 VINP.n268 VINP.n205 4.5005
R53862 VINP.n296 VINP.n205 4.5005
R53863 VINP.n267 VINP.n205 4.5005
R53864 VINP.n298 VINP.n205 4.5005
R53865 VINP.n266 VINP.n205 4.5005
R53866 VINP.n300 VINP.n205 4.5005
R53867 VINP.n265 VINP.n205 4.5005
R53868 VINP.n302 VINP.n205 4.5005
R53869 VINP.n264 VINP.n205 4.5005
R53870 VINP.n304 VINP.n205 4.5005
R53871 VINP.n263 VINP.n205 4.5005
R53872 VINP.n306 VINP.n205 4.5005
R53873 VINP.n262 VINP.n205 4.5005
R53874 VINP.n308 VINP.n205 4.5005
R53875 VINP.n261 VINP.n205 4.5005
R53876 VINP.n310 VINP.n205 4.5005
R53877 VINP.n260 VINP.n205 4.5005
R53878 VINP.n312 VINP.n205 4.5005
R53879 VINP.n259 VINP.n205 4.5005
R53880 VINP.n314 VINP.n205 4.5005
R53881 VINP.n258 VINP.n205 4.5005
R53882 VINP.n316 VINP.n205 4.5005
R53883 VINP.n257 VINP.n205 4.5005
R53884 VINP.n318 VINP.n205 4.5005
R53885 VINP.n256 VINP.n205 4.5005
R53886 VINP.n320 VINP.n205 4.5005
R53887 VINP.n255 VINP.n205 4.5005
R53888 VINP.n322 VINP.n205 4.5005
R53889 VINP.n254 VINP.n205 4.5005
R53890 VINP.n324 VINP.n205 4.5005
R53891 VINP.n253 VINP.n205 4.5005
R53892 VINP.n326 VINP.n205 4.5005
R53893 VINP.n252 VINP.n205 4.5005
R53894 VINP.n328 VINP.n205 4.5005
R53895 VINP.n251 VINP.n205 4.5005
R53896 VINP.n330 VINP.n205 4.5005
R53897 VINP.n250 VINP.n205 4.5005
R53898 VINP.n332 VINP.n205 4.5005
R53899 VINP.n249 VINP.n205 4.5005
R53900 VINP.n334 VINP.n205 4.5005
R53901 VINP.n248 VINP.n205 4.5005
R53902 VINP.n336 VINP.n205 4.5005
R53903 VINP.n247 VINP.n205 4.5005
R53904 VINP.n338 VINP.n205 4.5005
R53905 VINP.n246 VINP.n205 4.5005
R53906 VINP.n340 VINP.n205 4.5005
R53907 VINP.n245 VINP.n205 4.5005
R53908 VINP.n342 VINP.n205 4.5005
R53909 VINP.n244 VINP.n205 4.5005
R53910 VINP.n344 VINP.n205 4.5005
R53911 VINP.n243 VINP.n205 4.5005
R53912 VINP.n346 VINP.n205 4.5005
R53913 VINP.n242 VINP.n205 4.5005
R53914 VINP.n348 VINP.n205 4.5005
R53915 VINP.n241 VINP.n205 4.5005
R53916 VINP.n350 VINP.n205 4.5005
R53917 VINP.n240 VINP.n205 4.5005
R53918 VINP.n352 VINP.n205 4.5005
R53919 VINP.n239 VINP.n205 4.5005
R53920 VINP.n354 VINP.n205 4.5005
R53921 VINP.n238 VINP.n205 4.5005
R53922 VINP.n356 VINP.n205 4.5005
R53923 VINP.n237 VINP.n205 4.5005
R53924 VINP.n358 VINP.n205 4.5005
R53925 VINP.n236 VINP.n205 4.5005
R53926 VINP.n360 VINP.n205 4.5005
R53927 VINP.n235 VINP.n205 4.5005
R53928 VINP.n362 VINP.n205 4.5005
R53929 VINP.n234 VINP.n205 4.5005
R53930 VINP.n364 VINP.n205 4.5005
R53931 VINP.n233 VINP.n205 4.5005
R53932 VINP.n366 VINP.n205 4.5005
R53933 VINP.n232 VINP.n205 4.5005
R53934 VINP.n368 VINP.n205 4.5005
R53935 VINP.n231 VINP.n205 4.5005
R53936 VINP.n370 VINP.n205 4.5005
R53937 VINP.n230 VINP.n205 4.5005
R53938 VINP.n372 VINP.n205 4.5005
R53939 VINP.n229 VINP.n205 4.5005
R53940 VINP.n374 VINP.n205 4.5005
R53941 VINP.n228 VINP.n205 4.5005
R53942 VINP.n376 VINP.n205 4.5005
R53943 VINP.n227 VINP.n205 4.5005
R53944 VINP.n378 VINP.n205 4.5005
R53945 VINP.n226 VINP.n205 4.5005
R53946 VINP.n380 VINP.n205 4.5005
R53947 VINP.n225 VINP.n205 4.5005
R53948 VINP.n382 VINP.n205 4.5005
R53949 VINP.n224 VINP.n205 4.5005
R53950 VINP.n384 VINP.n205 4.5005
R53951 VINP.n223 VINP.n205 4.5005
R53952 VINP.n386 VINP.n205 4.5005
R53953 VINP.n222 VINP.n205 4.5005
R53954 VINP.n388 VINP.n205 4.5005
R53955 VINP.n221 VINP.n205 4.5005
R53956 VINP.n390 VINP.n205 4.5005
R53957 VINP.n220 VINP.n205 4.5005
R53958 VINP.n392 VINP.n205 4.5005
R53959 VINP.n219 VINP.n205 4.5005
R53960 VINP.n394 VINP.n205 4.5005
R53961 VINP.n218 VINP.n205 4.5005
R53962 VINP.n396 VINP.n205 4.5005
R53963 VINP.n217 VINP.n205 4.5005
R53964 VINP.n398 VINP.n205 4.5005
R53965 VINP.n216 VINP.n205 4.5005
R53966 VINP.n400 VINP.n205 4.5005
R53967 VINP.n215 VINP.n205 4.5005
R53968 VINP.n654 VINP.n205 4.5005
R53969 VINP.n656 VINP.n205 4.5005
R53970 VINP.n205 VINP.n0 4.5005
R53971 VINP.n278 VINP.n95 4.5005
R53972 VINP.n276 VINP.n95 4.5005
R53973 VINP.n280 VINP.n95 4.5005
R53974 VINP.n275 VINP.n95 4.5005
R53975 VINP.n282 VINP.n95 4.5005
R53976 VINP.n274 VINP.n95 4.5005
R53977 VINP.n284 VINP.n95 4.5005
R53978 VINP.n273 VINP.n95 4.5005
R53979 VINP.n286 VINP.n95 4.5005
R53980 VINP.n272 VINP.n95 4.5005
R53981 VINP.n288 VINP.n95 4.5005
R53982 VINP.n271 VINP.n95 4.5005
R53983 VINP.n290 VINP.n95 4.5005
R53984 VINP.n270 VINP.n95 4.5005
R53985 VINP.n292 VINP.n95 4.5005
R53986 VINP.n269 VINP.n95 4.5005
R53987 VINP.n294 VINP.n95 4.5005
R53988 VINP.n268 VINP.n95 4.5005
R53989 VINP.n296 VINP.n95 4.5005
R53990 VINP.n267 VINP.n95 4.5005
R53991 VINP.n298 VINP.n95 4.5005
R53992 VINP.n266 VINP.n95 4.5005
R53993 VINP.n300 VINP.n95 4.5005
R53994 VINP.n265 VINP.n95 4.5005
R53995 VINP.n302 VINP.n95 4.5005
R53996 VINP.n264 VINP.n95 4.5005
R53997 VINP.n304 VINP.n95 4.5005
R53998 VINP.n263 VINP.n95 4.5005
R53999 VINP.n306 VINP.n95 4.5005
R54000 VINP.n262 VINP.n95 4.5005
R54001 VINP.n308 VINP.n95 4.5005
R54002 VINP.n261 VINP.n95 4.5005
R54003 VINP.n310 VINP.n95 4.5005
R54004 VINP.n260 VINP.n95 4.5005
R54005 VINP.n312 VINP.n95 4.5005
R54006 VINP.n259 VINP.n95 4.5005
R54007 VINP.n314 VINP.n95 4.5005
R54008 VINP.n258 VINP.n95 4.5005
R54009 VINP.n316 VINP.n95 4.5005
R54010 VINP.n257 VINP.n95 4.5005
R54011 VINP.n318 VINP.n95 4.5005
R54012 VINP.n256 VINP.n95 4.5005
R54013 VINP.n320 VINP.n95 4.5005
R54014 VINP.n255 VINP.n95 4.5005
R54015 VINP.n322 VINP.n95 4.5005
R54016 VINP.n254 VINP.n95 4.5005
R54017 VINP.n324 VINP.n95 4.5005
R54018 VINP.n253 VINP.n95 4.5005
R54019 VINP.n326 VINP.n95 4.5005
R54020 VINP.n252 VINP.n95 4.5005
R54021 VINP.n328 VINP.n95 4.5005
R54022 VINP.n251 VINP.n95 4.5005
R54023 VINP.n330 VINP.n95 4.5005
R54024 VINP.n250 VINP.n95 4.5005
R54025 VINP.n332 VINP.n95 4.5005
R54026 VINP.n249 VINP.n95 4.5005
R54027 VINP.n334 VINP.n95 4.5005
R54028 VINP.n248 VINP.n95 4.5005
R54029 VINP.n336 VINP.n95 4.5005
R54030 VINP.n247 VINP.n95 4.5005
R54031 VINP.n338 VINP.n95 4.5005
R54032 VINP.n246 VINP.n95 4.5005
R54033 VINP.n340 VINP.n95 4.5005
R54034 VINP.n245 VINP.n95 4.5005
R54035 VINP.n342 VINP.n95 4.5005
R54036 VINP.n244 VINP.n95 4.5005
R54037 VINP.n344 VINP.n95 4.5005
R54038 VINP.n243 VINP.n95 4.5005
R54039 VINP.n346 VINP.n95 4.5005
R54040 VINP.n242 VINP.n95 4.5005
R54041 VINP.n348 VINP.n95 4.5005
R54042 VINP.n241 VINP.n95 4.5005
R54043 VINP.n350 VINP.n95 4.5005
R54044 VINP.n240 VINP.n95 4.5005
R54045 VINP.n352 VINP.n95 4.5005
R54046 VINP.n239 VINP.n95 4.5005
R54047 VINP.n354 VINP.n95 4.5005
R54048 VINP.n238 VINP.n95 4.5005
R54049 VINP.n356 VINP.n95 4.5005
R54050 VINP.n237 VINP.n95 4.5005
R54051 VINP.n358 VINP.n95 4.5005
R54052 VINP.n236 VINP.n95 4.5005
R54053 VINP.n360 VINP.n95 4.5005
R54054 VINP.n235 VINP.n95 4.5005
R54055 VINP.n362 VINP.n95 4.5005
R54056 VINP.n234 VINP.n95 4.5005
R54057 VINP.n364 VINP.n95 4.5005
R54058 VINP.n233 VINP.n95 4.5005
R54059 VINP.n366 VINP.n95 4.5005
R54060 VINP.n232 VINP.n95 4.5005
R54061 VINP.n368 VINP.n95 4.5005
R54062 VINP.n231 VINP.n95 4.5005
R54063 VINP.n370 VINP.n95 4.5005
R54064 VINP.n230 VINP.n95 4.5005
R54065 VINP.n372 VINP.n95 4.5005
R54066 VINP.n229 VINP.n95 4.5005
R54067 VINP.n374 VINP.n95 4.5005
R54068 VINP.n228 VINP.n95 4.5005
R54069 VINP.n376 VINP.n95 4.5005
R54070 VINP.n227 VINP.n95 4.5005
R54071 VINP.n378 VINP.n95 4.5005
R54072 VINP.n226 VINP.n95 4.5005
R54073 VINP.n380 VINP.n95 4.5005
R54074 VINP.n225 VINP.n95 4.5005
R54075 VINP.n382 VINP.n95 4.5005
R54076 VINP.n224 VINP.n95 4.5005
R54077 VINP.n384 VINP.n95 4.5005
R54078 VINP.n223 VINP.n95 4.5005
R54079 VINP.n386 VINP.n95 4.5005
R54080 VINP.n222 VINP.n95 4.5005
R54081 VINP.n388 VINP.n95 4.5005
R54082 VINP.n221 VINP.n95 4.5005
R54083 VINP.n390 VINP.n95 4.5005
R54084 VINP.n220 VINP.n95 4.5005
R54085 VINP.n392 VINP.n95 4.5005
R54086 VINP.n219 VINP.n95 4.5005
R54087 VINP.n394 VINP.n95 4.5005
R54088 VINP.n218 VINP.n95 4.5005
R54089 VINP.n396 VINP.n95 4.5005
R54090 VINP.n217 VINP.n95 4.5005
R54091 VINP.n398 VINP.n95 4.5005
R54092 VINP.n216 VINP.n95 4.5005
R54093 VINP.n400 VINP.n95 4.5005
R54094 VINP.n215 VINP.n95 4.5005
R54095 VINP.n654 VINP.n95 4.5005
R54096 VINP.n656 VINP.n95 4.5005
R54097 VINP.n95 VINP.n0 4.5005
R54098 VINP.n278 VINP.n206 4.5005
R54099 VINP.n276 VINP.n206 4.5005
R54100 VINP.n280 VINP.n206 4.5005
R54101 VINP.n275 VINP.n206 4.5005
R54102 VINP.n282 VINP.n206 4.5005
R54103 VINP.n274 VINP.n206 4.5005
R54104 VINP.n284 VINP.n206 4.5005
R54105 VINP.n273 VINP.n206 4.5005
R54106 VINP.n286 VINP.n206 4.5005
R54107 VINP.n272 VINP.n206 4.5005
R54108 VINP.n288 VINP.n206 4.5005
R54109 VINP.n271 VINP.n206 4.5005
R54110 VINP.n290 VINP.n206 4.5005
R54111 VINP.n270 VINP.n206 4.5005
R54112 VINP.n292 VINP.n206 4.5005
R54113 VINP.n269 VINP.n206 4.5005
R54114 VINP.n294 VINP.n206 4.5005
R54115 VINP.n268 VINP.n206 4.5005
R54116 VINP.n296 VINP.n206 4.5005
R54117 VINP.n267 VINP.n206 4.5005
R54118 VINP.n298 VINP.n206 4.5005
R54119 VINP.n266 VINP.n206 4.5005
R54120 VINP.n300 VINP.n206 4.5005
R54121 VINP.n265 VINP.n206 4.5005
R54122 VINP.n302 VINP.n206 4.5005
R54123 VINP.n264 VINP.n206 4.5005
R54124 VINP.n304 VINP.n206 4.5005
R54125 VINP.n263 VINP.n206 4.5005
R54126 VINP.n306 VINP.n206 4.5005
R54127 VINP.n262 VINP.n206 4.5005
R54128 VINP.n308 VINP.n206 4.5005
R54129 VINP.n261 VINP.n206 4.5005
R54130 VINP.n310 VINP.n206 4.5005
R54131 VINP.n260 VINP.n206 4.5005
R54132 VINP.n312 VINP.n206 4.5005
R54133 VINP.n259 VINP.n206 4.5005
R54134 VINP.n314 VINP.n206 4.5005
R54135 VINP.n258 VINP.n206 4.5005
R54136 VINP.n316 VINP.n206 4.5005
R54137 VINP.n257 VINP.n206 4.5005
R54138 VINP.n318 VINP.n206 4.5005
R54139 VINP.n256 VINP.n206 4.5005
R54140 VINP.n320 VINP.n206 4.5005
R54141 VINP.n255 VINP.n206 4.5005
R54142 VINP.n322 VINP.n206 4.5005
R54143 VINP.n254 VINP.n206 4.5005
R54144 VINP.n324 VINP.n206 4.5005
R54145 VINP.n253 VINP.n206 4.5005
R54146 VINP.n326 VINP.n206 4.5005
R54147 VINP.n252 VINP.n206 4.5005
R54148 VINP.n328 VINP.n206 4.5005
R54149 VINP.n251 VINP.n206 4.5005
R54150 VINP.n330 VINP.n206 4.5005
R54151 VINP.n250 VINP.n206 4.5005
R54152 VINP.n332 VINP.n206 4.5005
R54153 VINP.n249 VINP.n206 4.5005
R54154 VINP.n334 VINP.n206 4.5005
R54155 VINP.n248 VINP.n206 4.5005
R54156 VINP.n336 VINP.n206 4.5005
R54157 VINP.n247 VINP.n206 4.5005
R54158 VINP.n338 VINP.n206 4.5005
R54159 VINP.n246 VINP.n206 4.5005
R54160 VINP.n340 VINP.n206 4.5005
R54161 VINP.n245 VINP.n206 4.5005
R54162 VINP.n342 VINP.n206 4.5005
R54163 VINP.n244 VINP.n206 4.5005
R54164 VINP.n344 VINP.n206 4.5005
R54165 VINP.n243 VINP.n206 4.5005
R54166 VINP.n346 VINP.n206 4.5005
R54167 VINP.n242 VINP.n206 4.5005
R54168 VINP.n348 VINP.n206 4.5005
R54169 VINP.n241 VINP.n206 4.5005
R54170 VINP.n350 VINP.n206 4.5005
R54171 VINP.n240 VINP.n206 4.5005
R54172 VINP.n352 VINP.n206 4.5005
R54173 VINP.n239 VINP.n206 4.5005
R54174 VINP.n354 VINP.n206 4.5005
R54175 VINP.n238 VINP.n206 4.5005
R54176 VINP.n356 VINP.n206 4.5005
R54177 VINP.n237 VINP.n206 4.5005
R54178 VINP.n358 VINP.n206 4.5005
R54179 VINP.n236 VINP.n206 4.5005
R54180 VINP.n360 VINP.n206 4.5005
R54181 VINP.n235 VINP.n206 4.5005
R54182 VINP.n362 VINP.n206 4.5005
R54183 VINP.n234 VINP.n206 4.5005
R54184 VINP.n364 VINP.n206 4.5005
R54185 VINP.n233 VINP.n206 4.5005
R54186 VINP.n366 VINP.n206 4.5005
R54187 VINP.n232 VINP.n206 4.5005
R54188 VINP.n368 VINP.n206 4.5005
R54189 VINP.n231 VINP.n206 4.5005
R54190 VINP.n370 VINP.n206 4.5005
R54191 VINP.n230 VINP.n206 4.5005
R54192 VINP.n372 VINP.n206 4.5005
R54193 VINP.n229 VINP.n206 4.5005
R54194 VINP.n374 VINP.n206 4.5005
R54195 VINP.n228 VINP.n206 4.5005
R54196 VINP.n376 VINP.n206 4.5005
R54197 VINP.n227 VINP.n206 4.5005
R54198 VINP.n378 VINP.n206 4.5005
R54199 VINP.n226 VINP.n206 4.5005
R54200 VINP.n380 VINP.n206 4.5005
R54201 VINP.n225 VINP.n206 4.5005
R54202 VINP.n382 VINP.n206 4.5005
R54203 VINP.n224 VINP.n206 4.5005
R54204 VINP.n384 VINP.n206 4.5005
R54205 VINP.n223 VINP.n206 4.5005
R54206 VINP.n386 VINP.n206 4.5005
R54207 VINP.n222 VINP.n206 4.5005
R54208 VINP.n388 VINP.n206 4.5005
R54209 VINP.n221 VINP.n206 4.5005
R54210 VINP.n390 VINP.n206 4.5005
R54211 VINP.n220 VINP.n206 4.5005
R54212 VINP.n392 VINP.n206 4.5005
R54213 VINP.n219 VINP.n206 4.5005
R54214 VINP.n394 VINP.n206 4.5005
R54215 VINP.n218 VINP.n206 4.5005
R54216 VINP.n396 VINP.n206 4.5005
R54217 VINP.n217 VINP.n206 4.5005
R54218 VINP.n398 VINP.n206 4.5005
R54219 VINP.n216 VINP.n206 4.5005
R54220 VINP.n400 VINP.n206 4.5005
R54221 VINP.n215 VINP.n206 4.5005
R54222 VINP.n654 VINP.n206 4.5005
R54223 VINP.n656 VINP.n206 4.5005
R54224 VINP.n206 VINP.n0 4.5005
R54225 VINP.n278 VINP.n94 4.5005
R54226 VINP.n276 VINP.n94 4.5005
R54227 VINP.n280 VINP.n94 4.5005
R54228 VINP.n275 VINP.n94 4.5005
R54229 VINP.n282 VINP.n94 4.5005
R54230 VINP.n274 VINP.n94 4.5005
R54231 VINP.n284 VINP.n94 4.5005
R54232 VINP.n273 VINP.n94 4.5005
R54233 VINP.n286 VINP.n94 4.5005
R54234 VINP.n272 VINP.n94 4.5005
R54235 VINP.n288 VINP.n94 4.5005
R54236 VINP.n271 VINP.n94 4.5005
R54237 VINP.n290 VINP.n94 4.5005
R54238 VINP.n270 VINP.n94 4.5005
R54239 VINP.n292 VINP.n94 4.5005
R54240 VINP.n269 VINP.n94 4.5005
R54241 VINP.n294 VINP.n94 4.5005
R54242 VINP.n268 VINP.n94 4.5005
R54243 VINP.n296 VINP.n94 4.5005
R54244 VINP.n267 VINP.n94 4.5005
R54245 VINP.n298 VINP.n94 4.5005
R54246 VINP.n266 VINP.n94 4.5005
R54247 VINP.n300 VINP.n94 4.5005
R54248 VINP.n265 VINP.n94 4.5005
R54249 VINP.n302 VINP.n94 4.5005
R54250 VINP.n264 VINP.n94 4.5005
R54251 VINP.n304 VINP.n94 4.5005
R54252 VINP.n263 VINP.n94 4.5005
R54253 VINP.n306 VINP.n94 4.5005
R54254 VINP.n262 VINP.n94 4.5005
R54255 VINP.n308 VINP.n94 4.5005
R54256 VINP.n261 VINP.n94 4.5005
R54257 VINP.n310 VINP.n94 4.5005
R54258 VINP.n260 VINP.n94 4.5005
R54259 VINP.n312 VINP.n94 4.5005
R54260 VINP.n259 VINP.n94 4.5005
R54261 VINP.n314 VINP.n94 4.5005
R54262 VINP.n258 VINP.n94 4.5005
R54263 VINP.n316 VINP.n94 4.5005
R54264 VINP.n257 VINP.n94 4.5005
R54265 VINP.n318 VINP.n94 4.5005
R54266 VINP.n256 VINP.n94 4.5005
R54267 VINP.n320 VINP.n94 4.5005
R54268 VINP.n255 VINP.n94 4.5005
R54269 VINP.n322 VINP.n94 4.5005
R54270 VINP.n254 VINP.n94 4.5005
R54271 VINP.n324 VINP.n94 4.5005
R54272 VINP.n253 VINP.n94 4.5005
R54273 VINP.n326 VINP.n94 4.5005
R54274 VINP.n252 VINP.n94 4.5005
R54275 VINP.n328 VINP.n94 4.5005
R54276 VINP.n251 VINP.n94 4.5005
R54277 VINP.n330 VINP.n94 4.5005
R54278 VINP.n250 VINP.n94 4.5005
R54279 VINP.n332 VINP.n94 4.5005
R54280 VINP.n249 VINP.n94 4.5005
R54281 VINP.n334 VINP.n94 4.5005
R54282 VINP.n248 VINP.n94 4.5005
R54283 VINP.n336 VINP.n94 4.5005
R54284 VINP.n247 VINP.n94 4.5005
R54285 VINP.n338 VINP.n94 4.5005
R54286 VINP.n246 VINP.n94 4.5005
R54287 VINP.n340 VINP.n94 4.5005
R54288 VINP.n245 VINP.n94 4.5005
R54289 VINP.n342 VINP.n94 4.5005
R54290 VINP.n244 VINP.n94 4.5005
R54291 VINP.n344 VINP.n94 4.5005
R54292 VINP.n243 VINP.n94 4.5005
R54293 VINP.n346 VINP.n94 4.5005
R54294 VINP.n242 VINP.n94 4.5005
R54295 VINP.n348 VINP.n94 4.5005
R54296 VINP.n241 VINP.n94 4.5005
R54297 VINP.n350 VINP.n94 4.5005
R54298 VINP.n240 VINP.n94 4.5005
R54299 VINP.n352 VINP.n94 4.5005
R54300 VINP.n239 VINP.n94 4.5005
R54301 VINP.n354 VINP.n94 4.5005
R54302 VINP.n238 VINP.n94 4.5005
R54303 VINP.n356 VINP.n94 4.5005
R54304 VINP.n237 VINP.n94 4.5005
R54305 VINP.n358 VINP.n94 4.5005
R54306 VINP.n236 VINP.n94 4.5005
R54307 VINP.n360 VINP.n94 4.5005
R54308 VINP.n235 VINP.n94 4.5005
R54309 VINP.n362 VINP.n94 4.5005
R54310 VINP.n234 VINP.n94 4.5005
R54311 VINP.n364 VINP.n94 4.5005
R54312 VINP.n233 VINP.n94 4.5005
R54313 VINP.n366 VINP.n94 4.5005
R54314 VINP.n232 VINP.n94 4.5005
R54315 VINP.n368 VINP.n94 4.5005
R54316 VINP.n231 VINP.n94 4.5005
R54317 VINP.n370 VINP.n94 4.5005
R54318 VINP.n230 VINP.n94 4.5005
R54319 VINP.n372 VINP.n94 4.5005
R54320 VINP.n229 VINP.n94 4.5005
R54321 VINP.n374 VINP.n94 4.5005
R54322 VINP.n228 VINP.n94 4.5005
R54323 VINP.n376 VINP.n94 4.5005
R54324 VINP.n227 VINP.n94 4.5005
R54325 VINP.n378 VINP.n94 4.5005
R54326 VINP.n226 VINP.n94 4.5005
R54327 VINP.n380 VINP.n94 4.5005
R54328 VINP.n225 VINP.n94 4.5005
R54329 VINP.n382 VINP.n94 4.5005
R54330 VINP.n224 VINP.n94 4.5005
R54331 VINP.n384 VINP.n94 4.5005
R54332 VINP.n223 VINP.n94 4.5005
R54333 VINP.n386 VINP.n94 4.5005
R54334 VINP.n222 VINP.n94 4.5005
R54335 VINP.n388 VINP.n94 4.5005
R54336 VINP.n221 VINP.n94 4.5005
R54337 VINP.n390 VINP.n94 4.5005
R54338 VINP.n220 VINP.n94 4.5005
R54339 VINP.n392 VINP.n94 4.5005
R54340 VINP.n219 VINP.n94 4.5005
R54341 VINP.n394 VINP.n94 4.5005
R54342 VINP.n218 VINP.n94 4.5005
R54343 VINP.n396 VINP.n94 4.5005
R54344 VINP.n217 VINP.n94 4.5005
R54345 VINP.n398 VINP.n94 4.5005
R54346 VINP.n216 VINP.n94 4.5005
R54347 VINP.n400 VINP.n94 4.5005
R54348 VINP.n215 VINP.n94 4.5005
R54349 VINP.n654 VINP.n94 4.5005
R54350 VINP.n656 VINP.n94 4.5005
R54351 VINP.n94 VINP.n0 4.5005
R54352 VINP.n278 VINP.n207 4.5005
R54353 VINP.n276 VINP.n207 4.5005
R54354 VINP.n280 VINP.n207 4.5005
R54355 VINP.n275 VINP.n207 4.5005
R54356 VINP.n282 VINP.n207 4.5005
R54357 VINP.n274 VINP.n207 4.5005
R54358 VINP.n284 VINP.n207 4.5005
R54359 VINP.n273 VINP.n207 4.5005
R54360 VINP.n286 VINP.n207 4.5005
R54361 VINP.n272 VINP.n207 4.5005
R54362 VINP.n288 VINP.n207 4.5005
R54363 VINP.n271 VINP.n207 4.5005
R54364 VINP.n290 VINP.n207 4.5005
R54365 VINP.n270 VINP.n207 4.5005
R54366 VINP.n292 VINP.n207 4.5005
R54367 VINP.n269 VINP.n207 4.5005
R54368 VINP.n294 VINP.n207 4.5005
R54369 VINP.n268 VINP.n207 4.5005
R54370 VINP.n296 VINP.n207 4.5005
R54371 VINP.n267 VINP.n207 4.5005
R54372 VINP.n298 VINP.n207 4.5005
R54373 VINP.n266 VINP.n207 4.5005
R54374 VINP.n300 VINP.n207 4.5005
R54375 VINP.n265 VINP.n207 4.5005
R54376 VINP.n302 VINP.n207 4.5005
R54377 VINP.n264 VINP.n207 4.5005
R54378 VINP.n304 VINP.n207 4.5005
R54379 VINP.n263 VINP.n207 4.5005
R54380 VINP.n306 VINP.n207 4.5005
R54381 VINP.n262 VINP.n207 4.5005
R54382 VINP.n308 VINP.n207 4.5005
R54383 VINP.n261 VINP.n207 4.5005
R54384 VINP.n310 VINP.n207 4.5005
R54385 VINP.n260 VINP.n207 4.5005
R54386 VINP.n312 VINP.n207 4.5005
R54387 VINP.n259 VINP.n207 4.5005
R54388 VINP.n314 VINP.n207 4.5005
R54389 VINP.n258 VINP.n207 4.5005
R54390 VINP.n316 VINP.n207 4.5005
R54391 VINP.n257 VINP.n207 4.5005
R54392 VINP.n318 VINP.n207 4.5005
R54393 VINP.n256 VINP.n207 4.5005
R54394 VINP.n320 VINP.n207 4.5005
R54395 VINP.n255 VINP.n207 4.5005
R54396 VINP.n322 VINP.n207 4.5005
R54397 VINP.n254 VINP.n207 4.5005
R54398 VINP.n324 VINP.n207 4.5005
R54399 VINP.n253 VINP.n207 4.5005
R54400 VINP.n326 VINP.n207 4.5005
R54401 VINP.n252 VINP.n207 4.5005
R54402 VINP.n328 VINP.n207 4.5005
R54403 VINP.n251 VINP.n207 4.5005
R54404 VINP.n330 VINP.n207 4.5005
R54405 VINP.n250 VINP.n207 4.5005
R54406 VINP.n332 VINP.n207 4.5005
R54407 VINP.n249 VINP.n207 4.5005
R54408 VINP.n334 VINP.n207 4.5005
R54409 VINP.n248 VINP.n207 4.5005
R54410 VINP.n336 VINP.n207 4.5005
R54411 VINP.n247 VINP.n207 4.5005
R54412 VINP.n338 VINP.n207 4.5005
R54413 VINP.n246 VINP.n207 4.5005
R54414 VINP.n340 VINP.n207 4.5005
R54415 VINP.n245 VINP.n207 4.5005
R54416 VINP.n342 VINP.n207 4.5005
R54417 VINP.n244 VINP.n207 4.5005
R54418 VINP.n344 VINP.n207 4.5005
R54419 VINP.n243 VINP.n207 4.5005
R54420 VINP.n346 VINP.n207 4.5005
R54421 VINP.n242 VINP.n207 4.5005
R54422 VINP.n348 VINP.n207 4.5005
R54423 VINP.n241 VINP.n207 4.5005
R54424 VINP.n350 VINP.n207 4.5005
R54425 VINP.n240 VINP.n207 4.5005
R54426 VINP.n352 VINP.n207 4.5005
R54427 VINP.n239 VINP.n207 4.5005
R54428 VINP.n354 VINP.n207 4.5005
R54429 VINP.n238 VINP.n207 4.5005
R54430 VINP.n356 VINP.n207 4.5005
R54431 VINP.n237 VINP.n207 4.5005
R54432 VINP.n358 VINP.n207 4.5005
R54433 VINP.n236 VINP.n207 4.5005
R54434 VINP.n360 VINP.n207 4.5005
R54435 VINP.n235 VINP.n207 4.5005
R54436 VINP.n362 VINP.n207 4.5005
R54437 VINP.n234 VINP.n207 4.5005
R54438 VINP.n364 VINP.n207 4.5005
R54439 VINP.n233 VINP.n207 4.5005
R54440 VINP.n366 VINP.n207 4.5005
R54441 VINP.n232 VINP.n207 4.5005
R54442 VINP.n368 VINP.n207 4.5005
R54443 VINP.n231 VINP.n207 4.5005
R54444 VINP.n370 VINP.n207 4.5005
R54445 VINP.n230 VINP.n207 4.5005
R54446 VINP.n372 VINP.n207 4.5005
R54447 VINP.n229 VINP.n207 4.5005
R54448 VINP.n374 VINP.n207 4.5005
R54449 VINP.n228 VINP.n207 4.5005
R54450 VINP.n376 VINP.n207 4.5005
R54451 VINP.n227 VINP.n207 4.5005
R54452 VINP.n378 VINP.n207 4.5005
R54453 VINP.n226 VINP.n207 4.5005
R54454 VINP.n380 VINP.n207 4.5005
R54455 VINP.n225 VINP.n207 4.5005
R54456 VINP.n382 VINP.n207 4.5005
R54457 VINP.n224 VINP.n207 4.5005
R54458 VINP.n384 VINP.n207 4.5005
R54459 VINP.n223 VINP.n207 4.5005
R54460 VINP.n386 VINP.n207 4.5005
R54461 VINP.n222 VINP.n207 4.5005
R54462 VINP.n388 VINP.n207 4.5005
R54463 VINP.n221 VINP.n207 4.5005
R54464 VINP.n390 VINP.n207 4.5005
R54465 VINP.n220 VINP.n207 4.5005
R54466 VINP.n392 VINP.n207 4.5005
R54467 VINP.n219 VINP.n207 4.5005
R54468 VINP.n394 VINP.n207 4.5005
R54469 VINP.n218 VINP.n207 4.5005
R54470 VINP.n396 VINP.n207 4.5005
R54471 VINP.n217 VINP.n207 4.5005
R54472 VINP.n398 VINP.n207 4.5005
R54473 VINP.n216 VINP.n207 4.5005
R54474 VINP.n400 VINP.n207 4.5005
R54475 VINP.n215 VINP.n207 4.5005
R54476 VINP.n654 VINP.n207 4.5005
R54477 VINP.n656 VINP.n207 4.5005
R54478 VINP.n207 VINP.n0 4.5005
R54479 VINP.n278 VINP.n93 4.5005
R54480 VINP.n276 VINP.n93 4.5005
R54481 VINP.n280 VINP.n93 4.5005
R54482 VINP.n275 VINP.n93 4.5005
R54483 VINP.n282 VINP.n93 4.5005
R54484 VINP.n274 VINP.n93 4.5005
R54485 VINP.n284 VINP.n93 4.5005
R54486 VINP.n273 VINP.n93 4.5005
R54487 VINP.n286 VINP.n93 4.5005
R54488 VINP.n272 VINP.n93 4.5005
R54489 VINP.n288 VINP.n93 4.5005
R54490 VINP.n271 VINP.n93 4.5005
R54491 VINP.n290 VINP.n93 4.5005
R54492 VINP.n270 VINP.n93 4.5005
R54493 VINP.n292 VINP.n93 4.5005
R54494 VINP.n269 VINP.n93 4.5005
R54495 VINP.n294 VINP.n93 4.5005
R54496 VINP.n268 VINP.n93 4.5005
R54497 VINP.n296 VINP.n93 4.5005
R54498 VINP.n267 VINP.n93 4.5005
R54499 VINP.n298 VINP.n93 4.5005
R54500 VINP.n266 VINP.n93 4.5005
R54501 VINP.n300 VINP.n93 4.5005
R54502 VINP.n265 VINP.n93 4.5005
R54503 VINP.n302 VINP.n93 4.5005
R54504 VINP.n264 VINP.n93 4.5005
R54505 VINP.n304 VINP.n93 4.5005
R54506 VINP.n263 VINP.n93 4.5005
R54507 VINP.n306 VINP.n93 4.5005
R54508 VINP.n262 VINP.n93 4.5005
R54509 VINP.n308 VINP.n93 4.5005
R54510 VINP.n261 VINP.n93 4.5005
R54511 VINP.n310 VINP.n93 4.5005
R54512 VINP.n260 VINP.n93 4.5005
R54513 VINP.n312 VINP.n93 4.5005
R54514 VINP.n259 VINP.n93 4.5005
R54515 VINP.n314 VINP.n93 4.5005
R54516 VINP.n258 VINP.n93 4.5005
R54517 VINP.n316 VINP.n93 4.5005
R54518 VINP.n257 VINP.n93 4.5005
R54519 VINP.n318 VINP.n93 4.5005
R54520 VINP.n256 VINP.n93 4.5005
R54521 VINP.n320 VINP.n93 4.5005
R54522 VINP.n255 VINP.n93 4.5005
R54523 VINP.n322 VINP.n93 4.5005
R54524 VINP.n254 VINP.n93 4.5005
R54525 VINP.n324 VINP.n93 4.5005
R54526 VINP.n253 VINP.n93 4.5005
R54527 VINP.n326 VINP.n93 4.5005
R54528 VINP.n252 VINP.n93 4.5005
R54529 VINP.n328 VINP.n93 4.5005
R54530 VINP.n251 VINP.n93 4.5005
R54531 VINP.n330 VINP.n93 4.5005
R54532 VINP.n250 VINP.n93 4.5005
R54533 VINP.n332 VINP.n93 4.5005
R54534 VINP.n249 VINP.n93 4.5005
R54535 VINP.n334 VINP.n93 4.5005
R54536 VINP.n248 VINP.n93 4.5005
R54537 VINP.n336 VINP.n93 4.5005
R54538 VINP.n247 VINP.n93 4.5005
R54539 VINP.n338 VINP.n93 4.5005
R54540 VINP.n246 VINP.n93 4.5005
R54541 VINP.n340 VINP.n93 4.5005
R54542 VINP.n245 VINP.n93 4.5005
R54543 VINP.n342 VINP.n93 4.5005
R54544 VINP.n244 VINP.n93 4.5005
R54545 VINP.n344 VINP.n93 4.5005
R54546 VINP.n243 VINP.n93 4.5005
R54547 VINP.n346 VINP.n93 4.5005
R54548 VINP.n242 VINP.n93 4.5005
R54549 VINP.n348 VINP.n93 4.5005
R54550 VINP.n241 VINP.n93 4.5005
R54551 VINP.n350 VINP.n93 4.5005
R54552 VINP.n240 VINP.n93 4.5005
R54553 VINP.n352 VINP.n93 4.5005
R54554 VINP.n239 VINP.n93 4.5005
R54555 VINP.n354 VINP.n93 4.5005
R54556 VINP.n238 VINP.n93 4.5005
R54557 VINP.n356 VINP.n93 4.5005
R54558 VINP.n237 VINP.n93 4.5005
R54559 VINP.n358 VINP.n93 4.5005
R54560 VINP.n236 VINP.n93 4.5005
R54561 VINP.n360 VINP.n93 4.5005
R54562 VINP.n235 VINP.n93 4.5005
R54563 VINP.n362 VINP.n93 4.5005
R54564 VINP.n234 VINP.n93 4.5005
R54565 VINP.n364 VINP.n93 4.5005
R54566 VINP.n233 VINP.n93 4.5005
R54567 VINP.n366 VINP.n93 4.5005
R54568 VINP.n232 VINP.n93 4.5005
R54569 VINP.n368 VINP.n93 4.5005
R54570 VINP.n231 VINP.n93 4.5005
R54571 VINP.n370 VINP.n93 4.5005
R54572 VINP.n230 VINP.n93 4.5005
R54573 VINP.n372 VINP.n93 4.5005
R54574 VINP.n229 VINP.n93 4.5005
R54575 VINP.n374 VINP.n93 4.5005
R54576 VINP.n228 VINP.n93 4.5005
R54577 VINP.n376 VINP.n93 4.5005
R54578 VINP.n227 VINP.n93 4.5005
R54579 VINP.n378 VINP.n93 4.5005
R54580 VINP.n226 VINP.n93 4.5005
R54581 VINP.n380 VINP.n93 4.5005
R54582 VINP.n225 VINP.n93 4.5005
R54583 VINP.n382 VINP.n93 4.5005
R54584 VINP.n224 VINP.n93 4.5005
R54585 VINP.n384 VINP.n93 4.5005
R54586 VINP.n223 VINP.n93 4.5005
R54587 VINP.n386 VINP.n93 4.5005
R54588 VINP.n222 VINP.n93 4.5005
R54589 VINP.n388 VINP.n93 4.5005
R54590 VINP.n221 VINP.n93 4.5005
R54591 VINP.n390 VINP.n93 4.5005
R54592 VINP.n220 VINP.n93 4.5005
R54593 VINP.n392 VINP.n93 4.5005
R54594 VINP.n219 VINP.n93 4.5005
R54595 VINP.n394 VINP.n93 4.5005
R54596 VINP.n218 VINP.n93 4.5005
R54597 VINP.n396 VINP.n93 4.5005
R54598 VINP.n217 VINP.n93 4.5005
R54599 VINP.n398 VINP.n93 4.5005
R54600 VINP.n216 VINP.n93 4.5005
R54601 VINP.n400 VINP.n93 4.5005
R54602 VINP.n215 VINP.n93 4.5005
R54603 VINP.n654 VINP.n93 4.5005
R54604 VINP.n656 VINP.n93 4.5005
R54605 VINP.n93 VINP.n0 4.5005
R54606 VINP.n278 VINP.n208 4.5005
R54607 VINP.n276 VINP.n208 4.5005
R54608 VINP.n280 VINP.n208 4.5005
R54609 VINP.n275 VINP.n208 4.5005
R54610 VINP.n282 VINP.n208 4.5005
R54611 VINP.n274 VINP.n208 4.5005
R54612 VINP.n284 VINP.n208 4.5005
R54613 VINP.n273 VINP.n208 4.5005
R54614 VINP.n286 VINP.n208 4.5005
R54615 VINP.n272 VINP.n208 4.5005
R54616 VINP.n288 VINP.n208 4.5005
R54617 VINP.n271 VINP.n208 4.5005
R54618 VINP.n290 VINP.n208 4.5005
R54619 VINP.n270 VINP.n208 4.5005
R54620 VINP.n292 VINP.n208 4.5005
R54621 VINP.n269 VINP.n208 4.5005
R54622 VINP.n294 VINP.n208 4.5005
R54623 VINP.n268 VINP.n208 4.5005
R54624 VINP.n296 VINP.n208 4.5005
R54625 VINP.n267 VINP.n208 4.5005
R54626 VINP.n298 VINP.n208 4.5005
R54627 VINP.n266 VINP.n208 4.5005
R54628 VINP.n300 VINP.n208 4.5005
R54629 VINP.n265 VINP.n208 4.5005
R54630 VINP.n302 VINP.n208 4.5005
R54631 VINP.n264 VINP.n208 4.5005
R54632 VINP.n304 VINP.n208 4.5005
R54633 VINP.n263 VINP.n208 4.5005
R54634 VINP.n306 VINP.n208 4.5005
R54635 VINP.n262 VINP.n208 4.5005
R54636 VINP.n308 VINP.n208 4.5005
R54637 VINP.n261 VINP.n208 4.5005
R54638 VINP.n310 VINP.n208 4.5005
R54639 VINP.n260 VINP.n208 4.5005
R54640 VINP.n312 VINP.n208 4.5005
R54641 VINP.n259 VINP.n208 4.5005
R54642 VINP.n314 VINP.n208 4.5005
R54643 VINP.n258 VINP.n208 4.5005
R54644 VINP.n316 VINP.n208 4.5005
R54645 VINP.n257 VINP.n208 4.5005
R54646 VINP.n318 VINP.n208 4.5005
R54647 VINP.n256 VINP.n208 4.5005
R54648 VINP.n320 VINP.n208 4.5005
R54649 VINP.n255 VINP.n208 4.5005
R54650 VINP.n322 VINP.n208 4.5005
R54651 VINP.n254 VINP.n208 4.5005
R54652 VINP.n324 VINP.n208 4.5005
R54653 VINP.n253 VINP.n208 4.5005
R54654 VINP.n326 VINP.n208 4.5005
R54655 VINP.n252 VINP.n208 4.5005
R54656 VINP.n328 VINP.n208 4.5005
R54657 VINP.n251 VINP.n208 4.5005
R54658 VINP.n330 VINP.n208 4.5005
R54659 VINP.n250 VINP.n208 4.5005
R54660 VINP.n332 VINP.n208 4.5005
R54661 VINP.n249 VINP.n208 4.5005
R54662 VINP.n334 VINP.n208 4.5005
R54663 VINP.n248 VINP.n208 4.5005
R54664 VINP.n336 VINP.n208 4.5005
R54665 VINP.n247 VINP.n208 4.5005
R54666 VINP.n338 VINP.n208 4.5005
R54667 VINP.n246 VINP.n208 4.5005
R54668 VINP.n340 VINP.n208 4.5005
R54669 VINP.n245 VINP.n208 4.5005
R54670 VINP.n342 VINP.n208 4.5005
R54671 VINP.n244 VINP.n208 4.5005
R54672 VINP.n344 VINP.n208 4.5005
R54673 VINP.n243 VINP.n208 4.5005
R54674 VINP.n346 VINP.n208 4.5005
R54675 VINP.n242 VINP.n208 4.5005
R54676 VINP.n348 VINP.n208 4.5005
R54677 VINP.n241 VINP.n208 4.5005
R54678 VINP.n350 VINP.n208 4.5005
R54679 VINP.n240 VINP.n208 4.5005
R54680 VINP.n352 VINP.n208 4.5005
R54681 VINP.n239 VINP.n208 4.5005
R54682 VINP.n354 VINP.n208 4.5005
R54683 VINP.n238 VINP.n208 4.5005
R54684 VINP.n356 VINP.n208 4.5005
R54685 VINP.n237 VINP.n208 4.5005
R54686 VINP.n358 VINP.n208 4.5005
R54687 VINP.n236 VINP.n208 4.5005
R54688 VINP.n360 VINP.n208 4.5005
R54689 VINP.n235 VINP.n208 4.5005
R54690 VINP.n362 VINP.n208 4.5005
R54691 VINP.n234 VINP.n208 4.5005
R54692 VINP.n364 VINP.n208 4.5005
R54693 VINP.n233 VINP.n208 4.5005
R54694 VINP.n366 VINP.n208 4.5005
R54695 VINP.n232 VINP.n208 4.5005
R54696 VINP.n368 VINP.n208 4.5005
R54697 VINP.n231 VINP.n208 4.5005
R54698 VINP.n370 VINP.n208 4.5005
R54699 VINP.n230 VINP.n208 4.5005
R54700 VINP.n372 VINP.n208 4.5005
R54701 VINP.n229 VINP.n208 4.5005
R54702 VINP.n374 VINP.n208 4.5005
R54703 VINP.n228 VINP.n208 4.5005
R54704 VINP.n376 VINP.n208 4.5005
R54705 VINP.n227 VINP.n208 4.5005
R54706 VINP.n378 VINP.n208 4.5005
R54707 VINP.n226 VINP.n208 4.5005
R54708 VINP.n380 VINP.n208 4.5005
R54709 VINP.n225 VINP.n208 4.5005
R54710 VINP.n382 VINP.n208 4.5005
R54711 VINP.n224 VINP.n208 4.5005
R54712 VINP.n384 VINP.n208 4.5005
R54713 VINP.n223 VINP.n208 4.5005
R54714 VINP.n386 VINP.n208 4.5005
R54715 VINP.n222 VINP.n208 4.5005
R54716 VINP.n388 VINP.n208 4.5005
R54717 VINP.n221 VINP.n208 4.5005
R54718 VINP.n390 VINP.n208 4.5005
R54719 VINP.n220 VINP.n208 4.5005
R54720 VINP.n392 VINP.n208 4.5005
R54721 VINP.n219 VINP.n208 4.5005
R54722 VINP.n394 VINP.n208 4.5005
R54723 VINP.n218 VINP.n208 4.5005
R54724 VINP.n396 VINP.n208 4.5005
R54725 VINP.n217 VINP.n208 4.5005
R54726 VINP.n398 VINP.n208 4.5005
R54727 VINP.n216 VINP.n208 4.5005
R54728 VINP.n400 VINP.n208 4.5005
R54729 VINP.n215 VINP.n208 4.5005
R54730 VINP.n654 VINP.n208 4.5005
R54731 VINP.n656 VINP.n208 4.5005
R54732 VINP.n208 VINP.n0 4.5005
R54733 VINP.n278 VINP.n92 4.5005
R54734 VINP.n276 VINP.n92 4.5005
R54735 VINP.n280 VINP.n92 4.5005
R54736 VINP.n275 VINP.n92 4.5005
R54737 VINP.n282 VINP.n92 4.5005
R54738 VINP.n274 VINP.n92 4.5005
R54739 VINP.n284 VINP.n92 4.5005
R54740 VINP.n273 VINP.n92 4.5005
R54741 VINP.n286 VINP.n92 4.5005
R54742 VINP.n272 VINP.n92 4.5005
R54743 VINP.n288 VINP.n92 4.5005
R54744 VINP.n271 VINP.n92 4.5005
R54745 VINP.n290 VINP.n92 4.5005
R54746 VINP.n270 VINP.n92 4.5005
R54747 VINP.n292 VINP.n92 4.5005
R54748 VINP.n269 VINP.n92 4.5005
R54749 VINP.n294 VINP.n92 4.5005
R54750 VINP.n268 VINP.n92 4.5005
R54751 VINP.n296 VINP.n92 4.5005
R54752 VINP.n267 VINP.n92 4.5005
R54753 VINP.n298 VINP.n92 4.5005
R54754 VINP.n266 VINP.n92 4.5005
R54755 VINP.n300 VINP.n92 4.5005
R54756 VINP.n265 VINP.n92 4.5005
R54757 VINP.n302 VINP.n92 4.5005
R54758 VINP.n264 VINP.n92 4.5005
R54759 VINP.n304 VINP.n92 4.5005
R54760 VINP.n263 VINP.n92 4.5005
R54761 VINP.n306 VINP.n92 4.5005
R54762 VINP.n262 VINP.n92 4.5005
R54763 VINP.n308 VINP.n92 4.5005
R54764 VINP.n261 VINP.n92 4.5005
R54765 VINP.n310 VINP.n92 4.5005
R54766 VINP.n260 VINP.n92 4.5005
R54767 VINP.n312 VINP.n92 4.5005
R54768 VINP.n259 VINP.n92 4.5005
R54769 VINP.n314 VINP.n92 4.5005
R54770 VINP.n258 VINP.n92 4.5005
R54771 VINP.n316 VINP.n92 4.5005
R54772 VINP.n257 VINP.n92 4.5005
R54773 VINP.n318 VINP.n92 4.5005
R54774 VINP.n256 VINP.n92 4.5005
R54775 VINP.n320 VINP.n92 4.5005
R54776 VINP.n255 VINP.n92 4.5005
R54777 VINP.n322 VINP.n92 4.5005
R54778 VINP.n254 VINP.n92 4.5005
R54779 VINP.n324 VINP.n92 4.5005
R54780 VINP.n253 VINP.n92 4.5005
R54781 VINP.n326 VINP.n92 4.5005
R54782 VINP.n252 VINP.n92 4.5005
R54783 VINP.n328 VINP.n92 4.5005
R54784 VINP.n251 VINP.n92 4.5005
R54785 VINP.n330 VINP.n92 4.5005
R54786 VINP.n250 VINP.n92 4.5005
R54787 VINP.n332 VINP.n92 4.5005
R54788 VINP.n249 VINP.n92 4.5005
R54789 VINP.n334 VINP.n92 4.5005
R54790 VINP.n248 VINP.n92 4.5005
R54791 VINP.n336 VINP.n92 4.5005
R54792 VINP.n247 VINP.n92 4.5005
R54793 VINP.n338 VINP.n92 4.5005
R54794 VINP.n246 VINP.n92 4.5005
R54795 VINP.n340 VINP.n92 4.5005
R54796 VINP.n245 VINP.n92 4.5005
R54797 VINP.n342 VINP.n92 4.5005
R54798 VINP.n244 VINP.n92 4.5005
R54799 VINP.n344 VINP.n92 4.5005
R54800 VINP.n243 VINP.n92 4.5005
R54801 VINP.n346 VINP.n92 4.5005
R54802 VINP.n242 VINP.n92 4.5005
R54803 VINP.n348 VINP.n92 4.5005
R54804 VINP.n241 VINP.n92 4.5005
R54805 VINP.n350 VINP.n92 4.5005
R54806 VINP.n240 VINP.n92 4.5005
R54807 VINP.n352 VINP.n92 4.5005
R54808 VINP.n239 VINP.n92 4.5005
R54809 VINP.n354 VINP.n92 4.5005
R54810 VINP.n238 VINP.n92 4.5005
R54811 VINP.n356 VINP.n92 4.5005
R54812 VINP.n237 VINP.n92 4.5005
R54813 VINP.n358 VINP.n92 4.5005
R54814 VINP.n236 VINP.n92 4.5005
R54815 VINP.n360 VINP.n92 4.5005
R54816 VINP.n235 VINP.n92 4.5005
R54817 VINP.n362 VINP.n92 4.5005
R54818 VINP.n234 VINP.n92 4.5005
R54819 VINP.n364 VINP.n92 4.5005
R54820 VINP.n233 VINP.n92 4.5005
R54821 VINP.n366 VINP.n92 4.5005
R54822 VINP.n232 VINP.n92 4.5005
R54823 VINP.n368 VINP.n92 4.5005
R54824 VINP.n231 VINP.n92 4.5005
R54825 VINP.n370 VINP.n92 4.5005
R54826 VINP.n230 VINP.n92 4.5005
R54827 VINP.n372 VINP.n92 4.5005
R54828 VINP.n229 VINP.n92 4.5005
R54829 VINP.n374 VINP.n92 4.5005
R54830 VINP.n228 VINP.n92 4.5005
R54831 VINP.n376 VINP.n92 4.5005
R54832 VINP.n227 VINP.n92 4.5005
R54833 VINP.n378 VINP.n92 4.5005
R54834 VINP.n226 VINP.n92 4.5005
R54835 VINP.n380 VINP.n92 4.5005
R54836 VINP.n225 VINP.n92 4.5005
R54837 VINP.n382 VINP.n92 4.5005
R54838 VINP.n224 VINP.n92 4.5005
R54839 VINP.n384 VINP.n92 4.5005
R54840 VINP.n223 VINP.n92 4.5005
R54841 VINP.n386 VINP.n92 4.5005
R54842 VINP.n222 VINP.n92 4.5005
R54843 VINP.n388 VINP.n92 4.5005
R54844 VINP.n221 VINP.n92 4.5005
R54845 VINP.n390 VINP.n92 4.5005
R54846 VINP.n220 VINP.n92 4.5005
R54847 VINP.n392 VINP.n92 4.5005
R54848 VINP.n219 VINP.n92 4.5005
R54849 VINP.n394 VINP.n92 4.5005
R54850 VINP.n218 VINP.n92 4.5005
R54851 VINP.n396 VINP.n92 4.5005
R54852 VINP.n217 VINP.n92 4.5005
R54853 VINP.n398 VINP.n92 4.5005
R54854 VINP.n216 VINP.n92 4.5005
R54855 VINP.n400 VINP.n92 4.5005
R54856 VINP.n215 VINP.n92 4.5005
R54857 VINP.n654 VINP.n92 4.5005
R54858 VINP.n656 VINP.n92 4.5005
R54859 VINP.n92 VINP.n0 4.5005
R54860 VINP.n278 VINP.n209 4.5005
R54861 VINP.n276 VINP.n209 4.5005
R54862 VINP.n280 VINP.n209 4.5005
R54863 VINP.n275 VINP.n209 4.5005
R54864 VINP.n282 VINP.n209 4.5005
R54865 VINP.n274 VINP.n209 4.5005
R54866 VINP.n284 VINP.n209 4.5005
R54867 VINP.n273 VINP.n209 4.5005
R54868 VINP.n286 VINP.n209 4.5005
R54869 VINP.n272 VINP.n209 4.5005
R54870 VINP.n288 VINP.n209 4.5005
R54871 VINP.n271 VINP.n209 4.5005
R54872 VINP.n290 VINP.n209 4.5005
R54873 VINP.n270 VINP.n209 4.5005
R54874 VINP.n292 VINP.n209 4.5005
R54875 VINP.n269 VINP.n209 4.5005
R54876 VINP.n294 VINP.n209 4.5005
R54877 VINP.n268 VINP.n209 4.5005
R54878 VINP.n296 VINP.n209 4.5005
R54879 VINP.n267 VINP.n209 4.5005
R54880 VINP.n298 VINP.n209 4.5005
R54881 VINP.n266 VINP.n209 4.5005
R54882 VINP.n300 VINP.n209 4.5005
R54883 VINP.n265 VINP.n209 4.5005
R54884 VINP.n302 VINP.n209 4.5005
R54885 VINP.n264 VINP.n209 4.5005
R54886 VINP.n304 VINP.n209 4.5005
R54887 VINP.n263 VINP.n209 4.5005
R54888 VINP.n306 VINP.n209 4.5005
R54889 VINP.n262 VINP.n209 4.5005
R54890 VINP.n308 VINP.n209 4.5005
R54891 VINP.n261 VINP.n209 4.5005
R54892 VINP.n310 VINP.n209 4.5005
R54893 VINP.n260 VINP.n209 4.5005
R54894 VINP.n312 VINP.n209 4.5005
R54895 VINP.n259 VINP.n209 4.5005
R54896 VINP.n314 VINP.n209 4.5005
R54897 VINP.n258 VINP.n209 4.5005
R54898 VINP.n316 VINP.n209 4.5005
R54899 VINP.n257 VINP.n209 4.5005
R54900 VINP.n318 VINP.n209 4.5005
R54901 VINP.n256 VINP.n209 4.5005
R54902 VINP.n320 VINP.n209 4.5005
R54903 VINP.n255 VINP.n209 4.5005
R54904 VINP.n322 VINP.n209 4.5005
R54905 VINP.n254 VINP.n209 4.5005
R54906 VINP.n324 VINP.n209 4.5005
R54907 VINP.n253 VINP.n209 4.5005
R54908 VINP.n326 VINP.n209 4.5005
R54909 VINP.n252 VINP.n209 4.5005
R54910 VINP.n328 VINP.n209 4.5005
R54911 VINP.n251 VINP.n209 4.5005
R54912 VINP.n330 VINP.n209 4.5005
R54913 VINP.n250 VINP.n209 4.5005
R54914 VINP.n332 VINP.n209 4.5005
R54915 VINP.n249 VINP.n209 4.5005
R54916 VINP.n334 VINP.n209 4.5005
R54917 VINP.n248 VINP.n209 4.5005
R54918 VINP.n336 VINP.n209 4.5005
R54919 VINP.n247 VINP.n209 4.5005
R54920 VINP.n338 VINP.n209 4.5005
R54921 VINP.n246 VINP.n209 4.5005
R54922 VINP.n340 VINP.n209 4.5005
R54923 VINP.n245 VINP.n209 4.5005
R54924 VINP.n342 VINP.n209 4.5005
R54925 VINP.n244 VINP.n209 4.5005
R54926 VINP.n344 VINP.n209 4.5005
R54927 VINP.n243 VINP.n209 4.5005
R54928 VINP.n346 VINP.n209 4.5005
R54929 VINP.n242 VINP.n209 4.5005
R54930 VINP.n348 VINP.n209 4.5005
R54931 VINP.n241 VINP.n209 4.5005
R54932 VINP.n350 VINP.n209 4.5005
R54933 VINP.n240 VINP.n209 4.5005
R54934 VINP.n352 VINP.n209 4.5005
R54935 VINP.n239 VINP.n209 4.5005
R54936 VINP.n354 VINP.n209 4.5005
R54937 VINP.n238 VINP.n209 4.5005
R54938 VINP.n356 VINP.n209 4.5005
R54939 VINP.n237 VINP.n209 4.5005
R54940 VINP.n358 VINP.n209 4.5005
R54941 VINP.n236 VINP.n209 4.5005
R54942 VINP.n360 VINP.n209 4.5005
R54943 VINP.n235 VINP.n209 4.5005
R54944 VINP.n362 VINP.n209 4.5005
R54945 VINP.n234 VINP.n209 4.5005
R54946 VINP.n364 VINP.n209 4.5005
R54947 VINP.n233 VINP.n209 4.5005
R54948 VINP.n366 VINP.n209 4.5005
R54949 VINP.n232 VINP.n209 4.5005
R54950 VINP.n368 VINP.n209 4.5005
R54951 VINP.n231 VINP.n209 4.5005
R54952 VINP.n370 VINP.n209 4.5005
R54953 VINP.n230 VINP.n209 4.5005
R54954 VINP.n372 VINP.n209 4.5005
R54955 VINP.n229 VINP.n209 4.5005
R54956 VINP.n374 VINP.n209 4.5005
R54957 VINP.n228 VINP.n209 4.5005
R54958 VINP.n376 VINP.n209 4.5005
R54959 VINP.n227 VINP.n209 4.5005
R54960 VINP.n378 VINP.n209 4.5005
R54961 VINP.n226 VINP.n209 4.5005
R54962 VINP.n380 VINP.n209 4.5005
R54963 VINP.n225 VINP.n209 4.5005
R54964 VINP.n382 VINP.n209 4.5005
R54965 VINP.n224 VINP.n209 4.5005
R54966 VINP.n384 VINP.n209 4.5005
R54967 VINP.n223 VINP.n209 4.5005
R54968 VINP.n386 VINP.n209 4.5005
R54969 VINP.n222 VINP.n209 4.5005
R54970 VINP.n388 VINP.n209 4.5005
R54971 VINP.n221 VINP.n209 4.5005
R54972 VINP.n390 VINP.n209 4.5005
R54973 VINP.n220 VINP.n209 4.5005
R54974 VINP.n392 VINP.n209 4.5005
R54975 VINP.n219 VINP.n209 4.5005
R54976 VINP.n394 VINP.n209 4.5005
R54977 VINP.n218 VINP.n209 4.5005
R54978 VINP.n396 VINP.n209 4.5005
R54979 VINP.n217 VINP.n209 4.5005
R54980 VINP.n398 VINP.n209 4.5005
R54981 VINP.n216 VINP.n209 4.5005
R54982 VINP.n400 VINP.n209 4.5005
R54983 VINP.n215 VINP.n209 4.5005
R54984 VINP.n654 VINP.n209 4.5005
R54985 VINP.n656 VINP.n209 4.5005
R54986 VINP.n209 VINP.n0 4.5005
R54987 VINP.n278 VINP.n91 4.5005
R54988 VINP.n276 VINP.n91 4.5005
R54989 VINP.n280 VINP.n91 4.5005
R54990 VINP.n275 VINP.n91 4.5005
R54991 VINP.n282 VINP.n91 4.5005
R54992 VINP.n274 VINP.n91 4.5005
R54993 VINP.n284 VINP.n91 4.5005
R54994 VINP.n273 VINP.n91 4.5005
R54995 VINP.n286 VINP.n91 4.5005
R54996 VINP.n272 VINP.n91 4.5005
R54997 VINP.n288 VINP.n91 4.5005
R54998 VINP.n271 VINP.n91 4.5005
R54999 VINP.n290 VINP.n91 4.5005
R55000 VINP.n270 VINP.n91 4.5005
R55001 VINP.n292 VINP.n91 4.5005
R55002 VINP.n269 VINP.n91 4.5005
R55003 VINP.n294 VINP.n91 4.5005
R55004 VINP.n268 VINP.n91 4.5005
R55005 VINP.n296 VINP.n91 4.5005
R55006 VINP.n267 VINP.n91 4.5005
R55007 VINP.n298 VINP.n91 4.5005
R55008 VINP.n266 VINP.n91 4.5005
R55009 VINP.n300 VINP.n91 4.5005
R55010 VINP.n265 VINP.n91 4.5005
R55011 VINP.n302 VINP.n91 4.5005
R55012 VINP.n264 VINP.n91 4.5005
R55013 VINP.n304 VINP.n91 4.5005
R55014 VINP.n263 VINP.n91 4.5005
R55015 VINP.n306 VINP.n91 4.5005
R55016 VINP.n262 VINP.n91 4.5005
R55017 VINP.n308 VINP.n91 4.5005
R55018 VINP.n261 VINP.n91 4.5005
R55019 VINP.n310 VINP.n91 4.5005
R55020 VINP.n260 VINP.n91 4.5005
R55021 VINP.n312 VINP.n91 4.5005
R55022 VINP.n259 VINP.n91 4.5005
R55023 VINP.n314 VINP.n91 4.5005
R55024 VINP.n258 VINP.n91 4.5005
R55025 VINP.n316 VINP.n91 4.5005
R55026 VINP.n257 VINP.n91 4.5005
R55027 VINP.n318 VINP.n91 4.5005
R55028 VINP.n256 VINP.n91 4.5005
R55029 VINP.n320 VINP.n91 4.5005
R55030 VINP.n255 VINP.n91 4.5005
R55031 VINP.n322 VINP.n91 4.5005
R55032 VINP.n254 VINP.n91 4.5005
R55033 VINP.n324 VINP.n91 4.5005
R55034 VINP.n253 VINP.n91 4.5005
R55035 VINP.n326 VINP.n91 4.5005
R55036 VINP.n252 VINP.n91 4.5005
R55037 VINP.n328 VINP.n91 4.5005
R55038 VINP.n251 VINP.n91 4.5005
R55039 VINP.n330 VINP.n91 4.5005
R55040 VINP.n250 VINP.n91 4.5005
R55041 VINP.n332 VINP.n91 4.5005
R55042 VINP.n249 VINP.n91 4.5005
R55043 VINP.n334 VINP.n91 4.5005
R55044 VINP.n248 VINP.n91 4.5005
R55045 VINP.n336 VINP.n91 4.5005
R55046 VINP.n247 VINP.n91 4.5005
R55047 VINP.n338 VINP.n91 4.5005
R55048 VINP.n246 VINP.n91 4.5005
R55049 VINP.n340 VINP.n91 4.5005
R55050 VINP.n245 VINP.n91 4.5005
R55051 VINP.n342 VINP.n91 4.5005
R55052 VINP.n244 VINP.n91 4.5005
R55053 VINP.n344 VINP.n91 4.5005
R55054 VINP.n243 VINP.n91 4.5005
R55055 VINP.n346 VINP.n91 4.5005
R55056 VINP.n242 VINP.n91 4.5005
R55057 VINP.n348 VINP.n91 4.5005
R55058 VINP.n241 VINP.n91 4.5005
R55059 VINP.n350 VINP.n91 4.5005
R55060 VINP.n240 VINP.n91 4.5005
R55061 VINP.n352 VINP.n91 4.5005
R55062 VINP.n239 VINP.n91 4.5005
R55063 VINP.n354 VINP.n91 4.5005
R55064 VINP.n238 VINP.n91 4.5005
R55065 VINP.n356 VINP.n91 4.5005
R55066 VINP.n237 VINP.n91 4.5005
R55067 VINP.n358 VINP.n91 4.5005
R55068 VINP.n236 VINP.n91 4.5005
R55069 VINP.n360 VINP.n91 4.5005
R55070 VINP.n235 VINP.n91 4.5005
R55071 VINP.n362 VINP.n91 4.5005
R55072 VINP.n234 VINP.n91 4.5005
R55073 VINP.n364 VINP.n91 4.5005
R55074 VINP.n233 VINP.n91 4.5005
R55075 VINP.n366 VINP.n91 4.5005
R55076 VINP.n232 VINP.n91 4.5005
R55077 VINP.n368 VINP.n91 4.5005
R55078 VINP.n231 VINP.n91 4.5005
R55079 VINP.n370 VINP.n91 4.5005
R55080 VINP.n230 VINP.n91 4.5005
R55081 VINP.n372 VINP.n91 4.5005
R55082 VINP.n229 VINP.n91 4.5005
R55083 VINP.n374 VINP.n91 4.5005
R55084 VINP.n228 VINP.n91 4.5005
R55085 VINP.n376 VINP.n91 4.5005
R55086 VINP.n227 VINP.n91 4.5005
R55087 VINP.n378 VINP.n91 4.5005
R55088 VINP.n226 VINP.n91 4.5005
R55089 VINP.n380 VINP.n91 4.5005
R55090 VINP.n225 VINP.n91 4.5005
R55091 VINP.n382 VINP.n91 4.5005
R55092 VINP.n224 VINP.n91 4.5005
R55093 VINP.n384 VINP.n91 4.5005
R55094 VINP.n223 VINP.n91 4.5005
R55095 VINP.n386 VINP.n91 4.5005
R55096 VINP.n222 VINP.n91 4.5005
R55097 VINP.n388 VINP.n91 4.5005
R55098 VINP.n221 VINP.n91 4.5005
R55099 VINP.n390 VINP.n91 4.5005
R55100 VINP.n220 VINP.n91 4.5005
R55101 VINP.n392 VINP.n91 4.5005
R55102 VINP.n219 VINP.n91 4.5005
R55103 VINP.n394 VINP.n91 4.5005
R55104 VINP.n218 VINP.n91 4.5005
R55105 VINP.n396 VINP.n91 4.5005
R55106 VINP.n217 VINP.n91 4.5005
R55107 VINP.n398 VINP.n91 4.5005
R55108 VINP.n216 VINP.n91 4.5005
R55109 VINP.n400 VINP.n91 4.5005
R55110 VINP.n215 VINP.n91 4.5005
R55111 VINP.n654 VINP.n91 4.5005
R55112 VINP.n656 VINP.n91 4.5005
R55113 VINP.n91 VINP.n0 4.5005
R55114 VINP.n278 VINP.n210 4.5005
R55115 VINP.n276 VINP.n210 4.5005
R55116 VINP.n280 VINP.n210 4.5005
R55117 VINP.n275 VINP.n210 4.5005
R55118 VINP.n282 VINP.n210 4.5005
R55119 VINP.n274 VINP.n210 4.5005
R55120 VINP.n284 VINP.n210 4.5005
R55121 VINP.n273 VINP.n210 4.5005
R55122 VINP.n286 VINP.n210 4.5005
R55123 VINP.n272 VINP.n210 4.5005
R55124 VINP.n288 VINP.n210 4.5005
R55125 VINP.n271 VINP.n210 4.5005
R55126 VINP.n290 VINP.n210 4.5005
R55127 VINP.n270 VINP.n210 4.5005
R55128 VINP.n292 VINP.n210 4.5005
R55129 VINP.n269 VINP.n210 4.5005
R55130 VINP.n294 VINP.n210 4.5005
R55131 VINP.n268 VINP.n210 4.5005
R55132 VINP.n296 VINP.n210 4.5005
R55133 VINP.n267 VINP.n210 4.5005
R55134 VINP.n298 VINP.n210 4.5005
R55135 VINP.n266 VINP.n210 4.5005
R55136 VINP.n300 VINP.n210 4.5005
R55137 VINP.n265 VINP.n210 4.5005
R55138 VINP.n302 VINP.n210 4.5005
R55139 VINP.n264 VINP.n210 4.5005
R55140 VINP.n304 VINP.n210 4.5005
R55141 VINP.n263 VINP.n210 4.5005
R55142 VINP.n306 VINP.n210 4.5005
R55143 VINP.n262 VINP.n210 4.5005
R55144 VINP.n308 VINP.n210 4.5005
R55145 VINP.n261 VINP.n210 4.5005
R55146 VINP.n310 VINP.n210 4.5005
R55147 VINP.n260 VINP.n210 4.5005
R55148 VINP.n312 VINP.n210 4.5005
R55149 VINP.n259 VINP.n210 4.5005
R55150 VINP.n314 VINP.n210 4.5005
R55151 VINP.n258 VINP.n210 4.5005
R55152 VINP.n316 VINP.n210 4.5005
R55153 VINP.n257 VINP.n210 4.5005
R55154 VINP.n318 VINP.n210 4.5005
R55155 VINP.n256 VINP.n210 4.5005
R55156 VINP.n320 VINP.n210 4.5005
R55157 VINP.n255 VINP.n210 4.5005
R55158 VINP.n322 VINP.n210 4.5005
R55159 VINP.n254 VINP.n210 4.5005
R55160 VINP.n324 VINP.n210 4.5005
R55161 VINP.n253 VINP.n210 4.5005
R55162 VINP.n326 VINP.n210 4.5005
R55163 VINP.n252 VINP.n210 4.5005
R55164 VINP.n328 VINP.n210 4.5005
R55165 VINP.n251 VINP.n210 4.5005
R55166 VINP.n330 VINP.n210 4.5005
R55167 VINP.n250 VINP.n210 4.5005
R55168 VINP.n332 VINP.n210 4.5005
R55169 VINP.n249 VINP.n210 4.5005
R55170 VINP.n334 VINP.n210 4.5005
R55171 VINP.n248 VINP.n210 4.5005
R55172 VINP.n336 VINP.n210 4.5005
R55173 VINP.n247 VINP.n210 4.5005
R55174 VINP.n338 VINP.n210 4.5005
R55175 VINP.n246 VINP.n210 4.5005
R55176 VINP.n340 VINP.n210 4.5005
R55177 VINP.n245 VINP.n210 4.5005
R55178 VINP.n342 VINP.n210 4.5005
R55179 VINP.n244 VINP.n210 4.5005
R55180 VINP.n344 VINP.n210 4.5005
R55181 VINP.n243 VINP.n210 4.5005
R55182 VINP.n346 VINP.n210 4.5005
R55183 VINP.n242 VINP.n210 4.5005
R55184 VINP.n348 VINP.n210 4.5005
R55185 VINP.n241 VINP.n210 4.5005
R55186 VINP.n350 VINP.n210 4.5005
R55187 VINP.n240 VINP.n210 4.5005
R55188 VINP.n352 VINP.n210 4.5005
R55189 VINP.n239 VINP.n210 4.5005
R55190 VINP.n354 VINP.n210 4.5005
R55191 VINP.n238 VINP.n210 4.5005
R55192 VINP.n356 VINP.n210 4.5005
R55193 VINP.n237 VINP.n210 4.5005
R55194 VINP.n358 VINP.n210 4.5005
R55195 VINP.n236 VINP.n210 4.5005
R55196 VINP.n360 VINP.n210 4.5005
R55197 VINP.n235 VINP.n210 4.5005
R55198 VINP.n362 VINP.n210 4.5005
R55199 VINP.n234 VINP.n210 4.5005
R55200 VINP.n364 VINP.n210 4.5005
R55201 VINP.n233 VINP.n210 4.5005
R55202 VINP.n366 VINP.n210 4.5005
R55203 VINP.n232 VINP.n210 4.5005
R55204 VINP.n368 VINP.n210 4.5005
R55205 VINP.n231 VINP.n210 4.5005
R55206 VINP.n370 VINP.n210 4.5005
R55207 VINP.n230 VINP.n210 4.5005
R55208 VINP.n372 VINP.n210 4.5005
R55209 VINP.n229 VINP.n210 4.5005
R55210 VINP.n374 VINP.n210 4.5005
R55211 VINP.n228 VINP.n210 4.5005
R55212 VINP.n376 VINP.n210 4.5005
R55213 VINP.n227 VINP.n210 4.5005
R55214 VINP.n378 VINP.n210 4.5005
R55215 VINP.n226 VINP.n210 4.5005
R55216 VINP.n380 VINP.n210 4.5005
R55217 VINP.n225 VINP.n210 4.5005
R55218 VINP.n382 VINP.n210 4.5005
R55219 VINP.n224 VINP.n210 4.5005
R55220 VINP.n384 VINP.n210 4.5005
R55221 VINP.n223 VINP.n210 4.5005
R55222 VINP.n386 VINP.n210 4.5005
R55223 VINP.n222 VINP.n210 4.5005
R55224 VINP.n388 VINP.n210 4.5005
R55225 VINP.n221 VINP.n210 4.5005
R55226 VINP.n390 VINP.n210 4.5005
R55227 VINP.n220 VINP.n210 4.5005
R55228 VINP.n392 VINP.n210 4.5005
R55229 VINP.n219 VINP.n210 4.5005
R55230 VINP.n394 VINP.n210 4.5005
R55231 VINP.n218 VINP.n210 4.5005
R55232 VINP.n396 VINP.n210 4.5005
R55233 VINP.n217 VINP.n210 4.5005
R55234 VINP.n398 VINP.n210 4.5005
R55235 VINP.n216 VINP.n210 4.5005
R55236 VINP.n400 VINP.n210 4.5005
R55237 VINP.n215 VINP.n210 4.5005
R55238 VINP.n654 VINP.n210 4.5005
R55239 VINP.n656 VINP.n210 4.5005
R55240 VINP.n210 VINP.n0 4.5005
R55241 VINP.n278 VINP.n90 4.5005
R55242 VINP.n276 VINP.n90 4.5005
R55243 VINP.n280 VINP.n90 4.5005
R55244 VINP.n275 VINP.n90 4.5005
R55245 VINP.n282 VINP.n90 4.5005
R55246 VINP.n274 VINP.n90 4.5005
R55247 VINP.n284 VINP.n90 4.5005
R55248 VINP.n273 VINP.n90 4.5005
R55249 VINP.n286 VINP.n90 4.5005
R55250 VINP.n272 VINP.n90 4.5005
R55251 VINP.n288 VINP.n90 4.5005
R55252 VINP.n271 VINP.n90 4.5005
R55253 VINP.n290 VINP.n90 4.5005
R55254 VINP.n270 VINP.n90 4.5005
R55255 VINP.n292 VINP.n90 4.5005
R55256 VINP.n269 VINP.n90 4.5005
R55257 VINP.n294 VINP.n90 4.5005
R55258 VINP.n268 VINP.n90 4.5005
R55259 VINP.n296 VINP.n90 4.5005
R55260 VINP.n267 VINP.n90 4.5005
R55261 VINP.n298 VINP.n90 4.5005
R55262 VINP.n266 VINP.n90 4.5005
R55263 VINP.n300 VINP.n90 4.5005
R55264 VINP.n265 VINP.n90 4.5005
R55265 VINP.n302 VINP.n90 4.5005
R55266 VINP.n264 VINP.n90 4.5005
R55267 VINP.n304 VINP.n90 4.5005
R55268 VINP.n263 VINP.n90 4.5005
R55269 VINP.n306 VINP.n90 4.5005
R55270 VINP.n262 VINP.n90 4.5005
R55271 VINP.n308 VINP.n90 4.5005
R55272 VINP.n261 VINP.n90 4.5005
R55273 VINP.n310 VINP.n90 4.5005
R55274 VINP.n260 VINP.n90 4.5005
R55275 VINP.n312 VINP.n90 4.5005
R55276 VINP.n259 VINP.n90 4.5005
R55277 VINP.n314 VINP.n90 4.5005
R55278 VINP.n258 VINP.n90 4.5005
R55279 VINP.n316 VINP.n90 4.5005
R55280 VINP.n257 VINP.n90 4.5005
R55281 VINP.n318 VINP.n90 4.5005
R55282 VINP.n256 VINP.n90 4.5005
R55283 VINP.n320 VINP.n90 4.5005
R55284 VINP.n255 VINP.n90 4.5005
R55285 VINP.n322 VINP.n90 4.5005
R55286 VINP.n254 VINP.n90 4.5005
R55287 VINP.n324 VINP.n90 4.5005
R55288 VINP.n253 VINP.n90 4.5005
R55289 VINP.n326 VINP.n90 4.5005
R55290 VINP.n252 VINP.n90 4.5005
R55291 VINP.n328 VINP.n90 4.5005
R55292 VINP.n251 VINP.n90 4.5005
R55293 VINP.n330 VINP.n90 4.5005
R55294 VINP.n250 VINP.n90 4.5005
R55295 VINP.n332 VINP.n90 4.5005
R55296 VINP.n249 VINP.n90 4.5005
R55297 VINP.n334 VINP.n90 4.5005
R55298 VINP.n248 VINP.n90 4.5005
R55299 VINP.n336 VINP.n90 4.5005
R55300 VINP.n247 VINP.n90 4.5005
R55301 VINP.n338 VINP.n90 4.5005
R55302 VINP.n246 VINP.n90 4.5005
R55303 VINP.n340 VINP.n90 4.5005
R55304 VINP.n245 VINP.n90 4.5005
R55305 VINP.n342 VINP.n90 4.5005
R55306 VINP.n244 VINP.n90 4.5005
R55307 VINP.n344 VINP.n90 4.5005
R55308 VINP.n243 VINP.n90 4.5005
R55309 VINP.n346 VINP.n90 4.5005
R55310 VINP.n242 VINP.n90 4.5005
R55311 VINP.n348 VINP.n90 4.5005
R55312 VINP.n241 VINP.n90 4.5005
R55313 VINP.n350 VINP.n90 4.5005
R55314 VINP.n240 VINP.n90 4.5005
R55315 VINP.n352 VINP.n90 4.5005
R55316 VINP.n239 VINP.n90 4.5005
R55317 VINP.n354 VINP.n90 4.5005
R55318 VINP.n238 VINP.n90 4.5005
R55319 VINP.n356 VINP.n90 4.5005
R55320 VINP.n237 VINP.n90 4.5005
R55321 VINP.n358 VINP.n90 4.5005
R55322 VINP.n236 VINP.n90 4.5005
R55323 VINP.n360 VINP.n90 4.5005
R55324 VINP.n235 VINP.n90 4.5005
R55325 VINP.n362 VINP.n90 4.5005
R55326 VINP.n234 VINP.n90 4.5005
R55327 VINP.n364 VINP.n90 4.5005
R55328 VINP.n233 VINP.n90 4.5005
R55329 VINP.n366 VINP.n90 4.5005
R55330 VINP.n232 VINP.n90 4.5005
R55331 VINP.n368 VINP.n90 4.5005
R55332 VINP.n231 VINP.n90 4.5005
R55333 VINP.n370 VINP.n90 4.5005
R55334 VINP.n230 VINP.n90 4.5005
R55335 VINP.n372 VINP.n90 4.5005
R55336 VINP.n229 VINP.n90 4.5005
R55337 VINP.n374 VINP.n90 4.5005
R55338 VINP.n228 VINP.n90 4.5005
R55339 VINP.n376 VINP.n90 4.5005
R55340 VINP.n227 VINP.n90 4.5005
R55341 VINP.n378 VINP.n90 4.5005
R55342 VINP.n226 VINP.n90 4.5005
R55343 VINP.n380 VINP.n90 4.5005
R55344 VINP.n225 VINP.n90 4.5005
R55345 VINP.n382 VINP.n90 4.5005
R55346 VINP.n224 VINP.n90 4.5005
R55347 VINP.n384 VINP.n90 4.5005
R55348 VINP.n223 VINP.n90 4.5005
R55349 VINP.n386 VINP.n90 4.5005
R55350 VINP.n222 VINP.n90 4.5005
R55351 VINP.n388 VINP.n90 4.5005
R55352 VINP.n221 VINP.n90 4.5005
R55353 VINP.n390 VINP.n90 4.5005
R55354 VINP.n220 VINP.n90 4.5005
R55355 VINP.n392 VINP.n90 4.5005
R55356 VINP.n219 VINP.n90 4.5005
R55357 VINP.n394 VINP.n90 4.5005
R55358 VINP.n218 VINP.n90 4.5005
R55359 VINP.n396 VINP.n90 4.5005
R55360 VINP.n217 VINP.n90 4.5005
R55361 VINP.n398 VINP.n90 4.5005
R55362 VINP.n216 VINP.n90 4.5005
R55363 VINP.n400 VINP.n90 4.5005
R55364 VINP.n215 VINP.n90 4.5005
R55365 VINP.n654 VINP.n90 4.5005
R55366 VINP.n656 VINP.n90 4.5005
R55367 VINP.n90 VINP.n0 4.5005
R55368 VINP.n278 VINP.n211 4.5005
R55369 VINP.n276 VINP.n211 4.5005
R55370 VINP.n280 VINP.n211 4.5005
R55371 VINP.n275 VINP.n211 4.5005
R55372 VINP.n282 VINP.n211 4.5005
R55373 VINP.n274 VINP.n211 4.5005
R55374 VINP.n284 VINP.n211 4.5005
R55375 VINP.n273 VINP.n211 4.5005
R55376 VINP.n286 VINP.n211 4.5005
R55377 VINP.n272 VINP.n211 4.5005
R55378 VINP.n288 VINP.n211 4.5005
R55379 VINP.n271 VINP.n211 4.5005
R55380 VINP.n290 VINP.n211 4.5005
R55381 VINP.n270 VINP.n211 4.5005
R55382 VINP.n292 VINP.n211 4.5005
R55383 VINP.n269 VINP.n211 4.5005
R55384 VINP.n294 VINP.n211 4.5005
R55385 VINP.n268 VINP.n211 4.5005
R55386 VINP.n296 VINP.n211 4.5005
R55387 VINP.n267 VINP.n211 4.5005
R55388 VINP.n298 VINP.n211 4.5005
R55389 VINP.n266 VINP.n211 4.5005
R55390 VINP.n300 VINP.n211 4.5005
R55391 VINP.n265 VINP.n211 4.5005
R55392 VINP.n302 VINP.n211 4.5005
R55393 VINP.n264 VINP.n211 4.5005
R55394 VINP.n304 VINP.n211 4.5005
R55395 VINP.n263 VINP.n211 4.5005
R55396 VINP.n306 VINP.n211 4.5005
R55397 VINP.n262 VINP.n211 4.5005
R55398 VINP.n308 VINP.n211 4.5005
R55399 VINP.n261 VINP.n211 4.5005
R55400 VINP.n310 VINP.n211 4.5005
R55401 VINP.n260 VINP.n211 4.5005
R55402 VINP.n312 VINP.n211 4.5005
R55403 VINP.n259 VINP.n211 4.5005
R55404 VINP.n314 VINP.n211 4.5005
R55405 VINP.n258 VINP.n211 4.5005
R55406 VINP.n316 VINP.n211 4.5005
R55407 VINP.n257 VINP.n211 4.5005
R55408 VINP.n318 VINP.n211 4.5005
R55409 VINP.n256 VINP.n211 4.5005
R55410 VINP.n320 VINP.n211 4.5005
R55411 VINP.n255 VINP.n211 4.5005
R55412 VINP.n322 VINP.n211 4.5005
R55413 VINP.n254 VINP.n211 4.5005
R55414 VINP.n324 VINP.n211 4.5005
R55415 VINP.n253 VINP.n211 4.5005
R55416 VINP.n326 VINP.n211 4.5005
R55417 VINP.n252 VINP.n211 4.5005
R55418 VINP.n328 VINP.n211 4.5005
R55419 VINP.n251 VINP.n211 4.5005
R55420 VINP.n330 VINP.n211 4.5005
R55421 VINP.n250 VINP.n211 4.5005
R55422 VINP.n332 VINP.n211 4.5005
R55423 VINP.n249 VINP.n211 4.5005
R55424 VINP.n334 VINP.n211 4.5005
R55425 VINP.n248 VINP.n211 4.5005
R55426 VINP.n336 VINP.n211 4.5005
R55427 VINP.n247 VINP.n211 4.5005
R55428 VINP.n338 VINP.n211 4.5005
R55429 VINP.n246 VINP.n211 4.5005
R55430 VINP.n340 VINP.n211 4.5005
R55431 VINP.n245 VINP.n211 4.5005
R55432 VINP.n342 VINP.n211 4.5005
R55433 VINP.n244 VINP.n211 4.5005
R55434 VINP.n344 VINP.n211 4.5005
R55435 VINP.n243 VINP.n211 4.5005
R55436 VINP.n346 VINP.n211 4.5005
R55437 VINP.n242 VINP.n211 4.5005
R55438 VINP.n348 VINP.n211 4.5005
R55439 VINP.n241 VINP.n211 4.5005
R55440 VINP.n350 VINP.n211 4.5005
R55441 VINP.n240 VINP.n211 4.5005
R55442 VINP.n352 VINP.n211 4.5005
R55443 VINP.n239 VINP.n211 4.5005
R55444 VINP.n354 VINP.n211 4.5005
R55445 VINP.n238 VINP.n211 4.5005
R55446 VINP.n356 VINP.n211 4.5005
R55447 VINP.n237 VINP.n211 4.5005
R55448 VINP.n358 VINP.n211 4.5005
R55449 VINP.n236 VINP.n211 4.5005
R55450 VINP.n360 VINP.n211 4.5005
R55451 VINP.n235 VINP.n211 4.5005
R55452 VINP.n362 VINP.n211 4.5005
R55453 VINP.n234 VINP.n211 4.5005
R55454 VINP.n364 VINP.n211 4.5005
R55455 VINP.n233 VINP.n211 4.5005
R55456 VINP.n366 VINP.n211 4.5005
R55457 VINP.n232 VINP.n211 4.5005
R55458 VINP.n368 VINP.n211 4.5005
R55459 VINP.n231 VINP.n211 4.5005
R55460 VINP.n370 VINP.n211 4.5005
R55461 VINP.n230 VINP.n211 4.5005
R55462 VINP.n372 VINP.n211 4.5005
R55463 VINP.n229 VINP.n211 4.5005
R55464 VINP.n374 VINP.n211 4.5005
R55465 VINP.n228 VINP.n211 4.5005
R55466 VINP.n376 VINP.n211 4.5005
R55467 VINP.n227 VINP.n211 4.5005
R55468 VINP.n378 VINP.n211 4.5005
R55469 VINP.n226 VINP.n211 4.5005
R55470 VINP.n380 VINP.n211 4.5005
R55471 VINP.n225 VINP.n211 4.5005
R55472 VINP.n382 VINP.n211 4.5005
R55473 VINP.n224 VINP.n211 4.5005
R55474 VINP.n384 VINP.n211 4.5005
R55475 VINP.n223 VINP.n211 4.5005
R55476 VINP.n386 VINP.n211 4.5005
R55477 VINP.n222 VINP.n211 4.5005
R55478 VINP.n388 VINP.n211 4.5005
R55479 VINP.n221 VINP.n211 4.5005
R55480 VINP.n390 VINP.n211 4.5005
R55481 VINP.n220 VINP.n211 4.5005
R55482 VINP.n392 VINP.n211 4.5005
R55483 VINP.n219 VINP.n211 4.5005
R55484 VINP.n394 VINP.n211 4.5005
R55485 VINP.n218 VINP.n211 4.5005
R55486 VINP.n396 VINP.n211 4.5005
R55487 VINP.n217 VINP.n211 4.5005
R55488 VINP.n398 VINP.n211 4.5005
R55489 VINP.n216 VINP.n211 4.5005
R55490 VINP.n400 VINP.n211 4.5005
R55491 VINP.n215 VINP.n211 4.5005
R55492 VINP.n654 VINP.n211 4.5005
R55493 VINP.n656 VINP.n211 4.5005
R55494 VINP.n211 VINP.n0 4.5005
R55495 VINP.n278 VINP.n89 4.5005
R55496 VINP.n276 VINP.n89 4.5005
R55497 VINP.n280 VINP.n89 4.5005
R55498 VINP.n275 VINP.n89 4.5005
R55499 VINP.n282 VINP.n89 4.5005
R55500 VINP.n274 VINP.n89 4.5005
R55501 VINP.n284 VINP.n89 4.5005
R55502 VINP.n273 VINP.n89 4.5005
R55503 VINP.n286 VINP.n89 4.5005
R55504 VINP.n272 VINP.n89 4.5005
R55505 VINP.n288 VINP.n89 4.5005
R55506 VINP.n271 VINP.n89 4.5005
R55507 VINP.n290 VINP.n89 4.5005
R55508 VINP.n270 VINP.n89 4.5005
R55509 VINP.n292 VINP.n89 4.5005
R55510 VINP.n269 VINP.n89 4.5005
R55511 VINP.n294 VINP.n89 4.5005
R55512 VINP.n268 VINP.n89 4.5005
R55513 VINP.n296 VINP.n89 4.5005
R55514 VINP.n267 VINP.n89 4.5005
R55515 VINP.n298 VINP.n89 4.5005
R55516 VINP.n266 VINP.n89 4.5005
R55517 VINP.n300 VINP.n89 4.5005
R55518 VINP.n265 VINP.n89 4.5005
R55519 VINP.n302 VINP.n89 4.5005
R55520 VINP.n264 VINP.n89 4.5005
R55521 VINP.n304 VINP.n89 4.5005
R55522 VINP.n263 VINP.n89 4.5005
R55523 VINP.n306 VINP.n89 4.5005
R55524 VINP.n262 VINP.n89 4.5005
R55525 VINP.n308 VINP.n89 4.5005
R55526 VINP.n261 VINP.n89 4.5005
R55527 VINP.n310 VINP.n89 4.5005
R55528 VINP.n260 VINP.n89 4.5005
R55529 VINP.n312 VINP.n89 4.5005
R55530 VINP.n259 VINP.n89 4.5005
R55531 VINP.n314 VINP.n89 4.5005
R55532 VINP.n258 VINP.n89 4.5005
R55533 VINP.n316 VINP.n89 4.5005
R55534 VINP.n257 VINP.n89 4.5005
R55535 VINP.n318 VINP.n89 4.5005
R55536 VINP.n256 VINP.n89 4.5005
R55537 VINP.n320 VINP.n89 4.5005
R55538 VINP.n255 VINP.n89 4.5005
R55539 VINP.n322 VINP.n89 4.5005
R55540 VINP.n254 VINP.n89 4.5005
R55541 VINP.n324 VINP.n89 4.5005
R55542 VINP.n253 VINP.n89 4.5005
R55543 VINP.n326 VINP.n89 4.5005
R55544 VINP.n252 VINP.n89 4.5005
R55545 VINP.n328 VINP.n89 4.5005
R55546 VINP.n251 VINP.n89 4.5005
R55547 VINP.n330 VINP.n89 4.5005
R55548 VINP.n250 VINP.n89 4.5005
R55549 VINP.n332 VINP.n89 4.5005
R55550 VINP.n249 VINP.n89 4.5005
R55551 VINP.n334 VINP.n89 4.5005
R55552 VINP.n248 VINP.n89 4.5005
R55553 VINP.n336 VINP.n89 4.5005
R55554 VINP.n247 VINP.n89 4.5005
R55555 VINP.n338 VINP.n89 4.5005
R55556 VINP.n246 VINP.n89 4.5005
R55557 VINP.n340 VINP.n89 4.5005
R55558 VINP.n245 VINP.n89 4.5005
R55559 VINP.n342 VINP.n89 4.5005
R55560 VINP.n244 VINP.n89 4.5005
R55561 VINP.n344 VINP.n89 4.5005
R55562 VINP.n243 VINP.n89 4.5005
R55563 VINP.n346 VINP.n89 4.5005
R55564 VINP.n242 VINP.n89 4.5005
R55565 VINP.n348 VINP.n89 4.5005
R55566 VINP.n241 VINP.n89 4.5005
R55567 VINP.n350 VINP.n89 4.5005
R55568 VINP.n240 VINP.n89 4.5005
R55569 VINP.n352 VINP.n89 4.5005
R55570 VINP.n239 VINP.n89 4.5005
R55571 VINP.n354 VINP.n89 4.5005
R55572 VINP.n238 VINP.n89 4.5005
R55573 VINP.n356 VINP.n89 4.5005
R55574 VINP.n237 VINP.n89 4.5005
R55575 VINP.n358 VINP.n89 4.5005
R55576 VINP.n236 VINP.n89 4.5005
R55577 VINP.n360 VINP.n89 4.5005
R55578 VINP.n235 VINP.n89 4.5005
R55579 VINP.n362 VINP.n89 4.5005
R55580 VINP.n234 VINP.n89 4.5005
R55581 VINP.n364 VINP.n89 4.5005
R55582 VINP.n233 VINP.n89 4.5005
R55583 VINP.n366 VINP.n89 4.5005
R55584 VINP.n232 VINP.n89 4.5005
R55585 VINP.n368 VINP.n89 4.5005
R55586 VINP.n231 VINP.n89 4.5005
R55587 VINP.n370 VINP.n89 4.5005
R55588 VINP.n230 VINP.n89 4.5005
R55589 VINP.n372 VINP.n89 4.5005
R55590 VINP.n229 VINP.n89 4.5005
R55591 VINP.n374 VINP.n89 4.5005
R55592 VINP.n228 VINP.n89 4.5005
R55593 VINP.n376 VINP.n89 4.5005
R55594 VINP.n227 VINP.n89 4.5005
R55595 VINP.n378 VINP.n89 4.5005
R55596 VINP.n226 VINP.n89 4.5005
R55597 VINP.n380 VINP.n89 4.5005
R55598 VINP.n225 VINP.n89 4.5005
R55599 VINP.n382 VINP.n89 4.5005
R55600 VINP.n224 VINP.n89 4.5005
R55601 VINP.n384 VINP.n89 4.5005
R55602 VINP.n223 VINP.n89 4.5005
R55603 VINP.n386 VINP.n89 4.5005
R55604 VINP.n222 VINP.n89 4.5005
R55605 VINP.n388 VINP.n89 4.5005
R55606 VINP.n221 VINP.n89 4.5005
R55607 VINP.n390 VINP.n89 4.5005
R55608 VINP.n220 VINP.n89 4.5005
R55609 VINP.n392 VINP.n89 4.5005
R55610 VINP.n219 VINP.n89 4.5005
R55611 VINP.n394 VINP.n89 4.5005
R55612 VINP.n218 VINP.n89 4.5005
R55613 VINP.n396 VINP.n89 4.5005
R55614 VINP.n217 VINP.n89 4.5005
R55615 VINP.n398 VINP.n89 4.5005
R55616 VINP.n216 VINP.n89 4.5005
R55617 VINP.n400 VINP.n89 4.5005
R55618 VINP.n215 VINP.n89 4.5005
R55619 VINP.n654 VINP.n89 4.5005
R55620 VINP.n656 VINP.n89 4.5005
R55621 VINP.n89 VINP.n0 4.5005
R55622 VINP.n278 VINP.n212 4.5005
R55623 VINP.n276 VINP.n212 4.5005
R55624 VINP.n280 VINP.n212 4.5005
R55625 VINP.n275 VINP.n212 4.5005
R55626 VINP.n282 VINP.n212 4.5005
R55627 VINP.n274 VINP.n212 4.5005
R55628 VINP.n284 VINP.n212 4.5005
R55629 VINP.n273 VINP.n212 4.5005
R55630 VINP.n286 VINP.n212 4.5005
R55631 VINP.n272 VINP.n212 4.5005
R55632 VINP.n288 VINP.n212 4.5005
R55633 VINP.n271 VINP.n212 4.5005
R55634 VINP.n290 VINP.n212 4.5005
R55635 VINP.n270 VINP.n212 4.5005
R55636 VINP.n292 VINP.n212 4.5005
R55637 VINP.n269 VINP.n212 4.5005
R55638 VINP.n294 VINP.n212 4.5005
R55639 VINP.n268 VINP.n212 4.5005
R55640 VINP.n296 VINP.n212 4.5005
R55641 VINP.n267 VINP.n212 4.5005
R55642 VINP.n298 VINP.n212 4.5005
R55643 VINP.n266 VINP.n212 4.5005
R55644 VINP.n300 VINP.n212 4.5005
R55645 VINP.n265 VINP.n212 4.5005
R55646 VINP.n302 VINP.n212 4.5005
R55647 VINP.n264 VINP.n212 4.5005
R55648 VINP.n304 VINP.n212 4.5005
R55649 VINP.n263 VINP.n212 4.5005
R55650 VINP.n306 VINP.n212 4.5005
R55651 VINP.n262 VINP.n212 4.5005
R55652 VINP.n308 VINP.n212 4.5005
R55653 VINP.n261 VINP.n212 4.5005
R55654 VINP.n310 VINP.n212 4.5005
R55655 VINP.n260 VINP.n212 4.5005
R55656 VINP.n312 VINP.n212 4.5005
R55657 VINP.n259 VINP.n212 4.5005
R55658 VINP.n314 VINP.n212 4.5005
R55659 VINP.n258 VINP.n212 4.5005
R55660 VINP.n316 VINP.n212 4.5005
R55661 VINP.n257 VINP.n212 4.5005
R55662 VINP.n318 VINP.n212 4.5005
R55663 VINP.n256 VINP.n212 4.5005
R55664 VINP.n320 VINP.n212 4.5005
R55665 VINP.n255 VINP.n212 4.5005
R55666 VINP.n322 VINP.n212 4.5005
R55667 VINP.n254 VINP.n212 4.5005
R55668 VINP.n324 VINP.n212 4.5005
R55669 VINP.n253 VINP.n212 4.5005
R55670 VINP.n326 VINP.n212 4.5005
R55671 VINP.n252 VINP.n212 4.5005
R55672 VINP.n328 VINP.n212 4.5005
R55673 VINP.n251 VINP.n212 4.5005
R55674 VINP.n330 VINP.n212 4.5005
R55675 VINP.n250 VINP.n212 4.5005
R55676 VINP.n332 VINP.n212 4.5005
R55677 VINP.n249 VINP.n212 4.5005
R55678 VINP.n334 VINP.n212 4.5005
R55679 VINP.n248 VINP.n212 4.5005
R55680 VINP.n336 VINP.n212 4.5005
R55681 VINP.n247 VINP.n212 4.5005
R55682 VINP.n338 VINP.n212 4.5005
R55683 VINP.n246 VINP.n212 4.5005
R55684 VINP.n340 VINP.n212 4.5005
R55685 VINP.n245 VINP.n212 4.5005
R55686 VINP.n342 VINP.n212 4.5005
R55687 VINP.n244 VINP.n212 4.5005
R55688 VINP.n344 VINP.n212 4.5005
R55689 VINP.n243 VINP.n212 4.5005
R55690 VINP.n346 VINP.n212 4.5005
R55691 VINP.n242 VINP.n212 4.5005
R55692 VINP.n348 VINP.n212 4.5005
R55693 VINP.n241 VINP.n212 4.5005
R55694 VINP.n350 VINP.n212 4.5005
R55695 VINP.n240 VINP.n212 4.5005
R55696 VINP.n352 VINP.n212 4.5005
R55697 VINP.n239 VINP.n212 4.5005
R55698 VINP.n354 VINP.n212 4.5005
R55699 VINP.n238 VINP.n212 4.5005
R55700 VINP.n356 VINP.n212 4.5005
R55701 VINP.n237 VINP.n212 4.5005
R55702 VINP.n358 VINP.n212 4.5005
R55703 VINP.n236 VINP.n212 4.5005
R55704 VINP.n360 VINP.n212 4.5005
R55705 VINP.n235 VINP.n212 4.5005
R55706 VINP.n362 VINP.n212 4.5005
R55707 VINP.n234 VINP.n212 4.5005
R55708 VINP.n364 VINP.n212 4.5005
R55709 VINP.n233 VINP.n212 4.5005
R55710 VINP.n366 VINP.n212 4.5005
R55711 VINP.n232 VINP.n212 4.5005
R55712 VINP.n368 VINP.n212 4.5005
R55713 VINP.n231 VINP.n212 4.5005
R55714 VINP.n370 VINP.n212 4.5005
R55715 VINP.n230 VINP.n212 4.5005
R55716 VINP.n372 VINP.n212 4.5005
R55717 VINP.n229 VINP.n212 4.5005
R55718 VINP.n374 VINP.n212 4.5005
R55719 VINP.n228 VINP.n212 4.5005
R55720 VINP.n376 VINP.n212 4.5005
R55721 VINP.n227 VINP.n212 4.5005
R55722 VINP.n378 VINP.n212 4.5005
R55723 VINP.n226 VINP.n212 4.5005
R55724 VINP.n380 VINP.n212 4.5005
R55725 VINP.n225 VINP.n212 4.5005
R55726 VINP.n382 VINP.n212 4.5005
R55727 VINP.n224 VINP.n212 4.5005
R55728 VINP.n384 VINP.n212 4.5005
R55729 VINP.n223 VINP.n212 4.5005
R55730 VINP.n386 VINP.n212 4.5005
R55731 VINP.n222 VINP.n212 4.5005
R55732 VINP.n388 VINP.n212 4.5005
R55733 VINP.n221 VINP.n212 4.5005
R55734 VINP.n390 VINP.n212 4.5005
R55735 VINP.n220 VINP.n212 4.5005
R55736 VINP.n392 VINP.n212 4.5005
R55737 VINP.n219 VINP.n212 4.5005
R55738 VINP.n394 VINP.n212 4.5005
R55739 VINP.n218 VINP.n212 4.5005
R55740 VINP.n396 VINP.n212 4.5005
R55741 VINP.n217 VINP.n212 4.5005
R55742 VINP.n398 VINP.n212 4.5005
R55743 VINP.n216 VINP.n212 4.5005
R55744 VINP.n400 VINP.n212 4.5005
R55745 VINP.n215 VINP.n212 4.5005
R55746 VINP.n654 VINP.n212 4.5005
R55747 VINP.n656 VINP.n212 4.5005
R55748 VINP.n212 VINP.n0 4.5005
R55749 VINP.n278 VINP.n88 4.5005
R55750 VINP.n276 VINP.n88 4.5005
R55751 VINP.n280 VINP.n88 4.5005
R55752 VINP.n275 VINP.n88 4.5005
R55753 VINP.n282 VINP.n88 4.5005
R55754 VINP.n274 VINP.n88 4.5005
R55755 VINP.n284 VINP.n88 4.5005
R55756 VINP.n273 VINP.n88 4.5005
R55757 VINP.n286 VINP.n88 4.5005
R55758 VINP.n272 VINP.n88 4.5005
R55759 VINP.n288 VINP.n88 4.5005
R55760 VINP.n271 VINP.n88 4.5005
R55761 VINP.n290 VINP.n88 4.5005
R55762 VINP.n270 VINP.n88 4.5005
R55763 VINP.n292 VINP.n88 4.5005
R55764 VINP.n269 VINP.n88 4.5005
R55765 VINP.n294 VINP.n88 4.5005
R55766 VINP.n268 VINP.n88 4.5005
R55767 VINP.n296 VINP.n88 4.5005
R55768 VINP.n267 VINP.n88 4.5005
R55769 VINP.n298 VINP.n88 4.5005
R55770 VINP.n266 VINP.n88 4.5005
R55771 VINP.n300 VINP.n88 4.5005
R55772 VINP.n265 VINP.n88 4.5005
R55773 VINP.n302 VINP.n88 4.5005
R55774 VINP.n264 VINP.n88 4.5005
R55775 VINP.n304 VINP.n88 4.5005
R55776 VINP.n263 VINP.n88 4.5005
R55777 VINP.n306 VINP.n88 4.5005
R55778 VINP.n262 VINP.n88 4.5005
R55779 VINP.n308 VINP.n88 4.5005
R55780 VINP.n261 VINP.n88 4.5005
R55781 VINP.n310 VINP.n88 4.5005
R55782 VINP.n260 VINP.n88 4.5005
R55783 VINP.n312 VINP.n88 4.5005
R55784 VINP.n259 VINP.n88 4.5005
R55785 VINP.n314 VINP.n88 4.5005
R55786 VINP.n258 VINP.n88 4.5005
R55787 VINP.n316 VINP.n88 4.5005
R55788 VINP.n257 VINP.n88 4.5005
R55789 VINP.n318 VINP.n88 4.5005
R55790 VINP.n256 VINP.n88 4.5005
R55791 VINP.n320 VINP.n88 4.5005
R55792 VINP.n255 VINP.n88 4.5005
R55793 VINP.n322 VINP.n88 4.5005
R55794 VINP.n254 VINP.n88 4.5005
R55795 VINP.n324 VINP.n88 4.5005
R55796 VINP.n253 VINP.n88 4.5005
R55797 VINP.n326 VINP.n88 4.5005
R55798 VINP.n252 VINP.n88 4.5005
R55799 VINP.n328 VINP.n88 4.5005
R55800 VINP.n251 VINP.n88 4.5005
R55801 VINP.n330 VINP.n88 4.5005
R55802 VINP.n250 VINP.n88 4.5005
R55803 VINP.n332 VINP.n88 4.5005
R55804 VINP.n249 VINP.n88 4.5005
R55805 VINP.n334 VINP.n88 4.5005
R55806 VINP.n248 VINP.n88 4.5005
R55807 VINP.n336 VINP.n88 4.5005
R55808 VINP.n247 VINP.n88 4.5005
R55809 VINP.n338 VINP.n88 4.5005
R55810 VINP.n246 VINP.n88 4.5005
R55811 VINP.n340 VINP.n88 4.5005
R55812 VINP.n245 VINP.n88 4.5005
R55813 VINP.n342 VINP.n88 4.5005
R55814 VINP.n244 VINP.n88 4.5005
R55815 VINP.n344 VINP.n88 4.5005
R55816 VINP.n243 VINP.n88 4.5005
R55817 VINP.n346 VINP.n88 4.5005
R55818 VINP.n242 VINP.n88 4.5005
R55819 VINP.n348 VINP.n88 4.5005
R55820 VINP.n241 VINP.n88 4.5005
R55821 VINP.n350 VINP.n88 4.5005
R55822 VINP.n240 VINP.n88 4.5005
R55823 VINP.n352 VINP.n88 4.5005
R55824 VINP.n239 VINP.n88 4.5005
R55825 VINP.n354 VINP.n88 4.5005
R55826 VINP.n238 VINP.n88 4.5005
R55827 VINP.n356 VINP.n88 4.5005
R55828 VINP.n237 VINP.n88 4.5005
R55829 VINP.n358 VINP.n88 4.5005
R55830 VINP.n236 VINP.n88 4.5005
R55831 VINP.n360 VINP.n88 4.5005
R55832 VINP.n235 VINP.n88 4.5005
R55833 VINP.n362 VINP.n88 4.5005
R55834 VINP.n234 VINP.n88 4.5005
R55835 VINP.n364 VINP.n88 4.5005
R55836 VINP.n233 VINP.n88 4.5005
R55837 VINP.n366 VINP.n88 4.5005
R55838 VINP.n232 VINP.n88 4.5005
R55839 VINP.n368 VINP.n88 4.5005
R55840 VINP.n231 VINP.n88 4.5005
R55841 VINP.n370 VINP.n88 4.5005
R55842 VINP.n230 VINP.n88 4.5005
R55843 VINP.n372 VINP.n88 4.5005
R55844 VINP.n229 VINP.n88 4.5005
R55845 VINP.n374 VINP.n88 4.5005
R55846 VINP.n228 VINP.n88 4.5005
R55847 VINP.n376 VINP.n88 4.5005
R55848 VINP.n227 VINP.n88 4.5005
R55849 VINP.n378 VINP.n88 4.5005
R55850 VINP.n226 VINP.n88 4.5005
R55851 VINP.n380 VINP.n88 4.5005
R55852 VINP.n225 VINP.n88 4.5005
R55853 VINP.n382 VINP.n88 4.5005
R55854 VINP.n224 VINP.n88 4.5005
R55855 VINP.n384 VINP.n88 4.5005
R55856 VINP.n223 VINP.n88 4.5005
R55857 VINP.n386 VINP.n88 4.5005
R55858 VINP.n222 VINP.n88 4.5005
R55859 VINP.n388 VINP.n88 4.5005
R55860 VINP.n221 VINP.n88 4.5005
R55861 VINP.n390 VINP.n88 4.5005
R55862 VINP.n220 VINP.n88 4.5005
R55863 VINP.n392 VINP.n88 4.5005
R55864 VINP.n219 VINP.n88 4.5005
R55865 VINP.n394 VINP.n88 4.5005
R55866 VINP.n218 VINP.n88 4.5005
R55867 VINP.n396 VINP.n88 4.5005
R55868 VINP.n217 VINP.n88 4.5005
R55869 VINP.n398 VINP.n88 4.5005
R55870 VINP.n216 VINP.n88 4.5005
R55871 VINP.n400 VINP.n88 4.5005
R55872 VINP.n215 VINP.n88 4.5005
R55873 VINP.n654 VINP.n88 4.5005
R55874 VINP.n656 VINP.n88 4.5005
R55875 VINP.n88 VINP.n0 4.5005
R55876 VINP.n278 VINP.n213 4.5005
R55877 VINP.n276 VINP.n213 4.5005
R55878 VINP.n280 VINP.n213 4.5005
R55879 VINP.n275 VINP.n213 4.5005
R55880 VINP.n282 VINP.n213 4.5005
R55881 VINP.n274 VINP.n213 4.5005
R55882 VINP.n284 VINP.n213 4.5005
R55883 VINP.n273 VINP.n213 4.5005
R55884 VINP.n286 VINP.n213 4.5005
R55885 VINP.n272 VINP.n213 4.5005
R55886 VINP.n288 VINP.n213 4.5005
R55887 VINP.n271 VINP.n213 4.5005
R55888 VINP.n290 VINP.n213 4.5005
R55889 VINP.n270 VINP.n213 4.5005
R55890 VINP.n292 VINP.n213 4.5005
R55891 VINP.n269 VINP.n213 4.5005
R55892 VINP.n294 VINP.n213 4.5005
R55893 VINP.n268 VINP.n213 4.5005
R55894 VINP.n296 VINP.n213 4.5005
R55895 VINP.n267 VINP.n213 4.5005
R55896 VINP.n298 VINP.n213 4.5005
R55897 VINP.n266 VINP.n213 4.5005
R55898 VINP.n300 VINP.n213 4.5005
R55899 VINP.n265 VINP.n213 4.5005
R55900 VINP.n302 VINP.n213 4.5005
R55901 VINP.n264 VINP.n213 4.5005
R55902 VINP.n304 VINP.n213 4.5005
R55903 VINP.n263 VINP.n213 4.5005
R55904 VINP.n306 VINP.n213 4.5005
R55905 VINP.n262 VINP.n213 4.5005
R55906 VINP.n308 VINP.n213 4.5005
R55907 VINP.n261 VINP.n213 4.5005
R55908 VINP.n310 VINP.n213 4.5005
R55909 VINP.n260 VINP.n213 4.5005
R55910 VINP.n312 VINP.n213 4.5005
R55911 VINP.n259 VINP.n213 4.5005
R55912 VINP.n314 VINP.n213 4.5005
R55913 VINP.n258 VINP.n213 4.5005
R55914 VINP.n316 VINP.n213 4.5005
R55915 VINP.n257 VINP.n213 4.5005
R55916 VINP.n318 VINP.n213 4.5005
R55917 VINP.n256 VINP.n213 4.5005
R55918 VINP.n320 VINP.n213 4.5005
R55919 VINP.n255 VINP.n213 4.5005
R55920 VINP.n322 VINP.n213 4.5005
R55921 VINP.n254 VINP.n213 4.5005
R55922 VINP.n324 VINP.n213 4.5005
R55923 VINP.n253 VINP.n213 4.5005
R55924 VINP.n326 VINP.n213 4.5005
R55925 VINP.n252 VINP.n213 4.5005
R55926 VINP.n328 VINP.n213 4.5005
R55927 VINP.n251 VINP.n213 4.5005
R55928 VINP.n330 VINP.n213 4.5005
R55929 VINP.n250 VINP.n213 4.5005
R55930 VINP.n332 VINP.n213 4.5005
R55931 VINP.n249 VINP.n213 4.5005
R55932 VINP.n334 VINP.n213 4.5005
R55933 VINP.n248 VINP.n213 4.5005
R55934 VINP.n336 VINP.n213 4.5005
R55935 VINP.n247 VINP.n213 4.5005
R55936 VINP.n338 VINP.n213 4.5005
R55937 VINP.n246 VINP.n213 4.5005
R55938 VINP.n340 VINP.n213 4.5005
R55939 VINP.n245 VINP.n213 4.5005
R55940 VINP.n342 VINP.n213 4.5005
R55941 VINP.n244 VINP.n213 4.5005
R55942 VINP.n344 VINP.n213 4.5005
R55943 VINP.n243 VINP.n213 4.5005
R55944 VINP.n346 VINP.n213 4.5005
R55945 VINP.n242 VINP.n213 4.5005
R55946 VINP.n348 VINP.n213 4.5005
R55947 VINP.n241 VINP.n213 4.5005
R55948 VINP.n350 VINP.n213 4.5005
R55949 VINP.n240 VINP.n213 4.5005
R55950 VINP.n352 VINP.n213 4.5005
R55951 VINP.n239 VINP.n213 4.5005
R55952 VINP.n354 VINP.n213 4.5005
R55953 VINP.n238 VINP.n213 4.5005
R55954 VINP.n356 VINP.n213 4.5005
R55955 VINP.n237 VINP.n213 4.5005
R55956 VINP.n358 VINP.n213 4.5005
R55957 VINP.n236 VINP.n213 4.5005
R55958 VINP.n360 VINP.n213 4.5005
R55959 VINP.n235 VINP.n213 4.5005
R55960 VINP.n362 VINP.n213 4.5005
R55961 VINP.n234 VINP.n213 4.5005
R55962 VINP.n364 VINP.n213 4.5005
R55963 VINP.n233 VINP.n213 4.5005
R55964 VINP.n366 VINP.n213 4.5005
R55965 VINP.n232 VINP.n213 4.5005
R55966 VINP.n368 VINP.n213 4.5005
R55967 VINP.n231 VINP.n213 4.5005
R55968 VINP.n370 VINP.n213 4.5005
R55969 VINP.n230 VINP.n213 4.5005
R55970 VINP.n372 VINP.n213 4.5005
R55971 VINP.n229 VINP.n213 4.5005
R55972 VINP.n374 VINP.n213 4.5005
R55973 VINP.n228 VINP.n213 4.5005
R55974 VINP.n376 VINP.n213 4.5005
R55975 VINP.n227 VINP.n213 4.5005
R55976 VINP.n378 VINP.n213 4.5005
R55977 VINP.n226 VINP.n213 4.5005
R55978 VINP.n380 VINP.n213 4.5005
R55979 VINP.n225 VINP.n213 4.5005
R55980 VINP.n382 VINP.n213 4.5005
R55981 VINP.n224 VINP.n213 4.5005
R55982 VINP.n384 VINP.n213 4.5005
R55983 VINP.n223 VINP.n213 4.5005
R55984 VINP.n386 VINP.n213 4.5005
R55985 VINP.n222 VINP.n213 4.5005
R55986 VINP.n388 VINP.n213 4.5005
R55987 VINP.n221 VINP.n213 4.5005
R55988 VINP.n390 VINP.n213 4.5005
R55989 VINP.n220 VINP.n213 4.5005
R55990 VINP.n392 VINP.n213 4.5005
R55991 VINP.n219 VINP.n213 4.5005
R55992 VINP.n394 VINP.n213 4.5005
R55993 VINP.n218 VINP.n213 4.5005
R55994 VINP.n396 VINP.n213 4.5005
R55995 VINP.n217 VINP.n213 4.5005
R55996 VINP.n398 VINP.n213 4.5005
R55997 VINP.n216 VINP.n213 4.5005
R55998 VINP.n400 VINP.n213 4.5005
R55999 VINP.n215 VINP.n213 4.5005
R56000 VINP.n654 VINP.n213 4.5005
R56001 VINP.n656 VINP.n213 4.5005
R56002 VINP.n213 VINP.n0 4.5005
R56003 VINP.n278 VINP.n87 4.5005
R56004 VINP.n276 VINP.n87 4.5005
R56005 VINP.n280 VINP.n87 4.5005
R56006 VINP.n275 VINP.n87 4.5005
R56007 VINP.n282 VINP.n87 4.5005
R56008 VINP.n274 VINP.n87 4.5005
R56009 VINP.n284 VINP.n87 4.5005
R56010 VINP.n273 VINP.n87 4.5005
R56011 VINP.n286 VINP.n87 4.5005
R56012 VINP.n272 VINP.n87 4.5005
R56013 VINP.n288 VINP.n87 4.5005
R56014 VINP.n271 VINP.n87 4.5005
R56015 VINP.n290 VINP.n87 4.5005
R56016 VINP.n270 VINP.n87 4.5005
R56017 VINP.n292 VINP.n87 4.5005
R56018 VINP.n269 VINP.n87 4.5005
R56019 VINP.n294 VINP.n87 4.5005
R56020 VINP.n268 VINP.n87 4.5005
R56021 VINP.n296 VINP.n87 4.5005
R56022 VINP.n267 VINP.n87 4.5005
R56023 VINP.n298 VINP.n87 4.5005
R56024 VINP.n266 VINP.n87 4.5005
R56025 VINP.n300 VINP.n87 4.5005
R56026 VINP.n265 VINP.n87 4.5005
R56027 VINP.n302 VINP.n87 4.5005
R56028 VINP.n264 VINP.n87 4.5005
R56029 VINP.n304 VINP.n87 4.5005
R56030 VINP.n263 VINP.n87 4.5005
R56031 VINP.n306 VINP.n87 4.5005
R56032 VINP.n262 VINP.n87 4.5005
R56033 VINP.n308 VINP.n87 4.5005
R56034 VINP.n261 VINP.n87 4.5005
R56035 VINP.n310 VINP.n87 4.5005
R56036 VINP.n260 VINP.n87 4.5005
R56037 VINP.n312 VINP.n87 4.5005
R56038 VINP.n259 VINP.n87 4.5005
R56039 VINP.n314 VINP.n87 4.5005
R56040 VINP.n258 VINP.n87 4.5005
R56041 VINP.n316 VINP.n87 4.5005
R56042 VINP.n257 VINP.n87 4.5005
R56043 VINP.n318 VINP.n87 4.5005
R56044 VINP.n256 VINP.n87 4.5005
R56045 VINP.n320 VINP.n87 4.5005
R56046 VINP.n255 VINP.n87 4.5005
R56047 VINP.n322 VINP.n87 4.5005
R56048 VINP.n254 VINP.n87 4.5005
R56049 VINP.n324 VINP.n87 4.5005
R56050 VINP.n253 VINP.n87 4.5005
R56051 VINP.n326 VINP.n87 4.5005
R56052 VINP.n252 VINP.n87 4.5005
R56053 VINP.n328 VINP.n87 4.5005
R56054 VINP.n251 VINP.n87 4.5005
R56055 VINP.n330 VINP.n87 4.5005
R56056 VINP.n250 VINP.n87 4.5005
R56057 VINP.n332 VINP.n87 4.5005
R56058 VINP.n249 VINP.n87 4.5005
R56059 VINP.n334 VINP.n87 4.5005
R56060 VINP.n248 VINP.n87 4.5005
R56061 VINP.n336 VINP.n87 4.5005
R56062 VINP.n247 VINP.n87 4.5005
R56063 VINP.n338 VINP.n87 4.5005
R56064 VINP.n246 VINP.n87 4.5005
R56065 VINP.n340 VINP.n87 4.5005
R56066 VINP.n245 VINP.n87 4.5005
R56067 VINP.n342 VINP.n87 4.5005
R56068 VINP.n244 VINP.n87 4.5005
R56069 VINP.n344 VINP.n87 4.5005
R56070 VINP.n243 VINP.n87 4.5005
R56071 VINP.n346 VINP.n87 4.5005
R56072 VINP.n242 VINP.n87 4.5005
R56073 VINP.n348 VINP.n87 4.5005
R56074 VINP.n241 VINP.n87 4.5005
R56075 VINP.n350 VINP.n87 4.5005
R56076 VINP.n240 VINP.n87 4.5005
R56077 VINP.n352 VINP.n87 4.5005
R56078 VINP.n239 VINP.n87 4.5005
R56079 VINP.n354 VINP.n87 4.5005
R56080 VINP.n238 VINP.n87 4.5005
R56081 VINP.n356 VINP.n87 4.5005
R56082 VINP.n237 VINP.n87 4.5005
R56083 VINP.n358 VINP.n87 4.5005
R56084 VINP.n236 VINP.n87 4.5005
R56085 VINP.n360 VINP.n87 4.5005
R56086 VINP.n235 VINP.n87 4.5005
R56087 VINP.n362 VINP.n87 4.5005
R56088 VINP.n234 VINP.n87 4.5005
R56089 VINP.n364 VINP.n87 4.5005
R56090 VINP.n233 VINP.n87 4.5005
R56091 VINP.n366 VINP.n87 4.5005
R56092 VINP.n232 VINP.n87 4.5005
R56093 VINP.n368 VINP.n87 4.5005
R56094 VINP.n231 VINP.n87 4.5005
R56095 VINP.n370 VINP.n87 4.5005
R56096 VINP.n230 VINP.n87 4.5005
R56097 VINP.n372 VINP.n87 4.5005
R56098 VINP.n229 VINP.n87 4.5005
R56099 VINP.n374 VINP.n87 4.5005
R56100 VINP.n228 VINP.n87 4.5005
R56101 VINP.n376 VINP.n87 4.5005
R56102 VINP.n227 VINP.n87 4.5005
R56103 VINP.n378 VINP.n87 4.5005
R56104 VINP.n226 VINP.n87 4.5005
R56105 VINP.n380 VINP.n87 4.5005
R56106 VINP.n225 VINP.n87 4.5005
R56107 VINP.n382 VINP.n87 4.5005
R56108 VINP.n224 VINP.n87 4.5005
R56109 VINP.n384 VINP.n87 4.5005
R56110 VINP.n223 VINP.n87 4.5005
R56111 VINP.n386 VINP.n87 4.5005
R56112 VINP.n222 VINP.n87 4.5005
R56113 VINP.n388 VINP.n87 4.5005
R56114 VINP.n221 VINP.n87 4.5005
R56115 VINP.n390 VINP.n87 4.5005
R56116 VINP.n220 VINP.n87 4.5005
R56117 VINP.n392 VINP.n87 4.5005
R56118 VINP.n219 VINP.n87 4.5005
R56119 VINP.n394 VINP.n87 4.5005
R56120 VINP.n218 VINP.n87 4.5005
R56121 VINP.n396 VINP.n87 4.5005
R56122 VINP.n217 VINP.n87 4.5005
R56123 VINP.n398 VINP.n87 4.5005
R56124 VINP.n216 VINP.n87 4.5005
R56125 VINP.n400 VINP.n87 4.5005
R56126 VINP.n215 VINP.n87 4.5005
R56127 VINP.n654 VINP.n87 4.5005
R56128 VINP.n656 VINP.n87 4.5005
R56129 VINP.n87 VINP.n0 4.5005
R56130 VINP.n655 VINP.n278 4.5005
R56131 VINP.n655 VINP.n276 4.5005
R56132 VINP.n655 VINP.n280 4.5005
R56133 VINP.n655 VINP.n275 4.5005
R56134 VINP.n655 VINP.n282 4.5005
R56135 VINP.n655 VINP.n274 4.5005
R56136 VINP.n655 VINP.n284 4.5005
R56137 VINP.n655 VINP.n273 4.5005
R56138 VINP.n655 VINP.n286 4.5005
R56139 VINP.n655 VINP.n272 4.5005
R56140 VINP.n655 VINP.n288 4.5005
R56141 VINP.n655 VINP.n271 4.5005
R56142 VINP.n655 VINP.n290 4.5005
R56143 VINP.n655 VINP.n270 4.5005
R56144 VINP.n655 VINP.n292 4.5005
R56145 VINP.n655 VINP.n269 4.5005
R56146 VINP.n655 VINP.n294 4.5005
R56147 VINP.n655 VINP.n268 4.5005
R56148 VINP.n655 VINP.n296 4.5005
R56149 VINP.n655 VINP.n267 4.5005
R56150 VINP.n655 VINP.n298 4.5005
R56151 VINP.n655 VINP.n266 4.5005
R56152 VINP.n655 VINP.n300 4.5005
R56153 VINP.n655 VINP.n265 4.5005
R56154 VINP.n655 VINP.n302 4.5005
R56155 VINP.n655 VINP.n264 4.5005
R56156 VINP.n655 VINP.n304 4.5005
R56157 VINP.n655 VINP.n263 4.5005
R56158 VINP.n655 VINP.n306 4.5005
R56159 VINP.n655 VINP.n262 4.5005
R56160 VINP.n655 VINP.n308 4.5005
R56161 VINP.n655 VINP.n261 4.5005
R56162 VINP.n655 VINP.n310 4.5005
R56163 VINP.n655 VINP.n260 4.5005
R56164 VINP.n655 VINP.n312 4.5005
R56165 VINP.n655 VINP.n259 4.5005
R56166 VINP.n655 VINP.n314 4.5005
R56167 VINP.n655 VINP.n258 4.5005
R56168 VINP.n655 VINP.n316 4.5005
R56169 VINP.n655 VINP.n257 4.5005
R56170 VINP.n655 VINP.n318 4.5005
R56171 VINP.n655 VINP.n256 4.5005
R56172 VINP.n655 VINP.n320 4.5005
R56173 VINP.n655 VINP.n255 4.5005
R56174 VINP.n655 VINP.n322 4.5005
R56175 VINP.n655 VINP.n254 4.5005
R56176 VINP.n655 VINP.n324 4.5005
R56177 VINP.n655 VINP.n253 4.5005
R56178 VINP.n655 VINP.n326 4.5005
R56179 VINP.n655 VINP.n252 4.5005
R56180 VINP.n655 VINP.n328 4.5005
R56181 VINP.n655 VINP.n251 4.5005
R56182 VINP.n655 VINP.n330 4.5005
R56183 VINP.n655 VINP.n250 4.5005
R56184 VINP.n655 VINP.n332 4.5005
R56185 VINP.n655 VINP.n249 4.5005
R56186 VINP.n655 VINP.n334 4.5005
R56187 VINP.n655 VINP.n248 4.5005
R56188 VINP.n655 VINP.n336 4.5005
R56189 VINP.n655 VINP.n247 4.5005
R56190 VINP.n655 VINP.n338 4.5005
R56191 VINP.n655 VINP.n246 4.5005
R56192 VINP.n655 VINP.n340 4.5005
R56193 VINP.n655 VINP.n245 4.5005
R56194 VINP.n655 VINP.n342 4.5005
R56195 VINP.n655 VINP.n244 4.5005
R56196 VINP.n655 VINP.n344 4.5005
R56197 VINP.n655 VINP.n243 4.5005
R56198 VINP.n655 VINP.n346 4.5005
R56199 VINP.n655 VINP.n242 4.5005
R56200 VINP.n655 VINP.n348 4.5005
R56201 VINP.n655 VINP.n241 4.5005
R56202 VINP.n655 VINP.n350 4.5005
R56203 VINP.n655 VINP.n240 4.5005
R56204 VINP.n655 VINP.n352 4.5005
R56205 VINP.n655 VINP.n239 4.5005
R56206 VINP.n655 VINP.n354 4.5005
R56207 VINP.n655 VINP.n238 4.5005
R56208 VINP.n655 VINP.n356 4.5005
R56209 VINP.n655 VINP.n237 4.5005
R56210 VINP.n655 VINP.n358 4.5005
R56211 VINP.n655 VINP.n236 4.5005
R56212 VINP.n655 VINP.n360 4.5005
R56213 VINP.n655 VINP.n235 4.5005
R56214 VINP.n655 VINP.n362 4.5005
R56215 VINP.n655 VINP.n234 4.5005
R56216 VINP.n655 VINP.n364 4.5005
R56217 VINP.n655 VINP.n233 4.5005
R56218 VINP.n655 VINP.n366 4.5005
R56219 VINP.n655 VINP.n232 4.5005
R56220 VINP.n655 VINP.n368 4.5005
R56221 VINP.n655 VINP.n231 4.5005
R56222 VINP.n655 VINP.n370 4.5005
R56223 VINP.n655 VINP.n230 4.5005
R56224 VINP.n655 VINP.n372 4.5005
R56225 VINP.n655 VINP.n229 4.5005
R56226 VINP.n655 VINP.n374 4.5005
R56227 VINP.n655 VINP.n228 4.5005
R56228 VINP.n655 VINP.n376 4.5005
R56229 VINP.n655 VINP.n227 4.5005
R56230 VINP.n655 VINP.n378 4.5005
R56231 VINP.n655 VINP.n226 4.5005
R56232 VINP.n655 VINP.n380 4.5005
R56233 VINP.n655 VINP.n225 4.5005
R56234 VINP.n655 VINP.n382 4.5005
R56235 VINP.n655 VINP.n224 4.5005
R56236 VINP.n655 VINP.n384 4.5005
R56237 VINP.n655 VINP.n223 4.5005
R56238 VINP.n655 VINP.n386 4.5005
R56239 VINP.n655 VINP.n222 4.5005
R56240 VINP.n655 VINP.n388 4.5005
R56241 VINP.n655 VINP.n221 4.5005
R56242 VINP.n655 VINP.n390 4.5005
R56243 VINP.n655 VINP.n220 4.5005
R56244 VINP.n655 VINP.n392 4.5005
R56245 VINP.n655 VINP.n219 4.5005
R56246 VINP.n655 VINP.n394 4.5005
R56247 VINP.n655 VINP.n218 4.5005
R56248 VINP.n655 VINP.n396 4.5005
R56249 VINP.n655 VINP.n217 4.5005
R56250 VINP.n655 VINP.n398 4.5005
R56251 VINP.n655 VINP.n216 4.5005
R56252 VINP.n655 VINP.n400 4.5005
R56253 VINP.n655 VINP.n215 4.5005
R56254 VINP.n655 VINP.n654 4.5005
R56255 VINP.n656 VINP.n655 4.5005
R56256 VINP.n655 VINP.n0 4.5005
R56257 VINP.n278 VINP.n86 4.5005
R56258 VINP.n276 VINP.n86 4.5005
R56259 VINP.n280 VINP.n86 4.5005
R56260 VINP.n275 VINP.n86 4.5005
R56261 VINP.n282 VINP.n86 4.5005
R56262 VINP.n274 VINP.n86 4.5005
R56263 VINP.n284 VINP.n86 4.5005
R56264 VINP.n273 VINP.n86 4.5005
R56265 VINP.n286 VINP.n86 4.5005
R56266 VINP.n272 VINP.n86 4.5005
R56267 VINP.n288 VINP.n86 4.5005
R56268 VINP.n271 VINP.n86 4.5005
R56269 VINP.n290 VINP.n86 4.5005
R56270 VINP.n270 VINP.n86 4.5005
R56271 VINP.n292 VINP.n86 4.5005
R56272 VINP.n269 VINP.n86 4.5005
R56273 VINP.n294 VINP.n86 4.5005
R56274 VINP.n268 VINP.n86 4.5005
R56275 VINP.n296 VINP.n86 4.5005
R56276 VINP.n267 VINP.n86 4.5005
R56277 VINP.n298 VINP.n86 4.5005
R56278 VINP.n266 VINP.n86 4.5005
R56279 VINP.n300 VINP.n86 4.5005
R56280 VINP.n265 VINP.n86 4.5005
R56281 VINP.n302 VINP.n86 4.5005
R56282 VINP.n264 VINP.n86 4.5005
R56283 VINP.n304 VINP.n86 4.5005
R56284 VINP.n263 VINP.n86 4.5005
R56285 VINP.n306 VINP.n86 4.5005
R56286 VINP.n262 VINP.n86 4.5005
R56287 VINP.n308 VINP.n86 4.5005
R56288 VINP.n261 VINP.n86 4.5005
R56289 VINP.n310 VINP.n86 4.5005
R56290 VINP.n260 VINP.n86 4.5005
R56291 VINP.n312 VINP.n86 4.5005
R56292 VINP.n259 VINP.n86 4.5005
R56293 VINP.n314 VINP.n86 4.5005
R56294 VINP.n258 VINP.n86 4.5005
R56295 VINP.n316 VINP.n86 4.5005
R56296 VINP.n257 VINP.n86 4.5005
R56297 VINP.n318 VINP.n86 4.5005
R56298 VINP.n256 VINP.n86 4.5005
R56299 VINP.n320 VINP.n86 4.5005
R56300 VINP.n255 VINP.n86 4.5005
R56301 VINP.n322 VINP.n86 4.5005
R56302 VINP.n254 VINP.n86 4.5005
R56303 VINP.n324 VINP.n86 4.5005
R56304 VINP.n253 VINP.n86 4.5005
R56305 VINP.n326 VINP.n86 4.5005
R56306 VINP.n252 VINP.n86 4.5005
R56307 VINP.n328 VINP.n86 4.5005
R56308 VINP.n251 VINP.n86 4.5005
R56309 VINP.n330 VINP.n86 4.5005
R56310 VINP.n250 VINP.n86 4.5005
R56311 VINP.n332 VINP.n86 4.5005
R56312 VINP.n249 VINP.n86 4.5005
R56313 VINP.n334 VINP.n86 4.5005
R56314 VINP.n248 VINP.n86 4.5005
R56315 VINP.n336 VINP.n86 4.5005
R56316 VINP.n247 VINP.n86 4.5005
R56317 VINP.n338 VINP.n86 4.5005
R56318 VINP.n246 VINP.n86 4.5005
R56319 VINP.n340 VINP.n86 4.5005
R56320 VINP.n245 VINP.n86 4.5005
R56321 VINP.n342 VINP.n86 4.5005
R56322 VINP.n244 VINP.n86 4.5005
R56323 VINP.n344 VINP.n86 4.5005
R56324 VINP.n243 VINP.n86 4.5005
R56325 VINP.n346 VINP.n86 4.5005
R56326 VINP.n242 VINP.n86 4.5005
R56327 VINP.n348 VINP.n86 4.5005
R56328 VINP.n241 VINP.n86 4.5005
R56329 VINP.n350 VINP.n86 4.5005
R56330 VINP.n240 VINP.n86 4.5005
R56331 VINP.n352 VINP.n86 4.5005
R56332 VINP.n239 VINP.n86 4.5005
R56333 VINP.n354 VINP.n86 4.5005
R56334 VINP.n238 VINP.n86 4.5005
R56335 VINP.n356 VINP.n86 4.5005
R56336 VINP.n237 VINP.n86 4.5005
R56337 VINP.n358 VINP.n86 4.5005
R56338 VINP.n236 VINP.n86 4.5005
R56339 VINP.n360 VINP.n86 4.5005
R56340 VINP.n235 VINP.n86 4.5005
R56341 VINP.n362 VINP.n86 4.5005
R56342 VINP.n234 VINP.n86 4.5005
R56343 VINP.n364 VINP.n86 4.5005
R56344 VINP.n233 VINP.n86 4.5005
R56345 VINP.n366 VINP.n86 4.5005
R56346 VINP.n232 VINP.n86 4.5005
R56347 VINP.n368 VINP.n86 4.5005
R56348 VINP.n231 VINP.n86 4.5005
R56349 VINP.n370 VINP.n86 4.5005
R56350 VINP.n230 VINP.n86 4.5005
R56351 VINP.n372 VINP.n86 4.5005
R56352 VINP.n229 VINP.n86 4.5005
R56353 VINP.n374 VINP.n86 4.5005
R56354 VINP.n228 VINP.n86 4.5005
R56355 VINP.n376 VINP.n86 4.5005
R56356 VINP.n227 VINP.n86 4.5005
R56357 VINP.n378 VINP.n86 4.5005
R56358 VINP.n226 VINP.n86 4.5005
R56359 VINP.n380 VINP.n86 4.5005
R56360 VINP.n225 VINP.n86 4.5005
R56361 VINP.n382 VINP.n86 4.5005
R56362 VINP.n224 VINP.n86 4.5005
R56363 VINP.n384 VINP.n86 4.5005
R56364 VINP.n223 VINP.n86 4.5005
R56365 VINP.n386 VINP.n86 4.5005
R56366 VINP.n222 VINP.n86 4.5005
R56367 VINP.n388 VINP.n86 4.5005
R56368 VINP.n221 VINP.n86 4.5005
R56369 VINP.n390 VINP.n86 4.5005
R56370 VINP.n220 VINP.n86 4.5005
R56371 VINP.n392 VINP.n86 4.5005
R56372 VINP.n219 VINP.n86 4.5005
R56373 VINP.n394 VINP.n86 4.5005
R56374 VINP.n218 VINP.n86 4.5005
R56375 VINP.n396 VINP.n86 4.5005
R56376 VINP.n217 VINP.n86 4.5005
R56377 VINP.n398 VINP.n86 4.5005
R56378 VINP.n216 VINP.n86 4.5005
R56379 VINP.n400 VINP.n86 4.5005
R56380 VINP.n215 VINP.n86 4.5005
R56381 VINP.n654 VINP.n86 4.5005
R56382 VINP.n528 VINP.n86 4.5005
R56383 VINP.n656 VINP.n86 4.5005
R56384 VINP.n86 VINP.n0 4.5005
R56385 VINP.n462 VINP.n278 2.25083
R56386 VINP.n463 VINP.n461 2.25083
R56387 VINP.n463 VINP.n460 2.25083
R56388 VINP.n463 VINP.n459 2.25083
R56389 VINP.n463 VINP.n458 2.25083
R56390 VINP.n463 VINP.n457 2.25083
R56391 VINP.n463 VINP.n456 2.25083
R56392 VINP.n463 VINP.n455 2.25083
R56393 VINP.n463 VINP.n454 2.25083
R56394 VINP.n463 VINP.n453 2.25083
R56395 VINP.n463 VINP.n452 2.25083
R56396 VINP.n463 VINP.n451 2.25083
R56397 VINP.n463 VINP.n450 2.25083
R56398 VINP.n463 VINP.n449 2.25083
R56399 VINP.n463 VINP.n448 2.25083
R56400 VINP.n463 VINP.n447 2.25083
R56401 VINP.n463 VINP.n446 2.25083
R56402 VINP.n463 VINP.n445 2.25083
R56403 VINP.n463 VINP.n444 2.25083
R56404 VINP.n463 VINP.n443 2.25083
R56405 VINP.n463 VINP.n442 2.25083
R56406 VINP.n463 VINP.n441 2.25083
R56407 VINP.n463 VINP.n440 2.25083
R56408 VINP.n463 VINP.n439 2.25083
R56409 VINP.n463 VINP.n438 2.25083
R56410 VINP.n463 VINP.n437 2.25083
R56411 VINP.n463 VINP.n436 2.25083
R56412 VINP.n463 VINP.n435 2.25083
R56413 VINP.n463 VINP.n434 2.25083
R56414 VINP.n463 VINP.n433 2.25083
R56415 VINP.n463 VINP.n432 2.25083
R56416 VINP.n463 VINP.n431 2.25083
R56417 VINP.n463 VINP.n430 2.25083
R56418 VINP.n463 VINP.n429 2.25083
R56419 VINP.n463 VINP.n428 2.25083
R56420 VINP.n463 VINP.n427 2.25083
R56421 VINP.n463 VINP.n426 2.25083
R56422 VINP.n463 VINP.n425 2.25083
R56423 VINP.n463 VINP.n424 2.25083
R56424 VINP.n463 VINP.n423 2.25083
R56425 VINP.n463 VINP.n422 2.25083
R56426 VINP.n463 VINP.n421 2.25083
R56427 VINP.n463 VINP.n420 2.25083
R56428 VINP.n463 VINP.n419 2.25083
R56429 VINP.n463 VINP.n418 2.25083
R56430 VINP.n463 VINP.n417 2.25083
R56431 VINP.n463 VINP.n416 2.25083
R56432 VINP.n463 VINP.n415 2.25083
R56433 VINP.n463 VINP.n414 2.25083
R56434 VINP.n463 VINP.n413 2.25083
R56435 VINP.n463 VINP.n412 2.25083
R56436 VINP.n463 VINP.n411 2.25083
R56437 VINP.n463 VINP.n410 2.25083
R56438 VINP.n463 VINP.n409 2.25083
R56439 VINP.n463 VINP.n408 2.25083
R56440 VINP.n463 VINP.n407 2.25083
R56441 VINP.n463 VINP.n406 2.25083
R56442 VINP.n463 VINP.n405 2.25083
R56443 VINP.n463 VINP.n404 2.25083
R56444 VINP.n463 VINP.n403 2.25083
R56445 VINP.n463 VINP.n402 2.25083
R56446 VINP.n463 VINP.n401 2.25083
R56447 VINP.n464 VINP.n463 2.25083
R56448 VINP.n463 VINP.n150 2.25083
R56449 VINP.n463 VINP.n66 2.25083
R56450 VINP.n279 VINP.n151 2.25083
R56451 VINP.n281 VINP.n151 2.25083
R56452 VINP.n283 VINP.n151 2.25083
R56453 VINP.n285 VINP.n151 2.25083
R56454 VINP.n287 VINP.n151 2.25083
R56455 VINP.n289 VINP.n151 2.25083
R56456 VINP.n291 VINP.n151 2.25083
R56457 VINP.n293 VINP.n151 2.25083
R56458 VINP.n295 VINP.n151 2.25083
R56459 VINP.n297 VINP.n151 2.25083
R56460 VINP.n299 VINP.n151 2.25083
R56461 VINP.n301 VINP.n151 2.25083
R56462 VINP.n303 VINP.n151 2.25083
R56463 VINP.n305 VINP.n151 2.25083
R56464 VINP.n307 VINP.n151 2.25083
R56465 VINP.n309 VINP.n151 2.25083
R56466 VINP.n311 VINP.n151 2.25083
R56467 VINP.n313 VINP.n151 2.25083
R56468 VINP.n315 VINP.n151 2.25083
R56469 VINP.n317 VINP.n151 2.25083
R56470 VINP.n319 VINP.n151 2.25083
R56471 VINP.n321 VINP.n151 2.25083
R56472 VINP.n323 VINP.n151 2.25083
R56473 VINP.n325 VINP.n151 2.25083
R56474 VINP.n327 VINP.n151 2.25083
R56475 VINP.n329 VINP.n151 2.25083
R56476 VINP.n331 VINP.n151 2.25083
R56477 VINP.n333 VINP.n151 2.25083
R56478 VINP.n335 VINP.n151 2.25083
R56479 VINP.n337 VINP.n151 2.25083
R56480 VINP.n339 VINP.n151 2.25083
R56481 VINP.n341 VINP.n151 2.25083
R56482 VINP.n343 VINP.n151 2.25083
R56483 VINP.n345 VINP.n151 2.25083
R56484 VINP.n347 VINP.n151 2.25083
R56485 VINP.n349 VINP.n151 2.25083
R56486 VINP.n351 VINP.n151 2.25083
R56487 VINP.n353 VINP.n151 2.25083
R56488 VINP.n355 VINP.n151 2.25083
R56489 VINP.n357 VINP.n151 2.25083
R56490 VINP.n359 VINP.n151 2.25083
R56491 VINP.n361 VINP.n151 2.25083
R56492 VINP.n363 VINP.n151 2.25083
R56493 VINP.n365 VINP.n151 2.25083
R56494 VINP.n367 VINP.n151 2.25083
R56495 VINP.n369 VINP.n151 2.25083
R56496 VINP.n371 VINP.n151 2.25083
R56497 VINP.n373 VINP.n151 2.25083
R56498 VINP.n375 VINP.n151 2.25083
R56499 VINP.n377 VINP.n151 2.25083
R56500 VINP.n379 VINP.n151 2.25083
R56501 VINP.n381 VINP.n151 2.25083
R56502 VINP.n383 VINP.n151 2.25083
R56503 VINP.n385 VINP.n151 2.25083
R56504 VINP.n387 VINP.n151 2.25083
R56505 VINP.n389 VINP.n151 2.25083
R56506 VINP.n391 VINP.n151 2.25083
R56507 VINP.n393 VINP.n151 2.25083
R56508 VINP.n395 VINP.n151 2.25083
R56509 VINP.n397 VINP.n151 2.25083
R56510 VINP.n399 VINP.n151 2.25083
R56511 VINP.n465 VINP.n151 2.25083
R56512 VINP.n277 VINP.n149 2.25083
R56513 VINP.n657 VINP.n65 2.25083
R56514 VINP.n528 VINP.n466 2.25083
R56515 VINP.n657 VINP.n64 2.25083
R56516 VINP.n528 VINP.n467 2.25083
R56517 VINP.n657 VINP.n63 2.25083
R56518 VINP.n528 VINP.n468 2.25083
R56519 VINP.n657 VINP.n62 2.25083
R56520 VINP.n528 VINP.n469 2.25083
R56521 VINP.n657 VINP.n61 2.25083
R56522 VINP.n528 VINP.n470 2.25083
R56523 VINP.n657 VINP.n60 2.25083
R56524 VINP.n528 VINP.n471 2.25083
R56525 VINP.n657 VINP.n59 2.25083
R56526 VINP.n528 VINP.n472 2.25083
R56527 VINP.n657 VINP.n58 2.25083
R56528 VINP.n528 VINP.n473 2.25083
R56529 VINP.n657 VINP.n57 2.25083
R56530 VINP.n528 VINP.n474 2.25083
R56531 VINP.n657 VINP.n56 2.25083
R56532 VINP.n528 VINP.n475 2.25083
R56533 VINP.n657 VINP.n55 2.25083
R56534 VINP.n528 VINP.n476 2.25083
R56535 VINP.n657 VINP.n54 2.25083
R56536 VINP.n528 VINP.n477 2.25083
R56537 VINP.n657 VINP.n53 2.25083
R56538 VINP.n528 VINP.n478 2.25083
R56539 VINP.n657 VINP.n52 2.25083
R56540 VINP.n528 VINP.n479 2.25083
R56541 VINP.n657 VINP.n51 2.25083
R56542 VINP.n528 VINP.n480 2.25083
R56543 VINP.n657 VINP.n50 2.25083
R56544 VINP.n528 VINP.n481 2.25083
R56545 VINP.n657 VINP.n49 2.25083
R56546 VINP.n528 VINP.n482 2.25083
R56547 VINP.n657 VINP.n48 2.25083
R56548 VINP.n528 VINP.n483 2.25083
R56549 VINP.n657 VINP.n47 2.25083
R56550 VINP.n528 VINP.n484 2.25083
R56551 VINP.n657 VINP.n46 2.25083
R56552 VINP.n528 VINP.n485 2.25083
R56553 VINP.n657 VINP.n45 2.25083
R56554 VINP.n528 VINP.n486 2.25083
R56555 VINP.n657 VINP.n44 2.25083
R56556 VINP.n528 VINP.n487 2.25083
R56557 VINP.n657 VINP.n43 2.25083
R56558 VINP.n528 VINP.n488 2.25083
R56559 VINP.n657 VINP.n42 2.25083
R56560 VINP.n528 VINP.n489 2.25083
R56561 VINP.n657 VINP.n41 2.25083
R56562 VINP.n528 VINP.n490 2.25083
R56563 VINP.n657 VINP.n40 2.25083
R56564 VINP.n528 VINP.n491 2.25083
R56565 VINP.n657 VINP.n39 2.25083
R56566 VINP.n528 VINP.n492 2.25083
R56567 VINP.n657 VINP.n38 2.25083
R56568 VINP.n528 VINP.n493 2.25083
R56569 VINP.n657 VINP.n37 2.25083
R56570 VINP.n528 VINP.n494 2.25083
R56571 VINP.n657 VINP.n36 2.25083
R56572 VINP.n528 VINP.n495 2.25083
R56573 VINP.n657 VINP.n35 2.25083
R56574 VINP.n528 VINP.n496 2.25083
R56575 VINP.n657 VINP.n34 2.25083
R56576 VINP.n528 VINP.n497 2.25083
R56577 VINP.n657 VINP.n33 2.25083
R56578 VINP.n528 VINP.n498 2.25083
R56579 VINP.n657 VINP.n32 2.25083
R56580 VINP.n528 VINP.n499 2.25083
R56581 VINP.n657 VINP.n31 2.25083
R56582 VINP.n528 VINP.n500 2.25083
R56583 VINP.n657 VINP.n30 2.25083
R56584 VINP.n528 VINP.n501 2.25083
R56585 VINP.n657 VINP.n29 2.25083
R56586 VINP.n528 VINP.n502 2.25083
R56587 VINP.n657 VINP.n28 2.25083
R56588 VINP.n528 VINP.n503 2.25083
R56589 VINP.n657 VINP.n27 2.25083
R56590 VINP.n528 VINP.n504 2.25083
R56591 VINP.n657 VINP.n26 2.25083
R56592 VINP.n528 VINP.n505 2.25083
R56593 VINP.n657 VINP.n25 2.25083
R56594 VINP.n528 VINP.n506 2.25083
R56595 VINP.n657 VINP.n24 2.25083
R56596 VINP.n528 VINP.n507 2.25083
R56597 VINP.n657 VINP.n23 2.25083
R56598 VINP.n528 VINP.n508 2.25083
R56599 VINP.n657 VINP.n22 2.25083
R56600 VINP.n528 VINP.n509 2.25083
R56601 VINP.n657 VINP.n21 2.25083
R56602 VINP.n528 VINP.n510 2.25083
R56603 VINP.n657 VINP.n20 2.25083
R56604 VINP.n528 VINP.n511 2.25083
R56605 VINP.n657 VINP.n19 2.25083
R56606 VINP.n528 VINP.n512 2.25083
R56607 VINP.n657 VINP.n18 2.25083
R56608 VINP.n528 VINP.n513 2.25083
R56609 VINP.n657 VINP.n17 2.25083
R56610 VINP.n528 VINP.n514 2.25083
R56611 VINP.n657 VINP.n16 2.25083
R56612 VINP.n528 VINP.n515 2.25083
R56613 VINP.n657 VINP.n15 2.25083
R56614 VINP.n528 VINP.n516 2.25083
R56615 VINP.n657 VINP.n14 2.25083
R56616 VINP.n528 VINP.n517 2.25083
R56617 VINP.n657 VINP.n13 2.25083
R56618 VINP.n528 VINP.n518 2.25083
R56619 VINP.n657 VINP.n12 2.25083
R56620 VINP.n528 VINP.n519 2.25083
R56621 VINP.n657 VINP.n11 2.25083
R56622 VINP.n528 VINP.n520 2.25083
R56623 VINP.n657 VINP.n10 2.25083
R56624 VINP.n528 VINP.n521 2.25083
R56625 VINP.n657 VINP.n9 2.25083
R56626 VINP.n528 VINP.n522 2.25083
R56627 VINP.n657 VINP.n8 2.25083
R56628 VINP.n528 VINP.n523 2.25083
R56629 VINP.n657 VINP.n7 2.25083
R56630 VINP.n528 VINP.n524 2.25083
R56631 VINP.n657 VINP.n6 2.25083
R56632 VINP.n528 VINP.n525 2.25083
R56633 VINP.n657 VINP.n5 2.25083
R56634 VINP.n528 VINP.n526 2.25083
R56635 VINP.n657 VINP.n4 2.25083
R56636 VINP.n528 VINP.n527 2.25083
R56637 VINP.n657 VINP.n3 2.25083
R56638 VINP.n528 VINP.n214 2.25083
R56639 VINP.n657 VINP.n2 2.25083
R56640 VINP.n85 VINP.n84 0.0977
R56641 VINP.n84 VINP.n83 0.0977
R56642 VINP.n83 VINP.n82 0.0977
R56643 VINP.n82 VINP.n81 0.0977
R56644 VINP.n81 VINP.n80 0.0977
R56645 VINP.n80 VINP.n79 0.0977
R56646 VINP.n79 VINP.n78 0.0977
R56647 VINP.n78 VINP.n77 0.0977
R56648 VINP.n77 VINP.n76 0.0977
R56649 VINP.n76 VINP.n75 0.0977
R56650 VINP.n75 VINP.n74 0.0977
R56651 VINP.n74 VINP.n73 0.0977
R56652 VINP.n73 VINP.n72 0.0977
R56653 VINP.n72 VINP.n71 0.0977
R56654 VINP.n71 VINP.n70 0.0977
R56655 VINP.n70 VINP.n69 0.0977
R56656 VINP.n69 VINP.n68 0.0977
R56657 VINP.n68 VINP.n67 0.0977
R56658 VINP.n658 VINP.n0 0.0358487
R56659 VINP.n530 VINP.n278 0.0358487
R56660 VINP.n658 VINP.n657 0.0353837
R56661 VINP.n656 VINP.n1 0.0353837
R56662 VINP.n529 VINP.n528 0.0353837
R56663 VINP.n654 VINP.n653 0.0353837
R56664 VINP.n652 VINP.n215 0.0353837
R56665 VINP.n651 VINP.n400 0.0353837
R56666 VINP.n650 VINP.n216 0.0353837
R56667 VINP.n649 VINP.n398 0.0353837
R56668 VINP.n648 VINP.n217 0.0353837
R56669 VINP.n647 VINP.n396 0.0353837
R56670 VINP.n646 VINP.n218 0.0353837
R56671 VINP.n645 VINP.n394 0.0353837
R56672 VINP.n644 VINP.n219 0.0353837
R56673 VINP.n643 VINP.n392 0.0353837
R56674 VINP.n642 VINP.n220 0.0353837
R56675 VINP.n641 VINP.n390 0.0353837
R56676 VINP.n640 VINP.n221 0.0353837
R56677 VINP.n639 VINP.n388 0.0353837
R56678 VINP.n638 VINP.n222 0.0353837
R56679 VINP.n637 VINP.n386 0.0353837
R56680 VINP.n636 VINP.n223 0.0353837
R56681 VINP.n635 VINP.n384 0.0353837
R56682 VINP.n634 VINP.n224 0.0353837
R56683 VINP.n633 VINP.n382 0.0353837
R56684 VINP.n632 VINP.n225 0.0353837
R56685 VINP.n631 VINP.n380 0.0353837
R56686 VINP.n630 VINP.n226 0.0353837
R56687 VINP.n629 VINP.n378 0.0353837
R56688 VINP.n628 VINP.n227 0.0353837
R56689 VINP.n627 VINP.n376 0.0353837
R56690 VINP.n626 VINP.n228 0.0353837
R56691 VINP.n625 VINP.n374 0.0353837
R56692 VINP.n624 VINP.n229 0.0353837
R56693 VINP.n623 VINP.n372 0.0353837
R56694 VINP.n622 VINP.n230 0.0353837
R56695 VINP.n621 VINP.n370 0.0353837
R56696 VINP.n620 VINP.n231 0.0353837
R56697 VINP.n619 VINP.n368 0.0353837
R56698 VINP.n618 VINP.n232 0.0353837
R56699 VINP.n617 VINP.n366 0.0353837
R56700 VINP.n616 VINP.n233 0.0353837
R56701 VINP.n615 VINP.n364 0.0353837
R56702 VINP.n614 VINP.n234 0.0353837
R56703 VINP.n613 VINP.n362 0.0353837
R56704 VINP.n612 VINP.n235 0.0353837
R56705 VINP.n611 VINP.n360 0.0353837
R56706 VINP.n610 VINP.n236 0.0353837
R56707 VINP.n609 VINP.n358 0.0353837
R56708 VINP.n608 VINP.n237 0.0353837
R56709 VINP.n607 VINP.n356 0.0353837
R56710 VINP.n606 VINP.n238 0.0353837
R56711 VINP.n605 VINP.n354 0.0353837
R56712 VINP.n604 VINP.n239 0.0353837
R56713 VINP.n603 VINP.n352 0.0353837
R56714 VINP.n602 VINP.n240 0.0353837
R56715 VINP.n601 VINP.n350 0.0353837
R56716 VINP.n600 VINP.n241 0.0353837
R56717 VINP.n599 VINP.n348 0.0353837
R56718 VINP.n598 VINP.n242 0.0353837
R56719 VINP.n597 VINP.n346 0.0353837
R56720 VINP.n596 VINP.n243 0.0353837
R56721 VINP.n595 VINP.n344 0.0353837
R56722 VINP.n594 VINP.n244 0.0353837
R56723 VINP.n593 VINP.n342 0.0353837
R56724 VINP.n592 VINP.n245 0.0353837
R56725 VINP.n591 VINP.n340 0.0353837
R56726 VINP.n590 VINP.n246 0.0353837
R56727 VINP.n589 VINP.n338 0.0353837
R56728 VINP.n588 VINP.n247 0.0353837
R56729 VINP.n587 VINP.n336 0.0353837
R56730 VINP.n586 VINP.n248 0.0353837
R56731 VINP.n585 VINP.n334 0.0353837
R56732 VINP.n584 VINP.n249 0.0353837
R56733 VINP.n583 VINP.n332 0.0353837
R56734 VINP.n582 VINP.n250 0.0353837
R56735 VINP.n581 VINP.n330 0.0353837
R56736 VINP.n580 VINP.n251 0.0353837
R56737 VINP.n579 VINP.n328 0.0353837
R56738 VINP.n578 VINP.n252 0.0353837
R56739 VINP.n577 VINP.n326 0.0353837
R56740 VINP.n576 VINP.n253 0.0353837
R56741 VINP.n575 VINP.n324 0.0353837
R56742 VINP.n574 VINP.n254 0.0353837
R56743 VINP.n573 VINP.n322 0.0353837
R56744 VINP.n572 VINP.n255 0.0353837
R56745 VINP.n571 VINP.n320 0.0353837
R56746 VINP.n570 VINP.n256 0.0353837
R56747 VINP.n569 VINP.n318 0.0353837
R56748 VINP.n568 VINP.n257 0.0353837
R56749 VINP.n567 VINP.n316 0.0353837
R56750 VINP.n566 VINP.n258 0.0353837
R56751 VINP.n565 VINP.n314 0.0353837
R56752 VINP.n564 VINP.n259 0.0353837
R56753 VINP.n563 VINP.n312 0.0353837
R56754 VINP.n562 VINP.n260 0.0353837
R56755 VINP.n561 VINP.n310 0.0353837
R56756 VINP.n560 VINP.n261 0.0353837
R56757 VINP.n559 VINP.n308 0.0353837
R56758 VINP.n558 VINP.n262 0.0353837
R56759 VINP.n557 VINP.n306 0.0353837
R56760 VINP.n556 VINP.n263 0.0353837
R56761 VINP.n555 VINP.n304 0.0353837
R56762 VINP.n554 VINP.n264 0.0353837
R56763 VINP.n553 VINP.n302 0.0353837
R56764 VINP.n552 VINP.n265 0.0353837
R56765 VINP.n551 VINP.n300 0.0353837
R56766 VINP.n550 VINP.n266 0.0353837
R56767 VINP.n549 VINP.n298 0.0353837
R56768 VINP.n548 VINP.n267 0.0353837
R56769 VINP.n547 VINP.n296 0.0353837
R56770 VINP.n546 VINP.n268 0.0353837
R56771 VINP.n545 VINP.n294 0.0353837
R56772 VINP.n544 VINP.n269 0.0353837
R56773 VINP.n543 VINP.n292 0.0353837
R56774 VINP.n542 VINP.n270 0.0353837
R56775 VINP.n541 VINP.n290 0.0353837
R56776 VINP.n540 VINP.n271 0.0353837
R56777 VINP.n539 VINP.n288 0.0353837
R56778 VINP.n538 VINP.n272 0.0353837
R56779 VINP.n537 VINP.n286 0.0353837
R56780 VINP.n536 VINP.n273 0.0353837
R56781 VINP.n535 VINP.n284 0.0353837
R56782 VINP.n534 VINP.n274 0.0353837
R56783 VINP.n533 VINP.n282 0.0353837
R56784 VINP.n532 VINP.n275 0.0353837
R56785 VINP.n531 VINP.n280 0.0353837
R56786 VINP.n530 VINP.n276 0.0353837
R56787 VINP.n463 VINP.n462 0.00134872
R56788 VINP.n149 VINP.n65 0.00134872
R56789 VINP.n466 VINP.n152 0.00134872
R56790 VINP.n148 VINP.n64 0.00134872
R56791 VINP.n467 VINP.n153 0.00134872
R56792 VINP.n147 VINP.n63 0.00134872
R56793 VINP.n468 VINP.n154 0.00134872
R56794 VINP.n146 VINP.n62 0.00134872
R56795 VINP.n469 VINP.n155 0.00134872
R56796 VINP.n145 VINP.n61 0.00134872
R56797 VINP.n470 VINP.n156 0.00134872
R56798 VINP.n144 VINP.n60 0.00134872
R56799 VINP.n471 VINP.n157 0.00134872
R56800 VINP.n143 VINP.n59 0.00134872
R56801 VINP.n472 VINP.n158 0.00134872
R56802 VINP.n142 VINP.n58 0.00134872
R56803 VINP.n473 VINP.n159 0.00134872
R56804 VINP.n141 VINP.n57 0.00134872
R56805 VINP.n474 VINP.n160 0.00134872
R56806 VINP.n140 VINP.n56 0.00134872
R56807 VINP.n475 VINP.n161 0.00134872
R56808 VINP.n139 VINP.n55 0.00134872
R56809 VINP.n476 VINP.n162 0.00134872
R56810 VINP.n138 VINP.n54 0.00134872
R56811 VINP.n477 VINP.n163 0.00134872
R56812 VINP.n137 VINP.n53 0.00134872
R56813 VINP.n478 VINP.n164 0.00134872
R56814 VINP.n136 VINP.n52 0.00134872
R56815 VINP.n479 VINP.n165 0.00134872
R56816 VINP.n135 VINP.n51 0.00134872
R56817 VINP.n480 VINP.n166 0.00134872
R56818 VINP.n134 VINP.n50 0.00134872
R56819 VINP.n481 VINP.n167 0.00134872
R56820 VINP.n133 VINP.n49 0.00134872
R56821 VINP.n482 VINP.n168 0.00134872
R56822 VINP.n132 VINP.n48 0.00134872
R56823 VINP.n483 VINP.n169 0.00134872
R56824 VINP.n131 VINP.n47 0.00134872
R56825 VINP.n484 VINP.n170 0.00134872
R56826 VINP.n130 VINP.n46 0.00134872
R56827 VINP.n485 VINP.n171 0.00134872
R56828 VINP.n129 VINP.n45 0.00134872
R56829 VINP.n486 VINP.n172 0.00134872
R56830 VINP.n128 VINP.n44 0.00134872
R56831 VINP.n487 VINP.n173 0.00134872
R56832 VINP.n127 VINP.n43 0.00134872
R56833 VINP.n488 VINP.n174 0.00134872
R56834 VINP.n126 VINP.n42 0.00134872
R56835 VINP.n489 VINP.n175 0.00134872
R56836 VINP.n125 VINP.n41 0.00134872
R56837 VINP.n490 VINP.n176 0.00134872
R56838 VINP.n124 VINP.n40 0.00134872
R56839 VINP.n491 VINP.n177 0.00134872
R56840 VINP.n123 VINP.n39 0.00134872
R56841 VINP.n492 VINP.n178 0.00134872
R56842 VINP.n122 VINP.n38 0.00134872
R56843 VINP.n493 VINP.n179 0.00134872
R56844 VINP.n121 VINP.n37 0.00134872
R56845 VINP.n494 VINP.n180 0.00134872
R56846 VINP.n120 VINP.n36 0.00134872
R56847 VINP.n495 VINP.n181 0.00134872
R56848 VINP.n119 VINP.n35 0.00134872
R56849 VINP.n496 VINP.n182 0.00134872
R56850 VINP.n118 VINP.n34 0.00134872
R56851 VINP.n497 VINP.n183 0.00134872
R56852 VINP.n117 VINP.n33 0.00134872
R56853 VINP.n498 VINP.n184 0.00134872
R56854 VINP.n116 VINP.n32 0.00134872
R56855 VINP.n499 VINP.n185 0.00134872
R56856 VINP.n115 VINP.n31 0.00134872
R56857 VINP.n500 VINP.n186 0.00134872
R56858 VINP.n114 VINP.n30 0.00134872
R56859 VINP.n501 VINP.n187 0.00134872
R56860 VINP.n113 VINP.n29 0.00134872
R56861 VINP.n502 VINP.n188 0.00134872
R56862 VINP.n112 VINP.n28 0.00134872
R56863 VINP.n503 VINP.n189 0.00134872
R56864 VINP.n111 VINP.n27 0.00134872
R56865 VINP.n504 VINP.n190 0.00134872
R56866 VINP.n110 VINP.n26 0.00134872
R56867 VINP.n505 VINP.n191 0.00134872
R56868 VINP.n109 VINP.n25 0.00134872
R56869 VINP.n506 VINP.n192 0.00134872
R56870 VINP.n108 VINP.n24 0.00134872
R56871 VINP.n507 VINP.n193 0.00134872
R56872 VINP.n107 VINP.n23 0.00134872
R56873 VINP.n508 VINP.n194 0.00134872
R56874 VINP.n106 VINP.n22 0.00134872
R56875 VINP.n509 VINP.n195 0.00134872
R56876 VINP.n105 VINP.n21 0.00134872
R56877 VINP.n510 VINP.n196 0.00134872
R56878 VINP.n104 VINP.n20 0.00134872
R56879 VINP.n511 VINP.n197 0.00134872
R56880 VINP.n103 VINP.n19 0.00134872
R56881 VINP.n512 VINP.n198 0.00134872
R56882 VINP.n102 VINP.n18 0.00134872
R56883 VINP.n513 VINP.n199 0.00134872
R56884 VINP.n101 VINP.n17 0.00134872
R56885 VINP.n514 VINP.n200 0.00134872
R56886 VINP.n100 VINP.n16 0.00134872
R56887 VINP.n515 VINP.n201 0.00134872
R56888 VINP.n99 VINP.n15 0.00134872
R56889 VINP.n516 VINP.n202 0.00134872
R56890 VINP.n98 VINP.n14 0.00134872
R56891 VINP.n517 VINP.n203 0.00134872
R56892 VINP.n97 VINP.n13 0.00134872
R56893 VINP.n518 VINP.n204 0.00134872
R56894 VINP.n96 VINP.n12 0.00134872
R56895 VINP.n519 VINP.n205 0.00134872
R56896 VINP.n95 VINP.n11 0.00134872
R56897 VINP.n520 VINP.n206 0.00134872
R56898 VINP.n94 VINP.n10 0.00134872
R56899 VINP.n521 VINP.n207 0.00134872
R56900 VINP.n93 VINP.n9 0.00134872
R56901 VINP.n522 VINP.n208 0.00134872
R56902 VINP.n92 VINP.n8 0.00134872
R56903 VINP.n523 VINP.n209 0.00134872
R56904 VINP.n91 VINP.n7 0.00134872
R56905 VINP.n524 VINP.n210 0.00134872
R56906 VINP.n90 VINP.n6 0.00134872
R56907 VINP.n525 VINP.n211 0.00134872
R56908 VINP.n89 VINP.n5 0.00134872
R56909 VINP.n526 VINP.n212 0.00134872
R56910 VINP.n88 VINP.n4 0.00134872
R56911 VINP.n527 VINP.n213 0.00134872
R56912 VINP.n87 VINP.n3 0.00134872
R56913 VINP.n655 VINP.n214 0.00134872
R56914 VINP.n86 VINP.n2 0.00134872
R56915 VINP.n66 VINP.n0 0.00134872
R56916 VINP.n656 VINP.n150 0.00134872
R56917 VINP.n528 VINP.n465 0.00134872
R56918 VINP.n654 VINP.n464 0.00134872
R56919 VINP.n399 VINP.n215 0.00134872
R56920 VINP.n401 VINP.n400 0.00134872
R56921 VINP.n397 VINP.n216 0.00134872
R56922 VINP.n402 VINP.n398 0.00134872
R56923 VINP.n395 VINP.n217 0.00134872
R56924 VINP.n403 VINP.n396 0.00134872
R56925 VINP.n393 VINP.n218 0.00134872
R56926 VINP.n404 VINP.n394 0.00134872
R56927 VINP.n391 VINP.n219 0.00134872
R56928 VINP.n405 VINP.n392 0.00134872
R56929 VINP.n389 VINP.n220 0.00134872
R56930 VINP.n406 VINP.n390 0.00134872
R56931 VINP.n387 VINP.n221 0.00134872
R56932 VINP.n407 VINP.n388 0.00134872
R56933 VINP.n385 VINP.n222 0.00134872
R56934 VINP.n408 VINP.n386 0.00134872
R56935 VINP.n383 VINP.n223 0.00134872
R56936 VINP.n409 VINP.n384 0.00134872
R56937 VINP.n381 VINP.n224 0.00134872
R56938 VINP.n410 VINP.n382 0.00134872
R56939 VINP.n379 VINP.n225 0.00134872
R56940 VINP.n411 VINP.n380 0.00134872
R56941 VINP.n377 VINP.n226 0.00134872
R56942 VINP.n412 VINP.n378 0.00134872
R56943 VINP.n375 VINP.n227 0.00134872
R56944 VINP.n413 VINP.n376 0.00134872
R56945 VINP.n373 VINP.n228 0.00134872
R56946 VINP.n414 VINP.n374 0.00134872
R56947 VINP.n371 VINP.n229 0.00134872
R56948 VINP.n415 VINP.n372 0.00134872
R56949 VINP.n369 VINP.n230 0.00134872
R56950 VINP.n416 VINP.n370 0.00134872
R56951 VINP.n367 VINP.n231 0.00134872
R56952 VINP.n417 VINP.n368 0.00134872
R56953 VINP.n365 VINP.n232 0.00134872
R56954 VINP.n418 VINP.n366 0.00134872
R56955 VINP.n363 VINP.n233 0.00134872
R56956 VINP.n419 VINP.n364 0.00134872
R56957 VINP.n361 VINP.n234 0.00134872
R56958 VINP.n420 VINP.n362 0.00134872
R56959 VINP.n359 VINP.n235 0.00134872
R56960 VINP.n421 VINP.n360 0.00134872
R56961 VINP.n357 VINP.n236 0.00134872
R56962 VINP.n422 VINP.n358 0.00134872
R56963 VINP.n355 VINP.n237 0.00134872
R56964 VINP.n423 VINP.n356 0.00134872
R56965 VINP.n353 VINP.n238 0.00134872
R56966 VINP.n424 VINP.n354 0.00134872
R56967 VINP.n351 VINP.n239 0.00134872
R56968 VINP.n425 VINP.n352 0.00134872
R56969 VINP.n349 VINP.n240 0.00134872
R56970 VINP.n426 VINP.n350 0.00134872
R56971 VINP.n347 VINP.n241 0.00134872
R56972 VINP.n427 VINP.n348 0.00134872
R56973 VINP.n345 VINP.n242 0.00134872
R56974 VINP.n428 VINP.n346 0.00134872
R56975 VINP.n343 VINP.n243 0.00134872
R56976 VINP.n429 VINP.n344 0.00134872
R56977 VINP.n341 VINP.n244 0.00134872
R56978 VINP.n430 VINP.n342 0.00134872
R56979 VINP.n339 VINP.n245 0.00134872
R56980 VINP.n431 VINP.n340 0.00134872
R56981 VINP.n337 VINP.n246 0.00134872
R56982 VINP.n432 VINP.n338 0.00134872
R56983 VINP.n335 VINP.n247 0.00134872
R56984 VINP.n433 VINP.n336 0.00134872
R56985 VINP.n333 VINP.n248 0.00134872
R56986 VINP.n434 VINP.n334 0.00134872
R56987 VINP.n331 VINP.n249 0.00134872
R56988 VINP.n435 VINP.n332 0.00134872
R56989 VINP.n329 VINP.n250 0.00134872
R56990 VINP.n436 VINP.n330 0.00134872
R56991 VINP.n327 VINP.n251 0.00134872
R56992 VINP.n437 VINP.n328 0.00134872
R56993 VINP.n325 VINP.n252 0.00134872
R56994 VINP.n438 VINP.n326 0.00134872
R56995 VINP.n323 VINP.n253 0.00134872
R56996 VINP.n439 VINP.n324 0.00134872
R56997 VINP.n321 VINP.n254 0.00134872
R56998 VINP.n440 VINP.n322 0.00134872
R56999 VINP.n319 VINP.n255 0.00134872
R57000 VINP.n441 VINP.n320 0.00134872
R57001 VINP.n317 VINP.n256 0.00134872
R57002 VINP.n442 VINP.n318 0.00134872
R57003 VINP.n315 VINP.n257 0.00134872
R57004 VINP.n443 VINP.n316 0.00134872
R57005 VINP.n313 VINP.n258 0.00134872
R57006 VINP.n444 VINP.n314 0.00134872
R57007 VINP.n311 VINP.n259 0.00134872
R57008 VINP.n445 VINP.n312 0.00134872
R57009 VINP.n309 VINP.n260 0.00134872
R57010 VINP.n446 VINP.n310 0.00134872
R57011 VINP.n307 VINP.n261 0.00134872
R57012 VINP.n447 VINP.n308 0.00134872
R57013 VINP.n305 VINP.n262 0.00134872
R57014 VINP.n448 VINP.n306 0.00134872
R57015 VINP.n303 VINP.n263 0.00134872
R57016 VINP.n449 VINP.n304 0.00134872
R57017 VINP.n301 VINP.n264 0.00134872
R57018 VINP.n450 VINP.n302 0.00134872
R57019 VINP.n299 VINP.n265 0.00134872
R57020 VINP.n451 VINP.n300 0.00134872
R57021 VINP.n297 VINP.n266 0.00134872
R57022 VINP.n452 VINP.n298 0.00134872
R57023 VINP.n295 VINP.n267 0.00134872
R57024 VINP.n453 VINP.n296 0.00134872
R57025 VINP.n293 VINP.n268 0.00134872
R57026 VINP.n454 VINP.n294 0.00134872
R57027 VINP.n291 VINP.n269 0.00134872
R57028 VINP.n455 VINP.n292 0.00134872
R57029 VINP.n289 VINP.n270 0.00134872
R57030 VINP.n456 VINP.n290 0.00134872
R57031 VINP.n287 VINP.n271 0.00134872
R57032 VINP.n457 VINP.n288 0.00134872
R57033 VINP.n285 VINP.n272 0.00134872
R57034 VINP.n458 VINP.n286 0.00134872
R57035 VINP.n283 VINP.n273 0.00134872
R57036 VINP.n459 VINP.n284 0.00134872
R57037 VINP.n281 VINP.n274 0.00134872
R57038 VINP.n460 VINP.n282 0.00134872
R57039 VINP.n279 VINP.n275 0.00134872
R57040 VINP.n461 VINP.n280 0.00134872
R57041 VINP.n277 VINP.n276 0.00134872
R57042 VINP.n461 VINP.n276 0.00134872
R57043 VINP.n460 VINP.n275 0.00134872
R57044 VINP.n459 VINP.n274 0.00134872
R57045 VINP.n458 VINP.n273 0.00134872
R57046 VINP.n457 VINP.n272 0.00134872
R57047 VINP.n456 VINP.n271 0.00134872
R57048 VINP.n455 VINP.n270 0.00134872
R57049 VINP.n454 VINP.n269 0.00134872
R57050 VINP.n453 VINP.n268 0.00134872
R57051 VINP.n452 VINP.n267 0.00134872
R57052 VINP.n451 VINP.n266 0.00134872
R57053 VINP.n450 VINP.n265 0.00134872
R57054 VINP.n449 VINP.n264 0.00134872
R57055 VINP.n448 VINP.n263 0.00134872
R57056 VINP.n447 VINP.n262 0.00134872
R57057 VINP.n446 VINP.n261 0.00134872
R57058 VINP.n445 VINP.n260 0.00134872
R57059 VINP.n444 VINP.n259 0.00134872
R57060 VINP.n443 VINP.n258 0.00134872
R57061 VINP.n442 VINP.n257 0.00134872
R57062 VINP.n441 VINP.n256 0.00134872
R57063 VINP.n440 VINP.n255 0.00134872
R57064 VINP.n439 VINP.n254 0.00134872
R57065 VINP.n438 VINP.n253 0.00134872
R57066 VINP.n437 VINP.n252 0.00134872
R57067 VINP.n436 VINP.n251 0.00134872
R57068 VINP.n435 VINP.n250 0.00134872
R57069 VINP.n434 VINP.n249 0.00134872
R57070 VINP.n433 VINP.n248 0.00134872
R57071 VINP.n432 VINP.n247 0.00134872
R57072 VINP.n431 VINP.n246 0.00134872
R57073 VINP.n430 VINP.n245 0.00134872
R57074 VINP.n429 VINP.n244 0.00134872
R57075 VINP.n428 VINP.n243 0.00134872
R57076 VINP.n427 VINP.n242 0.00134872
R57077 VINP.n426 VINP.n241 0.00134872
R57078 VINP.n425 VINP.n240 0.00134872
R57079 VINP.n424 VINP.n239 0.00134872
R57080 VINP.n423 VINP.n238 0.00134872
R57081 VINP.n422 VINP.n237 0.00134872
R57082 VINP.n421 VINP.n236 0.00134872
R57083 VINP.n420 VINP.n235 0.00134872
R57084 VINP.n419 VINP.n234 0.00134872
R57085 VINP.n418 VINP.n233 0.00134872
R57086 VINP.n417 VINP.n232 0.00134872
R57087 VINP.n416 VINP.n231 0.00134872
R57088 VINP.n415 VINP.n230 0.00134872
R57089 VINP.n414 VINP.n229 0.00134872
R57090 VINP.n413 VINP.n228 0.00134872
R57091 VINP.n412 VINP.n227 0.00134872
R57092 VINP.n411 VINP.n226 0.00134872
R57093 VINP.n410 VINP.n225 0.00134872
R57094 VINP.n409 VINP.n224 0.00134872
R57095 VINP.n408 VINP.n223 0.00134872
R57096 VINP.n407 VINP.n222 0.00134872
R57097 VINP.n406 VINP.n221 0.00134872
R57098 VINP.n405 VINP.n220 0.00134872
R57099 VINP.n404 VINP.n219 0.00134872
R57100 VINP.n403 VINP.n218 0.00134872
R57101 VINP.n402 VINP.n217 0.00134872
R57102 VINP.n401 VINP.n216 0.00134872
R57103 VINP.n464 VINP.n215 0.00134872
R57104 VINP.n528 VINP.n150 0.00134872
R57105 VINP.n657 VINP.n66 0.00134872
R57106 VINP.n462 VINP.n151 0.00134872
R57107 VINP.n280 VINP.n279 0.00134872
R57108 VINP.n282 VINP.n281 0.00134872
R57109 VINP.n284 VINP.n283 0.00134872
R57110 VINP.n286 VINP.n285 0.00134872
R57111 VINP.n288 VINP.n287 0.00134872
R57112 VINP.n290 VINP.n289 0.00134872
R57113 VINP.n292 VINP.n291 0.00134872
R57114 VINP.n294 VINP.n293 0.00134872
R57115 VINP.n296 VINP.n295 0.00134872
R57116 VINP.n298 VINP.n297 0.00134872
R57117 VINP.n300 VINP.n299 0.00134872
R57118 VINP.n302 VINP.n301 0.00134872
R57119 VINP.n304 VINP.n303 0.00134872
R57120 VINP.n306 VINP.n305 0.00134872
R57121 VINP.n308 VINP.n307 0.00134872
R57122 VINP.n310 VINP.n309 0.00134872
R57123 VINP.n312 VINP.n311 0.00134872
R57124 VINP.n314 VINP.n313 0.00134872
R57125 VINP.n316 VINP.n315 0.00134872
R57126 VINP.n318 VINP.n317 0.00134872
R57127 VINP.n320 VINP.n319 0.00134872
R57128 VINP.n322 VINP.n321 0.00134872
R57129 VINP.n324 VINP.n323 0.00134872
R57130 VINP.n326 VINP.n325 0.00134872
R57131 VINP.n328 VINP.n327 0.00134872
R57132 VINP.n330 VINP.n329 0.00134872
R57133 VINP.n332 VINP.n331 0.00134872
R57134 VINP.n334 VINP.n333 0.00134872
R57135 VINP.n336 VINP.n335 0.00134872
R57136 VINP.n338 VINP.n337 0.00134872
R57137 VINP.n340 VINP.n339 0.00134872
R57138 VINP.n342 VINP.n341 0.00134872
R57139 VINP.n344 VINP.n343 0.00134872
R57140 VINP.n346 VINP.n345 0.00134872
R57141 VINP.n348 VINP.n347 0.00134872
R57142 VINP.n350 VINP.n349 0.00134872
R57143 VINP.n352 VINP.n351 0.00134872
R57144 VINP.n354 VINP.n353 0.00134872
R57145 VINP.n356 VINP.n355 0.00134872
R57146 VINP.n358 VINP.n357 0.00134872
R57147 VINP.n360 VINP.n359 0.00134872
R57148 VINP.n362 VINP.n361 0.00134872
R57149 VINP.n364 VINP.n363 0.00134872
R57150 VINP.n366 VINP.n365 0.00134872
R57151 VINP.n368 VINP.n367 0.00134872
R57152 VINP.n370 VINP.n369 0.00134872
R57153 VINP.n372 VINP.n371 0.00134872
R57154 VINP.n374 VINP.n373 0.00134872
R57155 VINP.n376 VINP.n375 0.00134872
R57156 VINP.n378 VINP.n377 0.00134872
R57157 VINP.n380 VINP.n379 0.00134872
R57158 VINP.n382 VINP.n381 0.00134872
R57159 VINP.n384 VINP.n383 0.00134872
R57160 VINP.n386 VINP.n385 0.00134872
R57161 VINP.n388 VINP.n387 0.00134872
R57162 VINP.n390 VINP.n389 0.00134872
R57163 VINP.n392 VINP.n391 0.00134872
R57164 VINP.n394 VINP.n393 0.00134872
R57165 VINP.n396 VINP.n395 0.00134872
R57166 VINP.n398 VINP.n397 0.00134872
R57167 VINP.n400 VINP.n399 0.00134872
R57168 VINP.n654 VINP.n465 0.00134872
R57169 VINP.n151 VINP.n65 0.00134872
R57170 VINP.n278 VINP.n277 0.00134872
R57171 VINP.n466 VINP.n149 0.00134872
R57172 VINP.n152 VINP.n64 0.00134872
R57173 VINP.n467 VINP.n148 0.00134872
R57174 VINP.n153 VINP.n63 0.00134872
R57175 VINP.n468 VINP.n147 0.00134872
R57176 VINP.n154 VINP.n62 0.00134872
R57177 VINP.n469 VINP.n146 0.00134872
R57178 VINP.n155 VINP.n61 0.00134872
R57179 VINP.n470 VINP.n145 0.00134872
R57180 VINP.n156 VINP.n60 0.00134872
R57181 VINP.n471 VINP.n144 0.00134872
R57182 VINP.n157 VINP.n59 0.00134872
R57183 VINP.n472 VINP.n143 0.00134872
R57184 VINP.n158 VINP.n58 0.00134872
R57185 VINP.n473 VINP.n142 0.00134872
R57186 VINP.n159 VINP.n57 0.00134872
R57187 VINP.n474 VINP.n141 0.00134872
R57188 VINP.n160 VINP.n56 0.00134872
R57189 VINP.n475 VINP.n140 0.00134872
R57190 VINP.n161 VINP.n55 0.00134872
R57191 VINP.n476 VINP.n139 0.00134872
R57192 VINP.n162 VINP.n54 0.00134872
R57193 VINP.n477 VINP.n138 0.00134872
R57194 VINP.n163 VINP.n53 0.00134872
R57195 VINP.n478 VINP.n137 0.00134872
R57196 VINP.n164 VINP.n52 0.00134872
R57197 VINP.n479 VINP.n136 0.00134872
R57198 VINP.n165 VINP.n51 0.00134872
R57199 VINP.n480 VINP.n135 0.00134872
R57200 VINP.n166 VINP.n50 0.00134872
R57201 VINP.n481 VINP.n134 0.00134872
R57202 VINP.n167 VINP.n49 0.00134872
R57203 VINP.n482 VINP.n133 0.00134872
R57204 VINP.n168 VINP.n48 0.00134872
R57205 VINP.n483 VINP.n132 0.00134872
R57206 VINP.n169 VINP.n47 0.00134872
R57207 VINP.n484 VINP.n131 0.00134872
R57208 VINP.n170 VINP.n46 0.00134872
R57209 VINP.n485 VINP.n130 0.00134872
R57210 VINP.n171 VINP.n45 0.00134872
R57211 VINP.n486 VINP.n129 0.00134872
R57212 VINP.n172 VINP.n44 0.00134872
R57213 VINP.n487 VINP.n128 0.00134872
R57214 VINP.n173 VINP.n43 0.00134872
R57215 VINP.n488 VINP.n127 0.00134872
R57216 VINP.n174 VINP.n42 0.00134872
R57217 VINP.n489 VINP.n126 0.00134872
R57218 VINP.n175 VINP.n41 0.00134872
R57219 VINP.n490 VINP.n125 0.00134872
R57220 VINP.n176 VINP.n40 0.00134872
R57221 VINP.n491 VINP.n124 0.00134872
R57222 VINP.n177 VINP.n39 0.00134872
R57223 VINP.n492 VINP.n123 0.00134872
R57224 VINP.n178 VINP.n38 0.00134872
R57225 VINP.n493 VINP.n122 0.00134872
R57226 VINP.n179 VINP.n37 0.00134872
R57227 VINP.n494 VINP.n121 0.00134872
R57228 VINP.n180 VINP.n36 0.00134872
R57229 VINP.n495 VINP.n120 0.00134872
R57230 VINP.n181 VINP.n35 0.00134872
R57231 VINP.n496 VINP.n119 0.00134872
R57232 VINP.n182 VINP.n34 0.00134872
R57233 VINP.n497 VINP.n118 0.00134872
R57234 VINP.n183 VINP.n33 0.00134872
R57235 VINP.n498 VINP.n117 0.00134872
R57236 VINP.n184 VINP.n32 0.00134872
R57237 VINP.n499 VINP.n116 0.00134872
R57238 VINP.n185 VINP.n31 0.00134872
R57239 VINP.n500 VINP.n115 0.00134872
R57240 VINP.n186 VINP.n30 0.00134872
R57241 VINP.n501 VINP.n114 0.00134872
R57242 VINP.n187 VINP.n29 0.00134872
R57243 VINP.n502 VINP.n113 0.00134872
R57244 VINP.n188 VINP.n28 0.00134872
R57245 VINP.n503 VINP.n112 0.00134872
R57246 VINP.n189 VINP.n27 0.00134872
R57247 VINP.n504 VINP.n111 0.00134872
R57248 VINP.n190 VINP.n26 0.00134872
R57249 VINP.n505 VINP.n110 0.00134872
R57250 VINP.n191 VINP.n25 0.00134872
R57251 VINP.n506 VINP.n109 0.00134872
R57252 VINP.n192 VINP.n24 0.00134872
R57253 VINP.n507 VINP.n108 0.00134872
R57254 VINP.n193 VINP.n23 0.00134872
R57255 VINP.n508 VINP.n107 0.00134872
R57256 VINP.n194 VINP.n22 0.00134872
R57257 VINP.n509 VINP.n106 0.00134872
R57258 VINP.n195 VINP.n21 0.00134872
R57259 VINP.n510 VINP.n105 0.00134872
R57260 VINP.n196 VINP.n20 0.00134872
R57261 VINP.n511 VINP.n104 0.00134872
R57262 VINP.n197 VINP.n19 0.00134872
R57263 VINP.n512 VINP.n103 0.00134872
R57264 VINP.n198 VINP.n18 0.00134872
R57265 VINP.n513 VINP.n102 0.00134872
R57266 VINP.n199 VINP.n17 0.00134872
R57267 VINP.n514 VINP.n101 0.00134872
R57268 VINP.n200 VINP.n16 0.00134872
R57269 VINP.n515 VINP.n100 0.00134872
R57270 VINP.n201 VINP.n15 0.00134872
R57271 VINP.n516 VINP.n99 0.00134872
R57272 VINP.n202 VINP.n14 0.00134872
R57273 VINP.n517 VINP.n98 0.00134872
R57274 VINP.n203 VINP.n13 0.00134872
R57275 VINP.n518 VINP.n97 0.00134872
R57276 VINP.n204 VINP.n12 0.00134872
R57277 VINP.n519 VINP.n96 0.00134872
R57278 VINP.n205 VINP.n11 0.00134872
R57279 VINP.n520 VINP.n95 0.00134872
R57280 VINP.n206 VINP.n10 0.00134872
R57281 VINP.n521 VINP.n94 0.00134872
R57282 VINP.n207 VINP.n9 0.00134872
R57283 VINP.n522 VINP.n93 0.00134872
R57284 VINP.n208 VINP.n8 0.00134872
R57285 VINP.n523 VINP.n92 0.00134872
R57286 VINP.n209 VINP.n7 0.00134872
R57287 VINP.n524 VINP.n91 0.00134872
R57288 VINP.n210 VINP.n6 0.00134872
R57289 VINP.n525 VINP.n90 0.00134872
R57290 VINP.n211 VINP.n5 0.00134872
R57291 VINP.n526 VINP.n89 0.00134872
R57292 VINP.n212 VINP.n4 0.00134872
R57293 VINP.n527 VINP.n88 0.00134872
R57294 VINP.n213 VINP.n3 0.00134872
R57295 VINP.n214 VINP.n87 0.00134872
R57296 VINP.n655 VINP.n2 0.00134872
R57297 VINP.n657 VINP.n656 0.0011975
R57298 VINP.n658 VINP.n1 0.000965
R57299 VINP.n529 VINP.n1 0.000965
R57300 VINP.n653 VINP.n529 0.000965
R57301 VINP.n653 VINP.n652 0.000965
R57302 VINP.n652 VINP.n651 0.000965
R57303 VINP.n651 VINP.n650 0.000965
R57304 VINP.n650 VINP.n649 0.000965
R57305 VINP.n649 VINP.n648 0.000965
R57306 VINP.n648 VINP.n647 0.000965
R57307 VINP.n647 VINP.n646 0.000965
R57308 VINP.n646 VINP.n645 0.000965
R57309 VINP.n645 VINP.n644 0.000965
R57310 VINP.n644 VINP.n643 0.000965
R57311 VINP.n643 VINP.n642 0.000965
R57312 VINP.n642 VINP.n641 0.000965
R57313 VINP.n641 VINP.n640 0.000965
R57314 VINP.n640 VINP.n639 0.000965
R57315 VINP.n639 VINP.n638 0.000965
R57316 VINP.n638 VINP.n637 0.000965
R57317 VINP.n637 VINP.n636 0.000965
R57318 VINP.n636 VINP.n635 0.000965
R57319 VINP.n635 VINP.n634 0.000965
R57320 VINP.n634 VINP.n633 0.000965
R57321 VINP.n633 VINP.n632 0.000965
R57322 VINP.n632 VINP.n631 0.000965
R57323 VINP.n631 VINP.n630 0.000965
R57324 VINP.n630 VINP.n629 0.000965
R57325 VINP.n629 VINP.n628 0.000965
R57326 VINP.n628 VINP.n627 0.000965
R57327 VINP.n627 VINP.n626 0.000965
R57328 VINP.n626 VINP.n625 0.000965
R57329 VINP.n625 VINP.n624 0.000965
R57330 VINP.n624 VINP.n623 0.000965
R57331 VINP.n623 VINP.n622 0.000965
R57332 VINP.n622 VINP.n621 0.000965
R57333 VINP.n621 VINP.n620 0.000965
R57334 VINP.n620 VINP.n619 0.000965
R57335 VINP.n619 VINP.n618 0.000965
R57336 VINP.n618 VINP.n617 0.000965
R57337 VINP.n617 VINP.n616 0.000965
R57338 VINP.n616 VINP.n615 0.000965
R57339 VINP.n615 VINP.n614 0.000965
R57340 VINP.n614 VINP.n613 0.000965
R57341 VINP.n613 VINP.n612 0.000965
R57342 VINP.n612 VINP.n611 0.000965
R57343 VINP.n611 VINP.n610 0.000965
R57344 VINP.n610 VINP.n609 0.000965
R57345 VINP.n609 VINP.n608 0.000965
R57346 VINP.n608 VINP.n607 0.000965
R57347 VINP.n607 VINP.n606 0.000965
R57348 VINP.n606 VINP.n605 0.000965
R57349 VINP.n605 VINP.n604 0.000965
R57350 VINP.n604 VINP.n603 0.000965
R57351 VINP.n603 VINP.n602 0.000965
R57352 VINP.n602 VINP.n601 0.000965
R57353 VINP.n601 VINP.n600 0.000965
R57354 VINP.n600 VINP.n599 0.000965
R57355 VINP.n599 VINP.n598 0.000965
R57356 VINP.n598 VINP.n597 0.000965
R57357 VINP.n597 VINP.n596 0.000965
R57358 VINP.n596 VINP.n595 0.000965
R57359 VINP.n595 VINP.n594 0.000965
R57360 VINP.n594 VINP.n593 0.000965
R57361 VINP.n593 VINP.n592 0.000965
R57362 VINP.n592 VINP.n591 0.000965
R57363 VINP.n591 VINP.n590 0.000965
R57364 VINP.n590 VINP.n589 0.000965
R57365 VINP.n589 VINP.n588 0.000965
R57366 VINP.n588 VINP.n587 0.000965
R57367 VINP.n587 VINP.n586 0.000965
R57368 VINP.n586 VINP.n585 0.000965
R57369 VINP.n585 VINP.n584 0.000965
R57370 VINP.n584 VINP.n583 0.000965
R57371 VINP.n583 VINP.n582 0.000965
R57372 VINP.n582 VINP.n581 0.000965
R57373 VINP.n581 VINP.n580 0.000965
R57374 VINP.n580 VINP.n579 0.000965
R57375 VINP.n579 VINP.n578 0.000965
R57376 VINP.n578 VINP.n577 0.000965
R57377 VINP.n577 VINP.n576 0.000965
R57378 VINP.n576 VINP.n575 0.000965
R57379 VINP.n574 VINP.n573 0.000965
R57380 VINP.n573 VINP.n572 0.000965
R57381 VINP.n572 VINP.n571 0.000965
R57382 VINP.n571 VINP.n570 0.000965
R57383 VINP.n570 VINP.n569 0.000965
R57384 VINP.n569 VINP.n568 0.000965
R57385 VINP.n568 VINP.n567 0.000965
R57386 VINP.n567 VINP.n566 0.000965
R57387 VINP.n566 VINP.n565 0.000965
R57388 VINP.n565 VINP.n564 0.000965
R57389 VINP.n564 VINP.n563 0.000965
R57390 VINP.n563 VINP.n562 0.000965
R57391 VINP.n562 VINP.n561 0.000965
R57392 VINP.n561 VINP.n560 0.000965
R57393 VINP.n560 VINP.n559 0.000965
R57394 VINP.n559 VINP.n558 0.000965
R57395 VINP.n558 VINP.n557 0.000965
R57396 VINP.n557 VINP.n556 0.000965
R57397 VINP.n556 VINP.n555 0.000965
R57398 VINP.n555 VINP.n554 0.000965
R57399 VINP.n554 VINP.n553 0.000965
R57400 VINP.n553 VINP.n552 0.000965
R57401 VINP.n552 VINP.n551 0.000965
R57402 VINP.n551 VINP.n550 0.000965
R57403 VINP.n550 VINP.n549 0.000965
R57404 VINP.n549 VINP.n548 0.000965
R57405 VINP.n548 VINP.n547 0.000965
R57406 VINP.n547 VINP.n546 0.000965
R57407 VINP.n546 VINP.n545 0.000965
R57408 VINP.n545 VINP.n544 0.000965
R57409 VINP.n544 VINP.n543 0.000965
R57410 VINP.n543 VINP.n542 0.000965
R57411 VINP.n542 VINP.n541 0.000965
R57412 VINP.n541 VINP.n540 0.000965
R57413 VINP.n540 VINP.n539 0.000965
R57414 VINP.n539 VINP.n538 0.000965
R57415 VINP.n538 VINP.n537 0.000965
R57416 VINP.n537 VINP.n536 0.000965
R57417 VINP.n536 VINP.n535 0.000965
R57418 VINP.n535 VINP.n534 0.000965
R57419 VINP.n534 VINP.n533 0.000965
R57420 VINP.n533 VINP.n532 0.000965
R57421 VINP.n532 VINP.n531 0.000965
R57422 VINP.n531 VINP.n530 0.000965
R57423 VINP.n575 VINP 0.00089
R57424 VINP VINP.n574 0.000575
R57425 w_1750_n43456.n33 w_1750_n43456.t78 270.493
R57426 w_1750_n43456.t76 w_1750_n43456.n31 270.493
R57427 w_1750_n43456.t29 w_1750_n43456.n42 270.493
R57428 w_1750_n43456.t13 w_1750_n43456.n43 270.493
R57429 w_1750_n43456.n31 w_1750_n43456.n9 235.089
R57430 w_1750_n43456.n31 w_1750_n43456.n10 235.089
R57431 w_1750_n43456.n33 w_1750_n43456.n10 235.089
R57432 w_1750_n43456.n33 w_1750_n43456.n9 235.089
R57433 w_1750_n43456.n48 w_1750_n43456.n43 235.089
R57434 w_1750_n43456.n46 w_1750_n43456.n43 235.089
R57435 w_1750_n43456.n46 w_1750_n43456.n42 235.089
R57436 w_1750_n43456.n48 w_1750_n43456.n42 235.089
R57437 w_1750_n43456.t78 w_1750_n43456.t54 169.28
R57438 w_1750_n43456.t54 w_1750_n43456.t58 169.28
R57439 w_1750_n43456.t58 w_1750_n43456.t70 169.28
R57440 w_1750_n43456.t70 w_1750_n43456.t80 169.28
R57441 w_1750_n43456.t80 w_1750_n43456.t62 169.28
R57442 w_1750_n43456.t62 w_1750_n43456.t72 169.28
R57443 w_1750_n43456.t72 w_1750_n43456.t46 169.28
R57444 w_1750_n43456.t46 w_1750_n43456.t56 169.28
R57445 w_1750_n43456.t56 w_1750_n43456.t64 169.28
R57446 w_1750_n43456.t48 w_1750_n43456.t44 169.28
R57447 w_1750_n43456.t44 w_1750_n43456.t66 169.28
R57448 w_1750_n43456.t66 w_1750_n43456.t82 169.28
R57449 w_1750_n43456.t82 w_1750_n43456.t50 169.28
R57450 w_1750_n43456.t50 w_1750_n43456.t74 169.28
R57451 w_1750_n43456.t74 w_1750_n43456.t68 169.28
R57452 w_1750_n43456.t68 w_1750_n43456.t52 169.28
R57453 w_1750_n43456.t52 w_1750_n43456.t60 169.28
R57454 w_1750_n43456.t60 w_1750_n43456.t76 169.28
R57455 w_1750_n43456.t3 w_1750_n43456.t29 169.28
R57456 w_1750_n43456.t31 w_1750_n43456.t3 169.28
R57457 w_1750_n43456.t21 w_1750_n43456.t31 169.28
R57458 w_1750_n43456.t11 w_1750_n43456.t21 169.28
R57459 w_1750_n43456.t41 w_1750_n43456.t11 169.28
R57460 w_1750_n43456.t17 w_1750_n43456.t41 169.28
R57461 w_1750_n43456.t5 w_1750_n43456.t17 169.28
R57462 w_1750_n43456.t37 w_1750_n43456.t5 169.28
R57463 w_1750_n43456.t27 w_1750_n43456.t37 169.28
R57464 w_1750_n43456.t15 w_1750_n43456.t33 169.28
R57465 w_1750_n43456.t33 w_1750_n43456.t19 169.28
R57466 w_1750_n43456.t19 w_1750_n43456.t9 169.28
R57467 w_1750_n43456.t9 w_1750_n43456.t35 169.28
R57468 w_1750_n43456.t35 w_1750_n43456.t25 169.28
R57469 w_1750_n43456.t25 w_1750_n43456.t39 169.28
R57470 w_1750_n43456.t39 w_1750_n43456.t7 169.28
R57471 w_1750_n43456.t7 w_1750_n43456.t23 169.28
R57472 w_1750_n43456.t23 w_1750_n43456.t13 169.28
R57473 w_1750_n43456.t64 w_1750_n43456.n32 84.64
R57474 w_1750_n43456.n32 w_1750_n43456.t48 84.64
R57475 w_1750_n43456.n47 w_1750_n43456.t27 84.64
R57476 w_1750_n43456.n47 w_1750_n43456.t15 84.64
R57477 w_1750_n43456.n3 w_1750_n43456.t2 9.53968
R57478 w_1750_n43456.n4 w_1750_n43456.t43 9.32226
R57479 w_1750_n43456.n3 w_1750_n43456.n2 7.97226
R57480 w_1750_n43456.n28 w_1750_n43456.n27 5.72126
R57481 w_1750_n43456.n26 w_1750_n43456.n25 5.72126
R57482 w_1750_n43456.n24 w_1750_n43456.n23 5.72126
R57483 w_1750_n43456.n22 w_1750_n43456.n21 5.72126
R57484 w_1750_n43456.n20 w_1750_n43456.n19 5.72126
R57485 w_1750_n43456.n18 w_1750_n43456.n17 5.72126
R57486 w_1750_n43456.n16 w_1750_n43456.n15 5.72126
R57487 w_1750_n43456.n14 w_1750_n43456.n13 5.72126
R57488 w_1750_n43456.n12 w_1750_n43456.n11 5.72126
R57489 w_1750_n43456.n6 w_1750_n43456.n5 5.72126
R57490 w_1750_n43456.n53 w_1750_n43456.n52 5.72126
R57491 w_1750_n43456.n55 w_1750_n43456.n54 5.72126
R57492 w_1750_n43456.n57 w_1750_n43456.n56 5.72126
R57493 w_1750_n43456.n59 w_1750_n43456.n58 5.72126
R57494 w_1750_n43456.n61 w_1750_n43456.n60 5.72126
R57495 w_1750_n43456.n63 w_1750_n43456.n62 5.72126
R57496 w_1750_n43456.n65 w_1750_n43456.n64 5.72126
R57497 w_1750_n43456.n1 w_1750_n43456.n0 5.72126
R57498 w_1750_n43456.n40 w_1750_n43456.n39 5.72126
R57499 w_1750_n43456.n67 w_1750_n43456.n66 5.72126
R57500 w_1750_n43456.n29 w_1750_n43456.n28 4.62855
R57501 w_1750_n43456.n41 w_1750_n43456.n40 4.62855
R57502 w_1750_n43456.n36 w_1750_n43456.n35 4.50143
R57503 w_1750_n43456.n51 w_1750_n43456.n50 4.50143
R57504 w_1750_n43456.n37 w_1750_n43456.n4 3.4391
R57505 w_1750_n43456.n30 w_1750_n43456.n8 3.35892
R57506 w_1750_n43456.n34 w_1750_n43456.n8 3.35892
R57507 w_1750_n43456.n45 w_1750_n43456.n38 3.35892
R57508 w_1750_n43456.n45 w_1750_n43456.n44 3.35892
R57509 w_1750_n43456.n35 w_1750_n43456.n7 3.05896
R57510 w_1750_n43456.n29 w_1750_n43456.n7 3.05896
R57511 w_1750_n43456.n49 w_1750_n43456.n41 3.05896
R57512 w_1750_n43456.n50 w_1750_n43456.n49 3.0566
R57513 w_1750_n43456.n31 w_1750_n43456.n30 0.9005
R57514 w_1750_n43456.n34 w_1750_n43456.n33 0.9005
R57515 w_1750_n43456.n43 w_1750_n43456.n38 0.9005
R57516 w_1750_n43456.n44 w_1750_n43456.n42 0.9005
R57517 w_1750_n43456.n27 w_1750_n43456.t61 0.6505
R57518 w_1750_n43456.n27 w_1750_n43456.t77 0.6505
R57519 w_1750_n43456.n25 w_1750_n43456.t69 0.6505
R57520 w_1750_n43456.n25 w_1750_n43456.t53 0.6505
R57521 w_1750_n43456.n23 w_1750_n43456.t51 0.6505
R57522 w_1750_n43456.n23 w_1750_n43456.t75 0.6505
R57523 w_1750_n43456.n21 w_1750_n43456.t67 0.6505
R57524 w_1750_n43456.n21 w_1750_n43456.t83 0.6505
R57525 w_1750_n43456.n19 w_1750_n43456.t49 0.6505
R57526 w_1750_n43456.n19 w_1750_n43456.t45 0.6505
R57527 w_1750_n43456.n17 w_1750_n43456.t57 0.6505
R57528 w_1750_n43456.n17 w_1750_n43456.t65 0.6505
R57529 w_1750_n43456.n15 w_1750_n43456.t73 0.6505
R57530 w_1750_n43456.n15 w_1750_n43456.t47 0.6505
R57531 w_1750_n43456.n13 w_1750_n43456.t81 0.6505
R57532 w_1750_n43456.n13 w_1750_n43456.t63 0.6505
R57533 w_1750_n43456.n11 w_1750_n43456.t59 0.6505
R57534 w_1750_n43456.n11 w_1750_n43456.t71 0.6505
R57535 w_1750_n43456.n5 w_1750_n43456.t79 0.6505
R57536 w_1750_n43456.n5 w_1750_n43456.t55 0.6505
R57537 w_1750_n43456.n52 w_1750_n43456.t24 0.6505
R57538 w_1750_n43456.n52 w_1750_n43456.t14 0.6505
R57539 w_1750_n43456.n54 w_1750_n43456.t40 0.6505
R57540 w_1750_n43456.n54 w_1750_n43456.t8 0.6505
R57541 w_1750_n43456.n56 w_1750_n43456.t36 0.6505
R57542 w_1750_n43456.n56 w_1750_n43456.t26 0.6505
R57543 w_1750_n43456.n58 w_1750_n43456.t20 0.6505
R57544 w_1750_n43456.n58 w_1750_n43456.t10 0.6505
R57545 w_1750_n43456.n60 w_1750_n43456.t16 0.6505
R57546 w_1750_n43456.n60 w_1750_n43456.t34 0.6505
R57547 w_1750_n43456.n62 w_1750_n43456.t38 0.6505
R57548 w_1750_n43456.n62 w_1750_n43456.t28 0.6505
R57549 w_1750_n43456.n64 w_1750_n43456.t18 0.6505
R57550 w_1750_n43456.n64 w_1750_n43456.t6 0.6505
R57551 w_1750_n43456.n0 w_1750_n43456.t32 0.6505
R57552 w_1750_n43456.n0 w_1750_n43456.t22 0.6505
R57553 w_1750_n43456.n39 w_1750_n43456.t30 0.6505
R57554 w_1750_n43456.n39 w_1750_n43456.t4 0.6505
R57555 w_1750_n43456.n2 w_1750_n43456.t0 0.6505
R57556 w_1750_n43456.n2 w_1750_n43456.t1 0.6505
R57557 w_1750_n43456.n67 w_1750_n43456.t12 0.6505
R57558 w_1750_n43456.t42 w_1750_n43456.n67 0.6505
R57559 w_1750_n43456.n50 w_1750_n43456.n38 0.302122
R57560 w_1750_n43456.n30 w_1750_n43456.n29 0.299754
R57561 w_1750_n43456.n35 w_1750_n43456.n34 0.299754
R57562 w_1750_n43456.n44 w_1750_n43456.n41 0.299754
R57563 w_1750_n43456.n37 w_1750_n43456.n36 0.22325
R57564 w_1750_n43456.n4 w_1750_n43456.n3 0.217926
R57565 w_1750_n43456.n51 w_1750_n43456.n37 0.206375
R57566 w_1750_n43456.n9 w_1750_n43456.n7 0.13175
R57567 w_1750_n43456.n32 w_1750_n43456.n9 0.13175
R57568 w_1750_n43456.n10 w_1750_n43456.n8 0.13175
R57569 w_1750_n43456.n32 w_1750_n43456.n10 0.13175
R57570 w_1750_n43456.n49 w_1750_n43456.n48 0.13175
R57571 w_1750_n43456.n48 w_1750_n43456.n47 0.13175
R57572 w_1750_n43456.n46 w_1750_n43456.n45 0.13175
R57573 w_1750_n43456.n47 w_1750_n43456.n46 0.13175
R57574 w_1750_n43456.n53 w_1750_n43456.n51 0.127625
R57575 w_1750_n43456.n36 w_1750_n43456.n6 0.127625
R57576 w_1750_n43456.n40 w_1750_n43456.n1 0.122
R57577 w_1750_n43456.n66 w_1750_n43456.n1 0.122
R57578 w_1750_n43456.n66 w_1750_n43456.n65 0.122
R57579 w_1750_n43456.n65 w_1750_n43456.n63 0.122
R57580 w_1750_n43456.n63 w_1750_n43456.n61 0.122
R57581 w_1750_n43456.n61 w_1750_n43456.n59 0.122
R57582 w_1750_n43456.n59 w_1750_n43456.n57 0.122
R57583 w_1750_n43456.n57 w_1750_n43456.n55 0.122
R57584 w_1750_n43456.n55 w_1750_n43456.n53 0.122
R57585 w_1750_n43456.n12 w_1750_n43456.n6 0.122
R57586 w_1750_n43456.n14 w_1750_n43456.n12 0.122
R57587 w_1750_n43456.n16 w_1750_n43456.n14 0.122
R57588 w_1750_n43456.n18 w_1750_n43456.n16 0.122
R57589 w_1750_n43456.n20 w_1750_n43456.n18 0.122
R57590 w_1750_n43456.n22 w_1750_n43456.n20 0.122
R57591 w_1750_n43456.n24 w_1750_n43456.n22 0.122
R57592 w_1750_n43456.n26 w_1750_n43456.n24 0.122
R57593 w_1750_n43456.n28 w_1750_n43456.n26 0.122
R57594 VINN.n67 VINN.t17 41.7362
R57595 VINN.n85 VINN.t16 41.638
R57596 VINN.n84 VINN.t8 41.638
R57597 VINN.n83 VINN.t4 41.638
R57598 VINN.n82 VINN.t12 41.638
R57599 VINN.n81 VINN.t15 41.638
R57600 VINN.n80 VINN.t3 41.638
R57601 VINN.n79 VINN.t19 41.638
R57602 VINN.n78 VINN.t11 41.638
R57603 VINN.n77 VINN.t0 41.638
R57604 VINN.n76 VINN.t2 41.638
R57605 VINN.n75 VINN.t10 41.638
R57606 VINN.n74 VINN.t6 41.638
R57607 VINN.n73 VINN.t1 41.638
R57608 VINN.n72 VINN.t14 41.638
R57609 VINN.n71 VINN.t9 41.638
R57610 VINN.n70 VINN.t18 41.638
R57611 VINN.n69 VINN.t13 41.638
R57612 VINN.n68 VINN.t7 41.638
R57613 VINN.n67 VINN.t5 41.638
R57614 VINN.n86 VINN.n85 10.6308
R57615 VINN.n276 VINN.n151 4.5005
R57616 VINN.n656 VINN.n151 4.5005
R57617 VINN.n151 VINN.n0 4.5005
R57618 VINN.n280 VINN.n149 4.5005
R57619 VINN.n275 VINN.n149 4.5005
R57620 VINN.n282 VINN.n149 4.5005
R57621 VINN.n274 VINN.n149 4.5005
R57622 VINN.n284 VINN.n149 4.5005
R57623 VINN.n273 VINN.n149 4.5005
R57624 VINN.n286 VINN.n149 4.5005
R57625 VINN.n272 VINN.n149 4.5005
R57626 VINN.n288 VINN.n149 4.5005
R57627 VINN.n271 VINN.n149 4.5005
R57628 VINN.n290 VINN.n149 4.5005
R57629 VINN.n270 VINN.n149 4.5005
R57630 VINN.n292 VINN.n149 4.5005
R57631 VINN.n269 VINN.n149 4.5005
R57632 VINN.n294 VINN.n149 4.5005
R57633 VINN.n268 VINN.n149 4.5005
R57634 VINN.n296 VINN.n149 4.5005
R57635 VINN.n267 VINN.n149 4.5005
R57636 VINN.n298 VINN.n149 4.5005
R57637 VINN.n266 VINN.n149 4.5005
R57638 VINN.n300 VINN.n149 4.5005
R57639 VINN.n265 VINN.n149 4.5005
R57640 VINN.n302 VINN.n149 4.5005
R57641 VINN.n264 VINN.n149 4.5005
R57642 VINN.n304 VINN.n149 4.5005
R57643 VINN.n263 VINN.n149 4.5005
R57644 VINN.n306 VINN.n149 4.5005
R57645 VINN.n262 VINN.n149 4.5005
R57646 VINN.n308 VINN.n149 4.5005
R57647 VINN.n261 VINN.n149 4.5005
R57648 VINN.n310 VINN.n149 4.5005
R57649 VINN.n260 VINN.n149 4.5005
R57650 VINN.n312 VINN.n149 4.5005
R57651 VINN.n259 VINN.n149 4.5005
R57652 VINN.n314 VINN.n149 4.5005
R57653 VINN.n258 VINN.n149 4.5005
R57654 VINN.n316 VINN.n149 4.5005
R57655 VINN.n257 VINN.n149 4.5005
R57656 VINN.n318 VINN.n149 4.5005
R57657 VINN.n256 VINN.n149 4.5005
R57658 VINN.n320 VINN.n149 4.5005
R57659 VINN.n255 VINN.n149 4.5005
R57660 VINN.n322 VINN.n149 4.5005
R57661 VINN.n254 VINN.n149 4.5005
R57662 VINN.n324 VINN.n149 4.5005
R57663 VINN.n253 VINN.n149 4.5005
R57664 VINN.n326 VINN.n149 4.5005
R57665 VINN.n252 VINN.n149 4.5005
R57666 VINN.n328 VINN.n149 4.5005
R57667 VINN.n251 VINN.n149 4.5005
R57668 VINN.n330 VINN.n149 4.5005
R57669 VINN.n250 VINN.n149 4.5005
R57670 VINN.n332 VINN.n149 4.5005
R57671 VINN.n249 VINN.n149 4.5005
R57672 VINN.n334 VINN.n149 4.5005
R57673 VINN.n248 VINN.n149 4.5005
R57674 VINN.n336 VINN.n149 4.5005
R57675 VINN.n247 VINN.n149 4.5005
R57676 VINN.n338 VINN.n149 4.5005
R57677 VINN.n246 VINN.n149 4.5005
R57678 VINN.n340 VINN.n149 4.5005
R57679 VINN.n245 VINN.n149 4.5005
R57680 VINN.n342 VINN.n149 4.5005
R57681 VINN.n244 VINN.n149 4.5005
R57682 VINN.n344 VINN.n149 4.5005
R57683 VINN.n243 VINN.n149 4.5005
R57684 VINN.n346 VINN.n149 4.5005
R57685 VINN.n242 VINN.n149 4.5005
R57686 VINN.n348 VINN.n149 4.5005
R57687 VINN.n241 VINN.n149 4.5005
R57688 VINN.n350 VINN.n149 4.5005
R57689 VINN.n240 VINN.n149 4.5005
R57690 VINN.n352 VINN.n149 4.5005
R57691 VINN.n239 VINN.n149 4.5005
R57692 VINN.n354 VINN.n149 4.5005
R57693 VINN.n238 VINN.n149 4.5005
R57694 VINN.n356 VINN.n149 4.5005
R57695 VINN.n237 VINN.n149 4.5005
R57696 VINN.n358 VINN.n149 4.5005
R57697 VINN.n236 VINN.n149 4.5005
R57698 VINN.n360 VINN.n149 4.5005
R57699 VINN.n235 VINN.n149 4.5005
R57700 VINN.n362 VINN.n149 4.5005
R57701 VINN.n234 VINN.n149 4.5005
R57702 VINN.n364 VINN.n149 4.5005
R57703 VINN.n233 VINN.n149 4.5005
R57704 VINN.n366 VINN.n149 4.5005
R57705 VINN.n232 VINN.n149 4.5005
R57706 VINN.n368 VINN.n149 4.5005
R57707 VINN.n231 VINN.n149 4.5005
R57708 VINN.n370 VINN.n149 4.5005
R57709 VINN.n230 VINN.n149 4.5005
R57710 VINN.n372 VINN.n149 4.5005
R57711 VINN.n229 VINN.n149 4.5005
R57712 VINN.n374 VINN.n149 4.5005
R57713 VINN.n228 VINN.n149 4.5005
R57714 VINN.n376 VINN.n149 4.5005
R57715 VINN.n227 VINN.n149 4.5005
R57716 VINN.n378 VINN.n149 4.5005
R57717 VINN.n226 VINN.n149 4.5005
R57718 VINN.n380 VINN.n149 4.5005
R57719 VINN.n225 VINN.n149 4.5005
R57720 VINN.n382 VINN.n149 4.5005
R57721 VINN.n224 VINN.n149 4.5005
R57722 VINN.n384 VINN.n149 4.5005
R57723 VINN.n223 VINN.n149 4.5005
R57724 VINN.n386 VINN.n149 4.5005
R57725 VINN.n222 VINN.n149 4.5005
R57726 VINN.n388 VINN.n149 4.5005
R57727 VINN.n221 VINN.n149 4.5005
R57728 VINN.n390 VINN.n149 4.5005
R57729 VINN.n220 VINN.n149 4.5005
R57730 VINN.n392 VINN.n149 4.5005
R57731 VINN.n219 VINN.n149 4.5005
R57732 VINN.n394 VINN.n149 4.5005
R57733 VINN.n218 VINN.n149 4.5005
R57734 VINN.n396 VINN.n149 4.5005
R57735 VINN.n217 VINN.n149 4.5005
R57736 VINN.n398 VINN.n149 4.5005
R57737 VINN.n216 VINN.n149 4.5005
R57738 VINN.n400 VINN.n149 4.5005
R57739 VINN.n215 VINN.n149 4.5005
R57740 VINN.n654 VINN.n149 4.5005
R57741 VINN.n656 VINN.n149 4.5005
R57742 VINN.n149 VINN.n0 4.5005
R57743 VINN.n278 VINN.n152 4.5005
R57744 VINN.n276 VINN.n152 4.5005
R57745 VINN.n280 VINN.n152 4.5005
R57746 VINN.n275 VINN.n152 4.5005
R57747 VINN.n282 VINN.n152 4.5005
R57748 VINN.n274 VINN.n152 4.5005
R57749 VINN.n284 VINN.n152 4.5005
R57750 VINN.n273 VINN.n152 4.5005
R57751 VINN.n286 VINN.n152 4.5005
R57752 VINN.n272 VINN.n152 4.5005
R57753 VINN.n288 VINN.n152 4.5005
R57754 VINN.n271 VINN.n152 4.5005
R57755 VINN.n290 VINN.n152 4.5005
R57756 VINN.n270 VINN.n152 4.5005
R57757 VINN.n292 VINN.n152 4.5005
R57758 VINN.n269 VINN.n152 4.5005
R57759 VINN.n294 VINN.n152 4.5005
R57760 VINN.n268 VINN.n152 4.5005
R57761 VINN.n296 VINN.n152 4.5005
R57762 VINN.n267 VINN.n152 4.5005
R57763 VINN.n298 VINN.n152 4.5005
R57764 VINN.n266 VINN.n152 4.5005
R57765 VINN.n300 VINN.n152 4.5005
R57766 VINN.n265 VINN.n152 4.5005
R57767 VINN.n302 VINN.n152 4.5005
R57768 VINN.n264 VINN.n152 4.5005
R57769 VINN.n304 VINN.n152 4.5005
R57770 VINN.n263 VINN.n152 4.5005
R57771 VINN.n306 VINN.n152 4.5005
R57772 VINN.n262 VINN.n152 4.5005
R57773 VINN.n308 VINN.n152 4.5005
R57774 VINN.n261 VINN.n152 4.5005
R57775 VINN.n310 VINN.n152 4.5005
R57776 VINN.n260 VINN.n152 4.5005
R57777 VINN.n312 VINN.n152 4.5005
R57778 VINN.n259 VINN.n152 4.5005
R57779 VINN.n314 VINN.n152 4.5005
R57780 VINN.n258 VINN.n152 4.5005
R57781 VINN.n316 VINN.n152 4.5005
R57782 VINN.n257 VINN.n152 4.5005
R57783 VINN.n318 VINN.n152 4.5005
R57784 VINN.n256 VINN.n152 4.5005
R57785 VINN.n320 VINN.n152 4.5005
R57786 VINN.n255 VINN.n152 4.5005
R57787 VINN.n322 VINN.n152 4.5005
R57788 VINN.n254 VINN.n152 4.5005
R57789 VINN.n324 VINN.n152 4.5005
R57790 VINN.n253 VINN.n152 4.5005
R57791 VINN.n326 VINN.n152 4.5005
R57792 VINN.n252 VINN.n152 4.5005
R57793 VINN.n328 VINN.n152 4.5005
R57794 VINN.n251 VINN.n152 4.5005
R57795 VINN.n330 VINN.n152 4.5005
R57796 VINN.n250 VINN.n152 4.5005
R57797 VINN.n332 VINN.n152 4.5005
R57798 VINN.n249 VINN.n152 4.5005
R57799 VINN.n334 VINN.n152 4.5005
R57800 VINN.n248 VINN.n152 4.5005
R57801 VINN.n336 VINN.n152 4.5005
R57802 VINN.n247 VINN.n152 4.5005
R57803 VINN.n338 VINN.n152 4.5005
R57804 VINN.n246 VINN.n152 4.5005
R57805 VINN.n340 VINN.n152 4.5005
R57806 VINN.n245 VINN.n152 4.5005
R57807 VINN.n342 VINN.n152 4.5005
R57808 VINN.n244 VINN.n152 4.5005
R57809 VINN.n344 VINN.n152 4.5005
R57810 VINN.n243 VINN.n152 4.5005
R57811 VINN.n346 VINN.n152 4.5005
R57812 VINN.n242 VINN.n152 4.5005
R57813 VINN.n348 VINN.n152 4.5005
R57814 VINN.n241 VINN.n152 4.5005
R57815 VINN.n350 VINN.n152 4.5005
R57816 VINN.n240 VINN.n152 4.5005
R57817 VINN.n352 VINN.n152 4.5005
R57818 VINN.n239 VINN.n152 4.5005
R57819 VINN.n354 VINN.n152 4.5005
R57820 VINN.n238 VINN.n152 4.5005
R57821 VINN.n356 VINN.n152 4.5005
R57822 VINN.n237 VINN.n152 4.5005
R57823 VINN.n358 VINN.n152 4.5005
R57824 VINN.n236 VINN.n152 4.5005
R57825 VINN.n360 VINN.n152 4.5005
R57826 VINN.n235 VINN.n152 4.5005
R57827 VINN.n362 VINN.n152 4.5005
R57828 VINN.n234 VINN.n152 4.5005
R57829 VINN.n364 VINN.n152 4.5005
R57830 VINN.n233 VINN.n152 4.5005
R57831 VINN.n366 VINN.n152 4.5005
R57832 VINN.n232 VINN.n152 4.5005
R57833 VINN.n368 VINN.n152 4.5005
R57834 VINN.n231 VINN.n152 4.5005
R57835 VINN.n370 VINN.n152 4.5005
R57836 VINN.n230 VINN.n152 4.5005
R57837 VINN.n372 VINN.n152 4.5005
R57838 VINN.n229 VINN.n152 4.5005
R57839 VINN.n374 VINN.n152 4.5005
R57840 VINN.n228 VINN.n152 4.5005
R57841 VINN.n376 VINN.n152 4.5005
R57842 VINN.n227 VINN.n152 4.5005
R57843 VINN.n378 VINN.n152 4.5005
R57844 VINN.n226 VINN.n152 4.5005
R57845 VINN.n380 VINN.n152 4.5005
R57846 VINN.n225 VINN.n152 4.5005
R57847 VINN.n382 VINN.n152 4.5005
R57848 VINN.n224 VINN.n152 4.5005
R57849 VINN.n384 VINN.n152 4.5005
R57850 VINN.n223 VINN.n152 4.5005
R57851 VINN.n386 VINN.n152 4.5005
R57852 VINN.n222 VINN.n152 4.5005
R57853 VINN.n388 VINN.n152 4.5005
R57854 VINN.n221 VINN.n152 4.5005
R57855 VINN.n390 VINN.n152 4.5005
R57856 VINN.n220 VINN.n152 4.5005
R57857 VINN.n392 VINN.n152 4.5005
R57858 VINN.n219 VINN.n152 4.5005
R57859 VINN.n394 VINN.n152 4.5005
R57860 VINN.n218 VINN.n152 4.5005
R57861 VINN.n396 VINN.n152 4.5005
R57862 VINN.n217 VINN.n152 4.5005
R57863 VINN.n398 VINN.n152 4.5005
R57864 VINN.n216 VINN.n152 4.5005
R57865 VINN.n400 VINN.n152 4.5005
R57866 VINN.n215 VINN.n152 4.5005
R57867 VINN.n654 VINN.n152 4.5005
R57868 VINN.n656 VINN.n152 4.5005
R57869 VINN.n152 VINN.n0 4.5005
R57870 VINN.n278 VINN.n148 4.5005
R57871 VINN.n276 VINN.n148 4.5005
R57872 VINN.n280 VINN.n148 4.5005
R57873 VINN.n275 VINN.n148 4.5005
R57874 VINN.n282 VINN.n148 4.5005
R57875 VINN.n274 VINN.n148 4.5005
R57876 VINN.n284 VINN.n148 4.5005
R57877 VINN.n273 VINN.n148 4.5005
R57878 VINN.n286 VINN.n148 4.5005
R57879 VINN.n272 VINN.n148 4.5005
R57880 VINN.n288 VINN.n148 4.5005
R57881 VINN.n271 VINN.n148 4.5005
R57882 VINN.n290 VINN.n148 4.5005
R57883 VINN.n270 VINN.n148 4.5005
R57884 VINN.n292 VINN.n148 4.5005
R57885 VINN.n269 VINN.n148 4.5005
R57886 VINN.n294 VINN.n148 4.5005
R57887 VINN.n268 VINN.n148 4.5005
R57888 VINN.n296 VINN.n148 4.5005
R57889 VINN.n267 VINN.n148 4.5005
R57890 VINN.n298 VINN.n148 4.5005
R57891 VINN.n266 VINN.n148 4.5005
R57892 VINN.n300 VINN.n148 4.5005
R57893 VINN.n265 VINN.n148 4.5005
R57894 VINN.n302 VINN.n148 4.5005
R57895 VINN.n264 VINN.n148 4.5005
R57896 VINN.n304 VINN.n148 4.5005
R57897 VINN.n263 VINN.n148 4.5005
R57898 VINN.n306 VINN.n148 4.5005
R57899 VINN.n262 VINN.n148 4.5005
R57900 VINN.n308 VINN.n148 4.5005
R57901 VINN.n261 VINN.n148 4.5005
R57902 VINN.n310 VINN.n148 4.5005
R57903 VINN.n260 VINN.n148 4.5005
R57904 VINN.n312 VINN.n148 4.5005
R57905 VINN.n259 VINN.n148 4.5005
R57906 VINN.n314 VINN.n148 4.5005
R57907 VINN.n258 VINN.n148 4.5005
R57908 VINN.n316 VINN.n148 4.5005
R57909 VINN.n257 VINN.n148 4.5005
R57910 VINN.n318 VINN.n148 4.5005
R57911 VINN.n256 VINN.n148 4.5005
R57912 VINN.n320 VINN.n148 4.5005
R57913 VINN.n255 VINN.n148 4.5005
R57914 VINN.n322 VINN.n148 4.5005
R57915 VINN.n254 VINN.n148 4.5005
R57916 VINN.n324 VINN.n148 4.5005
R57917 VINN.n253 VINN.n148 4.5005
R57918 VINN.n326 VINN.n148 4.5005
R57919 VINN.n252 VINN.n148 4.5005
R57920 VINN.n328 VINN.n148 4.5005
R57921 VINN.n251 VINN.n148 4.5005
R57922 VINN.n330 VINN.n148 4.5005
R57923 VINN.n250 VINN.n148 4.5005
R57924 VINN.n332 VINN.n148 4.5005
R57925 VINN.n249 VINN.n148 4.5005
R57926 VINN.n334 VINN.n148 4.5005
R57927 VINN.n248 VINN.n148 4.5005
R57928 VINN.n336 VINN.n148 4.5005
R57929 VINN.n247 VINN.n148 4.5005
R57930 VINN.n338 VINN.n148 4.5005
R57931 VINN.n246 VINN.n148 4.5005
R57932 VINN.n340 VINN.n148 4.5005
R57933 VINN.n245 VINN.n148 4.5005
R57934 VINN.n342 VINN.n148 4.5005
R57935 VINN.n244 VINN.n148 4.5005
R57936 VINN.n344 VINN.n148 4.5005
R57937 VINN.n243 VINN.n148 4.5005
R57938 VINN.n346 VINN.n148 4.5005
R57939 VINN.n242 VINN.n148 4.5005
R57940 VINN.n348 VINN.n148 4.5005
R57941 VINN.n241 VINN.n148 4.5005
R57942 VINN.n350 VINN.n148 4.5005
R57943 VINN.n240 VINN.n148 4.5005
R57944 VINN.n352 VINN.n148 4.5005
R57945 VINN.n239 VINN.n148 4.5005
R57946 VINN.n354 VINN.n148 4.5005
R57947 VINN.n238 VINN.n148 4.5005
R57948 VINN.n356 VINN.n148 4.5005
R57949 VINN.n237 VINN.n148 4.5005
R57950 VINN.n358 VINN.n148 4.5005
R57951 VINN.n236 VINN.n148 4.5005
R57952 VINN.n360 VINN.n148 4.5005
R57953 VINN.n235 VINN.n148 4.5005
R57954 VINN.n362 VINN.n148 4.5005
R57955 VINN.n234 VINN.n148 4.5005
R57956 VINN.n364 VINN.n148 4.5005
R57957 VINN.n233 VINN.n148 4.5005
R57958 VINN.n366 VINN.n148 4.5005
R57959 VINN.n232 VINN.n148 4.5005
R57960 VINN.n368 VINN.n148 4.5005
R57961 VINN.n231 VINN.n148 4.5005
R57962 VINN.n370 VINN.n148 4.5005
R57963 VINN.n230 VINN.n148 4.5005
R57964 VINN.n372 VINN.n148 4.5005
R57965 VINN.n229 VINN.n148 4.5005
R57966 VINN.n374 VINN.n148 4.5005
R57967 VINN.n228 VINN.n148 4.5005
R57968 VINN.n376 VINN.n148 4.5005
R57969 VINN.n227 VINN.n148 4.5005
R57970 VINN.n378 VINN.n148 4.5005
R57971 VINN.n226 VINN.n148 4.5005
R57972 VINN.n380 VINN.n148 4.5005
R57973 VINN.n225 VINN.n148 4.5005
R57974 VINN.n382 VINN.n148 4.5005
R57975 VINN.n224 VINN.n148 4.5005
R57976 VINN.n384 VINN.n148 4.5005
R57977 VINN.n223 VINN.n148 4.5005
R57978 VINN.n386 VINN.n148 4.5005
R57979 VINN.n222 VINN.n148 4.5005
R57980 VINN.n388 VINN.n148 4.5005
R57981 VINN.n221 VINN.n148 4.5005
R57982 VINN.n390 VINN.n148 4.5005
R57983 VINN.n220 VINN.n148 4.5005
R57984 VINN.n392 VINN.n148 4.5005
R57985 VINN.n219 VINN.n148 4.5005
R57986 VINN.n394 VINN.n148 4.5005
R57987 VINN.n218 VINN.n148 4.5005
R57988 VINN.n396 VINN.n148 4.5005
R57989 VINN.n217 VINN.n148 4.5005
R57990 VINN.n398 VINN.n148 4.5005
R57991 VINN.n216 VINN.n148 4.5005
R57992 VINN.n400 VINN.n148 4.5005
R57993 VINN.n215 VINN.n148 4.5005
R57994 VINN.n654 VINN.n148 4.5005
R57995 VINN.n656 VINN.n148 4.5005
R57996 VINN.n148 VINN.n0 4.5005
R57997 VINN.n278 VINN.n153 4.5005
R57998 VINN.n276 VINN.n153 4.5005
R57999 VINN.n280 VINN.n153 4.5005
R58000 VINN.n275 VINN.n153 4.5005
R58001 VINN.n282 VINN.n153 4.5005
R58002 VINN.n274 VINN.n153 4.5005
R58003 VINN.n284 VINN.n153 4.5005
R58004 VINN.n273 VINN.n153 4.5005
R58005 VINN.n286 VINN.n153 4.5005
R58006 VINN.n272 VINN.n153 4.5005
R58007 VINN.n288 VINN.n153 4.5005
R58008 VINN.n271 VINN.n153 4.5005
R58009 VINN.n290 VINN.n153 4.5005
R58010 VINN.n270 VINN.n153 4.5005
R58011 VINN.n292 VINN.n153 4.5005
R58012 VINN.n269 VINN.n153 4.5005
R58013 VINN.n294 VINN.n153 4.5005
R58014 VINN.n268 VINN.n153 4.5005
R58015 VINN.n296 VINN.n153 4.5005
R58016 VINN.n267 VINN.n153 4.5005
R58017 VINN.n298 VINN.n153 4.5005
R58018 VINN.n266 VINN.n153 4.5005
R58019 VINN.n300 VINN.n153 4.5005
R58020 VINN.n265 VINN.n153 4.5005
R58021 VINN.n302 VINN.n153 4.5005
R58022 VINN.n264 VINN.n153 4.5005
R58023 VINN.n304 VINN.n153 4.5005
R58024 VINN.n263 VINN.n153 4.5005
R58025 VINN.n306 VINN.n153 4.5005
R58026 VINN.n262 VINN.n153 4.5005
R58027 VINN.n308 VINN.n153 4.5005
R58028 VINN.n261 VINN.n153 4.5005
R58029 VINN.n310 VINN.n153 4.5005
R58030 VINN.n260 VINN.n153 4.5005
R58031 VINN.n312 VINN.n153 4.5005
R58032 VINN.n259 VINN.n153 4.5005
R58033 VINN.n314 VINN.n153 4.5005
R58034 VINN.n258 VINN.n153 4.5005
R58035 VINN.n316 VINN.n153 4.5005
R58036 VINN.n257 VINN.n153 4.5005
R58037 VINN.n318 VINN.n153 4.5005
R58038 VINN.n256 VINN.n153 4.5005
R58039 VINN.n320 VINN.n153 4.5005
R58040 VINN.n255 VINN.n153 4.5005
R58041 VINN.n322 VINN.n153 4.5005
R58042 VINN.n254 VINN.n153 4.5005
R58043 VINN.n324 VINN.n153 4.5005
R58044 VINN.n253 VINN.n153 4.5005
R58045 VINN.n326 VINN.n153 4.5005
R58046 VINN.n252 VINN.n153 4.5005
R58047 VINN.n328 VINN.n153 4.5005
R58048 VINN.n251 VINN.n153 4.5005
R58049 VINN.n330 VINN.n153 4.5005
R58050 VINN.n250 VINN.n153 4.5005
R58051 VINN.n332 VINN.n153 4.5005
R58052 VINN.n249 VINN.n153 4.5005
R58053 VINN.n334 VINN.n153 4.5005
R58054 VINN.n248 VINN.n153 4.5005
R58055 VINN.n336 VINN.n153 4.5005
R58056 VINN.n247 VINN.n153 4.5005
R58057 VINN.n338 VINN.n153 4.5005
R58058 VINN.n246 VINN.n153 4.5005
R58059 VINN.n340 VINN.n153 4.5005
R58060 VINN.n245 VINN.n153 4.5005
R58061 VINN.n342 VINN.n153 4.5005
R58062 VINN.n244 VINN.n153 4.5005
R58063 VINN.n344 VINN.n153 4.5005
R58064 VINN.n243 VINN.n153 4.5005
R58065 VINN.n346 VINN.n153 4.5005
R58066 VINN.n242 VINN.n153 4.5005
R58067 VINN.n348 VINN.n153 4.5005
R58068 VINN.n241 VINN.n153 4.5005
R58069 VINN.n350 VINN.n153 4.5005
R58070 VINN.n240 VINN.n153 4.5005
R58071 VINN.n352 VINN.n153 4.5005
R58072 VINN.n239 VINN.n153 4.5005
R58073 VINN.n354 VINN.n153 4.5005
R58074 VINN.n238 VINN.n153 4.5005
R58075 VINN.n356 VINN.n153 4.5005
R58076 VINN.n237 VINN.n153 4.5005
R58077 VINN.n358 VINN.n153 4.5005
R58078 VINN.n236 VINN.n153 4.5005
R58079 VINN.n360 VINN.n153 4.5005
R58080 VINN.n235 VINN.n153 4.5005
R58081 VINN.n362 VINN.n153 4.5005
R58082 VINN.n234 VINN.n153 4.5005
R58083 VINN.n364 VINN.n153 4.5005
R58084 VINN.n233 VINN.n153 4.5005
R58085 VINN.n366 VINN.n153 4.5005
R58086 VINN.n232 VINN.n153 4.5005
R58087 VINN.n368 VINN.n153 4.5005
R58088 VINN.n231 VINN.n153 4.5005
R58089 VINN.n370 VINN.n153 4.5005
R58090 VINN.n230 VINN.n153 4.5005
R58091 VINN.n372 VINN.n153 4.5005
R58092 VINN.n229 VINN.n153 4.5005
R58093 VINN.n374 VINN.n153 4.5005
R58094 VINN.n228 VINN.n153 4.5005
R58095 VINN.n376 VINN.n153 4.5005
R58096 VINN.n227 VINN.n153 4.5005
R58097 VINN.n378 VINN.n153 4.5005
R58098 VINN.n226 VINN.n153 4.5005
R58099 VINN.n380 VINN.n153 4.5005
R58100 VINN.n225 VINN.n153 4.5005
R58101 VINN.n382 VINN.n153 4.5005
R58102 VINN.n224 VINN.n153 4.5005
R58103 VINN.n384 VINN.n153 4.5005
R58104 VINN.n223 VINN.n153 4.5005
R58105 VINN.n386 VINN.n153 4.5005
R58106 VINN.n222 VINN.n153 4.5005
R58107 VINN.n388 VINN.n153 4.5005
R58108 VINN.n221 VINN.n153 4.5005
R58109 VINN.n390 VINN.n153 4.5005
R58110 VINN.n220 VINN.n153 4.5005
R58111 VINN.n392 VINN.n153 4.5005
R58112 VINN.n219 VINN.n153 4.5005
R58113 VINN.n394 VINN.n153 4.5005
R58114 VINN.n218 VINN.n153 4.5005
R58115 VINN.n396 VINN.n153 4.5005
R58116 VINN.n217 VINN.n153 4.5005
R58117 VINN.n398 VINN.n153 4.5005
R58118 VINN.n216 VINN.n153 4.5005
R58119 VINN.n400 VINN.n153 4.5005
R58120 VINN.n215 VINN.n153 4.5005
R58121 VINN.n654 VINN.n153 4.5005
R58122 VINN.n656 VINN.n153 4.5005
R58123 VINN.n153 VINN.n0 4.5005
R58124 VINN.n278 VINN.n147 4.5005
R58125 VINN.n276 VINN.n147 4.5005
R58126 VINN.n280 VINN.n147 4.5005
R58127 VINN.n275 VINN.n147 4.5005
R58128 VINN.n282 VINN.n147 4.5005
R58129 VINN.n274 VINN.n147 4.5005
R58130 VINN.n284 VINN.n147 4.5005
R58131 VINN.n273 VINN.n147 4.5005
R58132 VINN.n286 VINN.n147 4.5005
R58133 VINN.n272 VINN.n147 4.5005
R58134 VINN.n288 VINN.n147 4.5005
R58135 VINN.n271 VINN.n147 4.5005
R58136 VINN.n290 VINN.n147 4.5005
R58137 VINN.n270 VINN.n147 4.5005
R58138 VINN.n292 VINN.n147 4.5005
R58139 VINN.n269 VINN.n147 4.5005
R58140 VINN.n294 VINN.n147 4.5005
R58141 VINN.n268 VINN.n147 4.5005
R58142 VINN.n296 VINN.n147 4.5005
R58143 VINN.n267 VINN.n147 4.5005
R58144 VINN.n298 VINN.n147 4.5005
R58145 VINN.n266 VINN.n147 4.5005
R58146 VINN.n300 VINN.n147 4.5005
R58147 VINN.n265 VINN.n147 4.5005
R58148 VINN.n302 VINN.n147 4.5005
R58149 VINN.n264 VINN.n147 4.5005
R58150 VINN.n304 VINN.n147 4.5005
R58151 VINN.n263 VINN.n147 4.5005
R58152 VINN.n306 VINN.n147 4.5005
R58153 VINN.n262 VINN.n147 4.5005
R58154 VINN.n308 VINN.n147 4.5005
R58155 VINN.n261 VINN.n147 4.5005
R58156 VINN.n310 VINN.n147 4.5005
R58157 VINN.n260 VINN.n147 4.5005
R58158 VINN.n312 VINN.n147 4.5005
R58159 VINN.n259 VINN.n147 4.5005
R58160 VINN.n314 VINN.n147 4.5005
R58161 VINN.n258 VINN.n147 4.5005
R58162 VINN.n316 VINN.n147 4.5005
R58163 VINN.n257 VINN.n147 4.5005
R58164 VINN.n318 VINN.n147 4.5005
R58165 VINN.n256 VINN.n147 4.5005
R58166 VINN.n320 VINN.n147 4.5005
R58167 VINN.n255 VINN.n147 4.5005
R58168 VINN.n322 VINN.n147 4.5005
R58169 VINN.n254 VINN.n147 4.5005
R58170 VINN.n324 VINN.n147 4.5005
R58171 VINN.n253 VINN.n147 4.5005
R58172 VINN.n326 VINN.n147 4.5005
R58173 VINN.n252 VINN.n147 4.5005
R58174 VINN.n328 VINN.n147 4.5005
R58175 VINN.n251 VINN.n147 4.5005
R58176 VINN.n330 VINN.n147 4.5005
R58177 VINN.n250 VINN.n147 4.5005
R58178 VINN.n332 VINN.n147 4.5005
R58179 VINN.n249 VINN.n147 4.5005
R58180 VINN.n334 VINN.n147 4.5005
R58181 VINN.n248 VINN.n147 4.5005
R58182 VINN.n336 VINN.n147 4.5005
R58183 VINN.n247 VINN.n147 4.5005
R58184 VINN.n338 VINN.n147 4.5005
R58185 VINN.n246 VINN.n147 4.5005
R58186 VINN.n340 VINN.n147 4.5005
R58187 VINN.n245 VINN.n147 4.5005
R58188 VINN.n342 VINN.n147 4.5005
R58189 VINN.n244 VINN.n147 4.5005
R58190 VINN.n344 VINN.n147 4.5005
R58191 VINN.n243 VINN.n147 4.5005
R58192 VINN.n346 VINN.n147 4.5005
R58193 VINN.n242 VINN.n147 4.5005
R58194 VINN.n348 VINN.n147 4.5005
R58195 VINN.n241 VINN.n147 4.5005
R58196 VINN.n350 VINN.n147 4.5005
R58197 VINN.n240 VINN.n147 4.5005
R58198 VINN.n352 VINN.n147 4.5005
R58199 VINN.n239 VINN.n147 4.5005
R58200 VINN.n354 VINN.n147 4.5005
R58201 VINN.n238 VINN.n147 4.5005
R58202 VINN.n356 VINN.n147 4.5005
R58203 VINN.n237 VINN.n147 4.5005
R58204 VINN.n358 VINN.n147 4.5005
R58205 VINN.n236 VINN.n147 4.5005
R58206 VINN.n360 VINN.n147 4.5005
R58207 VINN.n235 VINN.n147 4.5005
R58208 VINN.n362 VINN.n147 4.5005
R58209 VINN.n234 VINN.n147 4.5005
R58210 VINN.n364 VINN.n147 4.5005
R58211 VINN.n233 VINN.n147 4.5005
R58212 VINN.n366 VINN.n147 4.5005
R58213 VINN.n232 VINN.n147 4.5005
R58214 VINN.n368 VINN.n147 4.5005
R58215 VINN.n231 VINN.n147 4.5005
R58216 VINN.n370 VINN.n147 4.5005
R58217 VINN.n230 VINN.n147 4.5005
R58218 VINN.n372 VINN.n147 4.5005
R58219 VINN.n229 VINN.n147 4.5005
R58220 VINN.n374 VINN.n147 4.5005
R58221 VINN.n228 VINN.n147 4.5005
R58222 VINN.n376 VINN.n147 4.5005
R58223 VINN.n227 VINN.n147 4.5005
R58224 VINN.n378 VINN.n147 4.5005
R58225 VINN.n226 VINN.n147 4.5005
R58226 VINN.n380 VINN.n147 4.5005
R58227 VINN.n225 VINN.n147 4.5005
R58228 VINN.n382 VINN.n147 4.5005
R58229 VINN.n224 VINN.n147 4.5005
R58230 VINN.n384 VINN.n147 4.5005
R58231 VINN.n223 VINN.n147 4.5005
R58232 VINN.n386 VINN.n147 4.5005
R58233 VINN.n222 VINN.n147 4.5005
R58234 VINN.n388 VINN.n147 4.5005
R58235 VINN.n221 VINN.n147 4.5005
R58236 VINN.n390 VINN.n147 4.5005
R58237 VINN.n220 VINN.n147 4.5005
R58238 VINN.n392 VINN.n147 4.5005
R58239 VINN.n219 VINN.n147 4.5005
R58240 VINN.n394 VINN.n147 4.5005
R58241 VINN.n218 VINN.n147 4.5005
R58242 VINN.n396 VINN.n147 4.5005
R58243 VINN.n217 VINN.n147 4.5005
R58244 VINN.n398 VINN.n147 4.5005
R58245 VINN.n216 VINN.n147 4.5005
R58246 VINN.n400 VINN.n147 4.5005
R58247 VINN.n215 VINN.n147 4.5005
R58248 VINN.n654 VINN.n147 4.5005
R58249 VINN.n656 VINN.n147 4.5005
R58250 VINN.n147 VINN.n0 4.5005
R58251 VINN.n278 VINN.n154 4.5005
R58252 VINN.n276 VINN.n154 4.5005
R58253 VINN.n280 VINN.n154 4.5005
R58254 VINN.n275 VINN.n154 4.5005
R58255 VINN.n282 VINN.n154 4.5005
R58256 VINN.n274 VINN.n154 4.5005
R58257 VINN.n284 VINN.n154 4.5005
R58258 VINN.n273 VINN.n154 4.5005
R58259 VINN.n286 VINN.n154 4.5005
R58260 VINN.n272 VINN.n154 4.5005
R58261 VINN.n288 VINN.n154 4.5005
R58262 VINN.n271 VINN.n154 4.5005
R58263 VINN.n290 VINN.n154 4.5005
R58264 VINN.n270 VINN.n154 4.5005
R58265 VINN.n292 VINN.n154 4.5005
R58266 VINN.n269 VINN.n154 4.5005
R58267 VINN.n294 VINN.n154 4.5005
R58268 VINN.n268 VINN.n154 4.5005
R58269 VINN.n296 VINN.n154 4.5005
R58270 VINN.n267 VINN.n154 4.5005
R58271 VINN.n298 VINN.n154 4.5005
R58272 VINN.n266 VINN.n154 4.5005
R58273 VINN.n300 VINN.n154 4.5005
R58274 VINN.n265 VINN.n154 4.5005
R58275 VINN.n302 VINN.n154 4.5005
R58276 VINN.n264 VINN.n154 4.5005
R58277 VINN.n304 VINN.n154 4.5005
R58278 VINN.n263 VINN.n154 4.5005
R58279 VINN.n306 VINN.n154 4.5005
R58280 VINN.n262 VINN.n154 4.5005
R58281 VINN.n308 VINN.n154 4.5005
R58282 VINN.n261 VINN.n154 4.5005
R58283 VINN.n310 VINN.n154 4.5005
R58284 VINN.n260 VINN.n154 4.5005
R58285 VINN.n312 VINN.n154 4.5005
R58286 VINN.n259 VINN.n154 4.5005
R58287 VINN.n314 VINN.n154 4.5005
R58288 VINN.n258 VINN.n154 4.5005
R58289 VINN.n316 VINN.n154 4.5005
R58290 VINN.n257 VINN.n154 4.5005
R58291 VINN.n318 VINN.n154 4.5005
R58292 VINN.n256 VINN.n154 4.5005
R58293 VINN.n320 VINN.n154 4.5005
R58294 VINN.n255 VINN.n154 4.5005
R58295 VINN.n322 VINN.n154 4.5005
R58296 VINN.n254 VINN.n154 4.5005
R58297 VINN.n324 VINN.n154 4.5005
R58298 VINN.n253 VINN.n154 4.5005
R58299 VINN.n326 VINN.n154 4.5005
R58300 VINN.n252 VINN.n154 4.5005
R58301 VINN.n328 VINN.n154 4.5005
R58302 VINN.n251 VINN.n154 4.5005
R58303 VINN.n330 VINN.n154 4.5005
R58304 VINN.n250 VINN.n154 4.5005
R58305 VINN.n332 VINN.n154 4.5005
R58306 VINN.n249 VINN.n154 4.5005
R58307 VINN.n334 VINN.n154 4.5005
R58308 VINN.n248 VINN.n154 4.5005
R58309 VINN.n336 VINN.n154 4.5005
R58310 VINN.n247 VINN.n154 4.5005
R58311 VINN.n338 VINN.n154 4.5005
R58312 VINN.n246 VINN.n154 4.5005
R58313 VINN.n340 VINN.n154 4.5005
R58314 VINN.n245 VINN.n154 4.5005
R58315 VINN.n342 VINN.n154 4.5005
R58316 VINN.n244 VINN.n154 4.5005
R58317 VINN.n344 VINN.n154 4.5005
R58318 VINN.n243 VINN.n154 4.5005
R58319 VINN.n346 VINN.n154 4.5005
R58320 VINN.n242 VINN.n154 4.5005
R58321 VINN.n348 VINN.n154 4.5005
R58322 VINN.n241 VINN.n154 4.5005
R58323 VINN.n350 VINN.n154 4.5005
R58324 VINN.n240 VINN.n154 4.5005
R58325 VINN.n352 VINN.n154 4.5005
R58326 VINN.n239 VINN.n154 4.5005
R58327 VINN.n354 VINN.n154 4.5005
R58328 VINN.n238 VINN.n154 4.5005
R58329 VINN.n356 VINN.n154 4.5005
R58330 VINN.n237 VINN.n154 4.5005
R58331 VINN.n358 VINN.n154 4.5005
R58332 VINN.n236 VINN.n154 4.5005
R58333 VINN.n360 VINN.n154 4.5005
R58334 VINN.n235 VINN.n154 4.5005
R58335 VINN.n362 VINN.n154 4.5005
R58336 VINN.n234 VINN.n154 4.5005
R58337 VINN.n364 VINN.n154 4.5005
R58338 VINN.n233 VINN.n154 4.5005
R58339 VINN.n366 VINN.n154 4.5005
R58340 VINN.n232 VINN.n154 4.5005
R58341 VINN.n368 VINN.n154 4.5005
R58342 VINN.n231 VINN.n154 4.5005
R58343 VINN.n370 VINN.n154 4.5005
R58344 VINN.n230 VINN.n154 4.5005
R58345 VINN.n372 VINN.n154 4.5005
R58346 VINN.n229 VINN.n154 4.5005
R58347 VINN.n374 VINN.n154 4.5005
R58348 VINN.n228 VINN.n154 4.5005
R58349 VINN.n376 VINN.n154 4.5005
R58350 VINN.n227 VINN.n154 4.5005
R58351 VINN.n378 VINN.n154 4.5005
R58352 VINN.n226 VINN.n154 4.5005
R58353 VINN.n380 VINN.n154 4.5005
R58354 VINN.n225 VINN.n154 4.5005
R58355 VINN.n382 VINN.n154 4.5005
R58356 VINN.n224 VINN.n154 4.5005
R58357 VINN.n384 VINN.n154 4.5005
R58358 VINN.n223 VINN.n154 4.5005
R58359 VINN.n386 VINN.n154 4.5005
R58360 VINN.n222 VINN.n154 4.5005
R58361 VINN.n388 VINN.n154 4.5005
R58362 VINN.n221 VINN.n154 4.5005
R58363 VINN.n390 VINN.n154 4.5005
R58364 VINN.n220 VINN.n154 4.5005
R58365 VINN.n392 VINN.n154 4.5005
R58366 VINN.n219 VINN.n154 4.5005
R58367 VINN.n394 VINN.n154 4.5005
R58368 VINN.n218 VINN.n154 4.5005
R58369 VINN.n396 VINN.n154 4.5005
R58370 VINN.n217 VINN.n154 4.5005
R58371 VINN.n398 VINN.n154 4.5005
R58372 VINN.n216 VINN.n154 4.5005
R58373 VINN.n400 VINN.n154 4.5005
R58374 VINN.n215 VINN.n154 4.5005
R58375 VINN.n654 VINN.n154 4.5005
R58376 VINN.n656 VINN.n154 4.5005
R58377 VINN.n154 VINN.n0 4.5005
R58378 VINN.n278 VINN.n146 4.5005
R58379 VINN.n276 VINN.n146 4.5005
R58380 VINN.n280 VINN.n146 4.5005
R58381 VINN.n275 VINN.n146 4.5005
R58382 VINN.n282 VINN.n146 4.5005
R58383 VINN.n274 VINN.n146 4.5005
R58384 VINN.n284 VINN.n146 4.5005
R58385 VINN.n273 VINN.n146 4.5005
R58386 VINN.n286 VINN.n146 4.5005
R58387 VINN.n272 VINN.n146 4.5005
R58388 VINN.n288 VINN.n146 4.5005
R58389 VINN.n271 VINN.n146 4.5005
R58390 VINN.n290 VINN.n146 4.5005
R58391 VINN.n270 VINN.n146 4.5005
R58392 VINN.n292 VINN.n146 4.5005
R58393 VINN.n269 VINN.n146 4.5005
R58394 VINN.n294 VINN.n146 4.5005
R58395 VINN.n268 VINN.n146 4.5005
R58396 VINN.n296 VINN.n146 4.5005
R58397 VINN.n267 VINN.n146 4.5005
R58398 VINN.n298 VINN.n146 4.5005
R58399 VINN.n266 VINN.n146 4.5005
R58400 VINN.n300 VINN.n146 4.5005
R58401 VINN.n265 VINN.n146 4.5005
R58402 VINN.n302 VINN.n146 4.5005
R58403 VINN.n264 VINN.n146 4.5005
R58404 VINN.n304 VINN.n146 4.5005
R58405 VINN.n263 VINN.n146 4.5005
R58406 VINN.n306 VINN.n146 4.5005
R58407 VINN.n262 VINN.n146 4.5005
R58408 VINN.n308 VINN.n146 4.5005
R58409 VINN.n261 VINN.n146 4.5005
R58410 VINN.n310 VINN.n146 4.5005
R58411 VINN.n260 VINN.n146 4.5005
R58412 VINN.n312 VINN.n146 4.5005
R58413 VINN.n259 VINN.n146 4.5005
R58414 VINN.n314 VINN.n146 4.5005
R58415 VINN.n258 VINN.n146 4.5005
R58416 VINN.n316 VINN.n146 4.5005
R58417 VINN.n257 VINN.n146 4.5005
R58418 VINN.n318 VINN.n146 4.5005
R58419 VINN.n256 VINN.n146 4.5005
R58420 VINN.n320 VINN.n146 4.5005
R58421 VINN.n255 VINN.n146 4.5005
R58422 VINN.n322 VINN.n146 4.5005
R58423 VINN.n254 VINN.n146 4.5005
R58424 VINN.n324 VINN.n146 4.5005
R58425 VINN.n253 VINN.n146 4.5005
R58426 VINN.n326 VINN.n146 4.5005
R58427 VINN.n252 VINN.n146 4.5005
R58428 VINN.n328 VINN.n146 4.5005
R58429 VINN.n251 VINN.n146 4.5005
R58430 VINN.n330 VINN.n146 4.5005
R58431 VINN.n250 VINN.n146 4.5005
R58432 VINN.n332 VINN.n146 4.5005
R58433 VINN.n249 VINN.n146 4.5005
R58434 VINN.n334 VINN.n146 4.5005
R58435 VINN.n248 VINN.n146 4.5005
R58436 VINN.n336 VINN.n146 4.5005
R58437 VINN.n247 VINN.n146 4.5005
R58438 VINN.n338 VINN.n146 4.5005
R58439 VINN.n246 VINN.n146 4.5005
R58440 VINN.n340 VINN.n146 4.5005
R58441 VINN.n245 VINN.n146 4.5005
R58442 VINN.n342 VINN.n146 4.5005
R58443 VINN.n244 VINN.n146 4.5005
R58444 VINN.n344 VINN.n146 4.5005
R58445 VINN.n243 VINN.n146 4.5005
R58446 VINN.n346 VINN.n146 4.5005
R58447 VINN.n242 VINN.n146 4.5005
R58448 VINN.n348 VINN.n146 4.5005
R58449 VINN.n241 VINN.n146 4.5005
R58450 VINN.n350 VINN.n146 4.5005
R58451 VINN.n240 VINN.n146 4.5005
R58452 VINN.n352 VINN.n146 4.5005
R58453 VINN.n239 VINN.n146 4.5005
R58454 VINN.n354 VINN.n146 4.5005
R58455 VINN.n238 VINN.n146 4.5005
R58456 VINN.n356 VINN.n146 4.5005
R58457 VINN.n237 VINN.n146 4.5005
R58458 VINN.n358 VINN.n146 4.5005
R58459 VINN.n236 VINN.n146 4.5005
R58460 VINN.n360 VINN.n146 4.5005
R58461 VINN.n235 VINN.n146 4.5005
R58462 VINN.n362 VINN.n146 4.5005
R58463 VINN.n234 VINN.n146 4.5005
R58464 VINN.n364 VINN.n146 4.5005
R58465 VINN.n233 VINN.n146 4.5005
R58466 VINN.n366 VINN.n146 4.5005
R58467 VINN.n232 VINN.n146 4.5005
R58468 VINN.n368 VINN.n146 4.5005
R58469 VINN.n231 VINN.n146 4.5005
R58470 VINN.n370 VINN.n146 4.5005
R58471 VINN.n230 VINN.n146 4.5005
R58472 VINN.n372 VINN.n146 4.5005
R58473 VINN.n229 VINN.n146 4.5005
R58474 VINN.n374 VINN.n146 4.5005
R58475 VINN.n228 VINN.n146 4.5005
R58476 VINN.n376 VINN.n146 4.5005
R58477 VINN.n227 VINN.n146 4.5005
R58478 VINN.n378 VINN.n146 4.5005
R58479 VINN.n226 VINN.n146 4.5005
R58480 VINN.n380 VINN.n146 4.5005
R58481 VINN.n225 VINN.n146 4.5005
R58482 VINN.n382 VINN.n146 4.5005
R58483 VINN.n224 VINN.n146 4.5005
R58484 VINN.n384 VINN.n146 4.5005
R58485 VINN.n223 VINN.n146 4.5005
R58486 VINN.n386 VINN.n146 4.5005
R58487 VINN.n222 VINN.n146 4.5005
R58488 VINN.n388 VINN.n146 4.5005
R58489 VINN.n221 VINN.n146 4.5005
R58490 VINN.n390 VINN.n146 4.5005
R58491 VINN.n220 VINN.n146 4.5005
R58492 VINN.n392 VINN.n146 4.5005
R58493 VINN.n219 VINN.n146 4.5005
R58494 VINN.n394 VINN.n146 4.5005
R58495 VINN.n218 VINN.n146 4.5005
R58496 VINN.n396 VINN.n146 4.5005
R58497 VINN.n217 VINN.n146 4.5005
R58498 VINN.n398 VINN.n146 4.5005
R58499 VINN.n216 VINN.n146 4.5005
R58500 VINN.n400 VINN.n146 4.5005
R58501 VINN.n215 VINN.n146 4.5005
R58502 VINN.n654 VINN.n146 4.5005
R58503 VINN.n656 VINN.n146 4.5005
R58504 VINN.n146 VINN.n0 4.5005
R58505 VINN.n278 VINN.n155 4.5005
R58506 VINN.n276 VINN.n155 4.5005
R58507 VINN.n280 VINN.n155 4.5005
R58508 VINN.n275 VINN.n155 4.5005
R58509 VINN.n282 VINN.n155 4.5005
R58510 VINN.n274 VINN.n155 4.5005
R58511 VINN.n284 VINN.n155 4.5005
R58512 VINN.n273 VINN.n155 4.5005
R58513 VINN.n286 VINN.n155 4.5005
R58514 VINN.n272 VINN.n155 4.5005
R58515 VINN.n288 VINN.n155 4.5005
R58516 VINN.n271 VINN.n155 4.5005
R58517 VINN.n290 VINN.n155 4.5005
R58518 VINN.n270 VINN.n155 4.5005
R58519 VINN.n292 VINN.n155 4.5005
R58520 VINN.n269 VINN.n155 4.5005
R58521 VINN.n294 VINN.n155 4.5005
R58522 VINN.n268 VINN.n155 4.5005
R58523 VINN.n296 VINN.n155 4.5005
R58524 VINN.n267 VINN.n155 4.5005
R58525 VINN.n298 VINN.n155 4.5005
R58526 VINN.n266 VINN.n155 4.5005
R58527 VINN.n300 VINN.n155 4.5005
R58528 VINN.n265 VINN.n155 4.5005
R58529 VINN.n302 VINN.n155 4.5005
R58530 VINN.n264 VINN.n155 4.5005
R58531 VINN.n304 VINN.n155 4.5005
R58532 VINN.n263 VINN.n155 4.5005
R58533 VINN.n306 VINN.n155 4.5005
R58534 VINN.n262 VINN.n155 4.5005
R58535 VINN.n308 VINN.n155 4.5005
R58536 VINN.n261 VINN.n155 4.5005
R58537 VINN.n310 VINN.n155 4.5005
R58538 VINN.n260 VINN.n155 4.5005
R58539 VINN.n312 VINN.n155 4.5005
R58540 VINN.n259 VINN.n155 4.5005
R58541 VINN.n314 VINN.n155 4.5005
R58542 VINN.n258 VINN.n155 4.5005
R58543 VINN.n316 VINN.n155 4.5005
R58544 VINN.n257 VINN.n155 4.5005
R58545 VINN.n318 VINN.n155 4.5005
R58546 VINN.n256 VINN.n155 4.5005
R58547 VINN.n320 VINN.n155 4.5005
R58548 VINN.n255 VINN.n155 4.5005
R58549 VINN.n322 VINN.n155 4.5005
R58550 VINN.n254 VINN.n155 4.5005
R58551 VINN.n324 VINN.n155 4.5005
R58552 VINN.n253 VINN.n155 4.5005
R58553 VINN.n326 VINN.n155 4.5005
R58554 VINN.n252 VINN.n155 4.5005
R58555 VINN.n328 VINN.n155 4.5005
R58556 VINN.n251 VINN.n155 4.5005
R58557 VINN.n330 VINN.n155 4.5005
R58558 VINN.n250 VINN.n155 4.5005
R58559 VINN.n332 VINN.n155 4.5005
R58560 VINN.n249 VINN.n155 4.5005
R58561 VINN.n334 VINN.n155 4.5005
R58562 VINN.n248 VINN.n155 4.5005
R58563 VINN.n336 VINN.n155 4.5005
R58564 VINN.n247 VINN.n155 4.5005
R58565 VINN.n338 VINN.n155 4.5005
R58566 VINN.n246 VINN.n155 4.5005
R58567 VINN.n340 VINN.n155 4.5005
R58568 VINN.n245 VINN.n155 4.5005
R58569 VINN.n342 VINN.n155 4.5005
R58570 VINN.n244 VINN.n155 4.5005
R58571 VINN.n344 VINN.n155 4.5005
R58572 VINN.n243 VINN.n155 4.5005
R58573 VINN.n346 VINN.n155 4.5005
R58574 VINN.n242 VINN.n155 4.5005
R58575 VINN.n348 VINN.n155 4.5005
R58576 VINN.n241 VINN.n155 4.5005
R58577 VINN.n350 VINN.n155 4.5005
R58578 VINN.n240 VINN.n155 4.5005
R58579 VINN.n352 VINN.n155 4.5005
R58580 VINN.n239 VINN.n155 4.5005
R58581 VINN.n354 VINN.n155 4.5005
R58582 VINN.n238 VINN.n155 4.5005
R58583 VINN.n356 VINN.n155 4.5005
R58584 VINN.n237 VINN.n155 4.5005
R58585 VINN.n358 VINN.n155 4.5005
R58586 VINN.n236 VINN.n155 4.5005
R58587 VINN.n360 VINN.n155 4.5005
R58588 VINN.n235 VINN.n155 4.5005
R58589 VINN.n362 VINN.n155 4.5005
R58590 VINN.n234 VINN.n155 4.5005
R58591 VINN.n364 VINN.n155 4.5005
R58592 VINN.n233 VINN.n155 4.5005
R58593 VINN.n366 VINN.n155 4.5005
R58594 VINN.n232 VINN.n155 4.5005
R58595 VINN.n368 VINN.n155 4.5005
R58596 VINN.n231 VINN.n155 4.5005
R58597 VINN.n370 VINN.n155 4.5005
R58598 VINN.n230 VINN.n155 4.5005
R58599 VINN.n372 VINN.n155 4.5005
R58600 VINN.n229 VINN.n155 4.5005
R58601 VINN.n374 VINN.n155 4.5005
R58602 VINN.n228 VINN.n155 4.5005
R58603 VINN.n376 VINN.n155 4.5005
R58604 VINN.n227 VINN.n155 4.5005
R58605 VINN.n378 VINN.n155 4.5005
R58606 VINN.n226 VINN.n155 4.5005
R58607 VINN.n380 VINN.n155 4.5005
R58608 VINN.n225 VINN.n155 4.5005
R58609 VINN.n382 VINN.n155 4.5005
R58610 VINN.n224 VINN.n155 4.5005
R58611 VINN.n384 VINN.n155 4.5005
R58612 VINN.n223 VINN.n155 4.5005
R58613 VINN.n386 VINN.n155 4.5005
R58614 VINN.n222 VINN.n155 4.5005
R58615 VINN.n388 VINN.n155 4.5005
R58616 VINN.n221 VINN.n155 4.5005
R58617 VINN.n390 VINN.n155 4.5005
R58618 VINN.n220 VINN.n155 4.5005
R58619 VINN.n392 VINN.n155 4.5005
R58620 VINN.n219 VINN.n155 4.5005
R58621 VINN.n394 VINN.n155 4.5005
R58622 VINN.n218 VINN.n155 4.5005
R58623 VINN.n396 VINN.n155 4.5005
R58624 VINN.n217 VINN.n155 4.5005
R58625 VINN.n398 VINN.n155 4.5005
R58626 VINN.n216 VINN.n155 4.5005
R58627 VINN.n400 VINN.n155 4.5005
R58628 VINN.n215 VINN.n155 4.5005
R58629 VINN.n654 VINN.n155 4.5005
R58630 VINN.n656 VINN.n155 4.5005
R58631 VINN.n155 VINN.n0 4.5005
R58632 VINN.n278 VINN.n145 4.5005
R58633 VINN.n276 VINN.n145 4.5005
R58634 VINN.n280 VINN.n145 4.5005
R58635 VINN.n275 VINN.n145 4.5005
R58636 VINN.n282 VINN.n145 4.5005
R58637 VINN.n274 VINN.n145 4.5005
R58638 VINN.n284 VINN.n145 4.5005
R58639 VINN.n273 VINN.n145 4.5005
R58640 VINN.n286 VINN.n145 4.5005
R58641 VINN.n272 VINN.n145 4.5005
R58642 VINN.n288 VINN.n145 4.5005
R58643 VINN.n271 VINN.n145 4.5005
R58644 VINN.n290 VINN.n145 4.5005
R58645 VINN.n270 VINN.n145 4.5005
R58646 VINN.n292 VINN.n145 4.5005
R58647 VINN.n269 VINN.n145 4.5005
R58648 VINN.n294 VINN.n145 4.5005
R58649 VINN.n268 VINN.n145 4.5005
R58650 VINN.n296 VINN.n145 4.5005
R58651 VINN.n267 VINN.n145 4.5005
R58652 VINN.n298 VINN.n145 4.5005
R58653 VINN.n266 VINN.n145 4.5005
R58654 VINN.n300 VINN.n145 4.5005
R58655 VINN.n265 VINN.n145 4.5005
R58656 VINN.n302 VINN.n145 4.5005
R58657 VINN.n264 VINN.n145 4.5005
R58658 VINN.n304 VINN.n145 4.5005
R58659 VINN.n263 VINN.n145 4.5005
R58660 VINN.n306 VINN.n145 4.5005
R58661 VINN.n262 VINN.n145 4.5005
R58662 VINN.n308 VINN.n145 4.5005
R58663 VINN.n261 VINN.n145 4.5005
R58664 VINN.n310 VINN.n145 4.5005
R58665 VINN.n260 VINN.n145 4.5005
R58666 VINN.n312 VINN.n145 4.5005
R58667 VINN.n259 VINN.n145 4.5005
R58668 VINN.n314 VINN.n145 4.5005
R58669 VINN.n258 VINN.n145 4.5005
R58670 VINN.n316 VINN.n145 4.5005
R58671 VINN.n257 VINN.n145 4.5005
R58672 VINN.n318 VINN.n145 4.5005
R58673 VINN.n256 VINN.n145 4.5005
R58674 VINN.n320 VINN.n145 4.5005
R58675 VINN.n255 VINN.n145 4.5005
R58676 VINN.n322 VINN.n145 4.5005
R58677 VINN.n254 VINN.n145 4.5005
R58678 VINN.n324 VINN.n145 4.5005
R58679 VINN.n253 VINN.n145 4.5005
R58680 VINN.n326 VINN.n145 4.5005
R58681 VINN.n252 VINN.n145 4.5005
R58682 VINN.n328 VINN.n145 4.5005
R58683 VINN.n251 VINN.n145 4.5005
R58684 VINN.n330 VINN.n145 4.5005
R58685 VINN.n250 VINN.n145 4.5005
R58686 VINN.n332 VINN.n145 4.5005
R58687 VINN.n249 VINN.n145 4.5005
R58688 VINN.n334 VINN.n145 4.5005
R58689 VINN.n248 VINN.n145 4.5005
R58690 VINN.n336 VINN.n145 4.5005
R58691 VINN.n247 VINN.n145 4.5005
R58692 VINN.n338 VINN.n145 4.5005
R58693 VINN.n246 VINN.n145 4.5005
R58694 VINN.n340 VINN.n145 4.5005
R58695 VINN.n245 VINN.n145 4.5005
R58696 VINN.n342 VINN.n145 4.5005
R58697 VINN.n244 VINN.n145 4.5005
R58698 VINN.n344 VINN.n145 4.5005
R58699 VINN.n243 VINN.n145 4.5005
R58700 VINN.n346 VINN.n145 4.5005
R58701 VINN.n242 VINN.n145 4.5005
R58702 VINN.n348 VINN.n145 4.5005
R58703 VINN.n241 VINN.n145 4.5005
R58704 VINN.n350 VINN.n145 4.5005
R58705 VINN.n240 VINN.n145 4.5005
R58706 VINN.n352 VINN.n145 4.5005
R58707 VINN.n239 VINN.n145 4.5005
R58708 VINN.n354 VINN.n145 4.5005
R58709 VINN.n238 VINN.n145 4.5005
R58710 VINN.n356 VINN.n145 4.5005
R58711 VINN.n237 VINN.n145 4.5005
R58712 VINN.n358 VINN.n145 4.5005
R58713 VINN.n236 VINN.n145 4.5005
R58714 VINN.n360 VINN.n145 4.5005
R58715 VINN.n235 VINN.n145 4.5005
R58716 VINN.n362 VINN.n145 4.5005
R58717 VINN.n234 VINN.n145 4.5005
R58718 VINN.n364 VINN.n145 4.5005
R58719 VINN.n233 VINN.n145 4.5005
R58720 VINN.n366 VINN.n145 4.5005
R58721 VINN.n232 VINN.n145 4.5005
R58722 VINN.n368 VINN.n145 4.5005
R58723 VINN.n231 VINN.n145 4.5005
R58724 VINN.n370 VINN.n145 4.5005
R58725 VINN.n230 VINN.n145 4.5005
R58726 VINN.n372 VINN.n145 4.5005
R58727 VINN.n229 VINN.n145 4.5005
R58728 VINN.n374 VINN.n145 4.5005
R58729 VINN.n228 VINN.n145 4.5005
R58730 VINN.n376 VINN.n145 4.5005
R58731 VINN.n227 VINN.n145 4.5005
R58732 VINN.n378 VINN.n145 4.5005
R58733 VINN.n226 VINN.n145 4.5005
R58734 VINN.n380 VINN.n145 4.5005
R58735 VINN.n225 VINN.n145 4.5005
R58736 VINN.n382 VINN.n145 4.5005
R58737 VINN.n224 VINN.n145 4.5005
R58738 VINN.n384 VINN.n145 4.5005
R58739 VINN.n223 VINN.n145 4.5005
R58740 VINN.n386 VINN.n145 4.5005
R58741 VINN.n222 VINN.n145 4.5005
R58742 VINN.n388 VINN.n145 4.5005
R58743 VINN.n221 VINN.n145 4.5005
R58744 VINN.n390 VINN.n145 4.5005
R58745 VINN.n220 VINN.n145 4.5005
R58746 VINN.n392 VINN.n145 4.5005
R58747 VINN.n219 VINN.n145 4.5005
R58748 VINN.n394 VINN.n145 4.5005
R58749 VINN.n218 VINN.n145 4.5005
R58750 VINN.n396 VINN.n145 4.5005
R58751 VINN.n217 VINN.n145 4.5005
R58752 VINN.n398 VINN.n145 4.5005
R58753 VINN.n216 VINN.n145 4.5005
R58754 VINN.n400 VINN.n145 4.5005
R58755 VINN.n215 VINN.n145 4.5005
R58756 VINN.n654 VINN.n145 4.5005
R58757 VINN.n656 VINN.n145 4.5005
R58758 VINN.n145 VINN.n0 4.5005
R58759 VINN.n278 VINN.n156 4.5005
R58760 VINN.n276 VINN.n156 4.5005
R58761 VINN.n280 VINN.n156 4.5005
R58762 VINN.n275 VINN.n156 4.5005
R58763 VINN.n282 VINN.n156 4.5005
R58764 VINN.n274 VINN.n156 4.5005
R58765 VINN.n284 VINN.n156 4.5005
R58766 VINN.n273 VINN.n156 4.5005
R58767 VINN.n286 VINN.n156 4.5005
R58768 VINN.n272 VINN.n156 4.5005
R58769 VINN.n288 VINN.n156 4.5005
R58770 VINN.n271 VINN.n156 4.5005
R58771 VINN.n290 VINN.n156 4.5005
R58772 VINN.n270 VINN.n156 4.5005
R58773 VINN.n292 VINN.n156 4.5005
R58774 VINN.n269 VINN.n156 4.5005
R58775 VINN.n294 VINN.n156 4.5005
R58776 VINN.n268 VINN.n156 4.5005
R58777 VINN.n296 VINN.n156 4.5005
R58778 VINN.n267 VINN.n156 4.5005
R58779 VINN.n298 VINN.n156 4.5005
R58780 VINN.n266 VINN.n156 4.5005
R58781 VINN.n300 VINN.n156 4.5005
R58782 VINN.n265 VINN.n156 4.5005
R58783 VINN.n302 VINN.n156 4.5005
R58784 VINN.n264 VINN.n156 4.5005
R58785 VINN.n304 VINN.n156 4.5005
R58786 VINN.n263 VINN.n156 4.5005
R58787 VINN.n306 VINN.n156 4.5005
R58788 VINN.n262 VINN.n156 4.5005
R58789 VINN.n308 VINN.n156 4.5005
R58790 VINN.n261 VINN.n156 4.5005
R58791 VINN.n310 VINN.n156 4.5005
R58792 VINN.n260 VINN.n156 4.5005
R58793 VINN.n312 VINN.n156 4.5005
R58794 VINN.n259 VINN.n156 4.5005
R58795 VINN.n314 VINN.n156 4.5005
R58796 VINN.n258 VINN.n156 4.5005
R58797 VINN.n316 VINN.n156 4.5005
R58798 VINN.n257 VINN.n156 4.5005
R58799 VINN.n318 VINN.n156 4.5005
R58800 VINN.n256 VINN.n156 4.5005
R58801 VINN.n320 VINN.n156 4.5005
R58802 VINN.n255 VINN.n156 4.5005
R58803 VINN.n322 VINN.n156 4.5005
R58804 VINN.n254 VINN.n156 4.5005
R58805 VINN.n324 VINN.n156 4.5005
R58806 VINN.n253 VINN.n156 4.5005
R58807 VINN.n326 VINN.n156 4.5005
R58808 VINN.n252 VINN.n156 4.5005
R58809 VINN.n328 VINN.n156 4.5005
R58810 VINN.n251 VINN.n156 4.5005
R58811 VINN.n330 VINN.n156 4.5005
R58812 VINN.n250 VINN.n156 4.5005
R58813 VINN.n332 VINN.n156 4.5005
R58814 VINN.n249 VINN.n156 4.5005
R58815 VINN.n334 VINN.n156 4.5005
R58816 VINN.n248 VINN.n156 4.5005
R58817 VINN.n336 VINN.n156 4.5005
R58818 VINN.n247 VINN.n156 4.5005
R58819 VINN.n338 VINN.n156 4.5005
R58820 VINN.n246 VINN.n156 4.5005
R58821 VINN.n340 VINN.n156 4.5005
R58822 VINN.n245 VINN.n156 4.5005
R58823 VINN.n342 VINN.n156 4.5005
R58824 VINN.n244 VINN.n156 4.5005
R58825 VINN.n344 VINN.n156 4.5005
R58826 VINN.n243 VINN.n156 4.5005
R58827 VINN.n346 VINN.n156 4.5005
R58828 VINN.n242 VINN.n156 4.5005
R58829 VINN.n348 VINN.n156 4.5005
R58830 VINN.n241 VINN.n156 4.5005
R58831 VINN.n350 VINN.n156 4.5005
R58832 VINN.n240 VINN.n156 4.5005
R58833 VINN.n352 VINN.n156 4.5005
R58834 VINN.n239 VINN.n156 4.5005
R58835 VINN.n354 VINN.n156 4.5005
R58836 VINN.n238 VINN.n156 4.5005
R58837 VINN.n356 VINN.n156 4.5005
R58838 VINN.n237 VINN.n156 4.5005
R58839 VINN.n358 VINN.n156 4.5005
R58840 VINN.n236 VINN.n156 4.5005
R58841 VINN.n360 VINN.n156 4.5005
R58842 VINN.n235 VINN.n156 4.5005
R58843 VINN.n362 VINN.n156 4.5005
R58844 VINN.n234 VINN.n156 4.5005
R58845 VINN.n364 VINN.n156 4.5005
R58846 VINN.n233 VINN.n156 4.5005
R58847 VINN.n366 VINN.n156 4.5005
R58848 VINN.n232 VINN.n156 4.5005
R58849 VINN.n368 VINN.n156 4.5005
R58850 VINN.n231 VINN.n156 4.5005
R58851 VINN.n370 VINN.n156 4.5005
R58852 VINN.n230 VINN.n156 4.5005
R58853 VINN.n372 VINN.n156 4.5005
R58854 VINN.n229 VINN.n156 4.5005
R58855 VINN.n374 VINN.n156 4.5005
R58856 VINN.n228 VINN.n156 4.5005
R58857 VINN.n376 VINN.n156 4.5005
R58858 VINN.n227 VINN.n156 4.5005
R58859 VINN.n378 VINN.n156 4.5005
R58860 VINN.n226 VINN.n156 4.5005
R58861 VINN.n380 VINN.n156 4.5005
R58862 VINN.n225 VINN.n156 4.5005
R58863 VINN.n382 VINN.n156 4.5005
R58864 VINN.n224 VINN.n156 4.5005
R58865 VINN.n384 VINN.n156 4.5005
R58866 VINN.n223 VINN.n156 4.5005
R58867 VINN.n386 VINN.n156 4.5005
R58868 VINN.n222 VINN.n156 4.5005
R58869 VINN.n388 VINN.n156 4.5005
R58870 VINN.n221 VINN.n156 4.5005
R58871 VINN.n390 VINN.n156 4.5005
R58872 VINN.n220 VINN.n156 4.5005
R58873 VINN.n392 VINN.n156 4.5005
R58874 VINN.n219 VINN.n156 4.5005
R58875 VINN.n394 VINN.n156 4.5005
R58876 VINN.n218 VINN.n156 4.5005
R58877 VINN.n396 VINN.n156 4.5005
R58878 VINN.n217 VINN.n156 4.5005
R58879 VINN.n398 VINN.n156 4.5005
R58880 VINN.n216 VINN.n156 4.5005
R58881 VINN.n400 VINN.n156 4.5005
R58882 VINN.n215 VINN.n156 4.5005
R58883 VINN.n654 VINN.n156 4.5005
R58884 VINN.n656 VINN.n156 4.5005
R58885 VINN.n156 VINN.n0 4.5005
R58886 VINN.n278 VINN.n144 4.5005
R58887 VINN.n276 VINN.n144 4.5005
R58888 VINN.n280 VINN.n144 4.5005
R58889 VINN.n275 VINN.n144 4.5005
R58890 VINN.n282 VINN.n144 4.5005
R58891 VINN.n274 VINN.n144 4.5005
R58892 VINN.n284 VINN.n144 4.5005
R58893 VINN.n273 VINN.n144 4.5005
R58894 VINN.n286 VINN.n144 4.5005
R58895 VINN.n272 VINN.n144 4.5005
R58896 VINN.n288 VINN.n144 4.5005
R58897 VINN.n271 VINN.n144 4.5005
R58898 VINN.n290 VINN.n144 4.5005
R58899 VINN.n270 VINN.n144 4.5005
R58900 VINN.n292 VINN.n144 4.5005
R58901 VINN.n269 VINN.n144 4.5005
R58902 VINN.n294 VINN.n144 4.5005
R58903 VINN.n268 VINN.n144 4.5005
R58904 VINN.n296 VINN.n144 4.5005
R58905 VINN.n267 VINN.n144 4.5005
R58906 VINN.n298 VINN.n144 4.5005
R58907 VINN.n266 VINN.n144 4.5005
R58908 VINN.n300 VINN.n144 4.5005
R58909 VINN.n265 VINN.n144 4.5005
R58910 VINN.n302 VINN.n144 4.5005
R58911 VINN.n264 VINN.n144 4.5005
R58912 VINN.n304 VINN.n144 4.5005
R58913 VINN.n263 VINN.n144 4.5005
R58914 VINN.n306 VINN.n144 4.5005
R58915 VINN.n262 VINN.n144 4.5005
R58916 VINN.n308 VINN.n144 4.5005
R58917 VINN.n261 VINN.n144 4.5005
R58918 VINN.n310 VINN.n144 4.5005
R58919 VINN.n260 VINN.n144 4.5005
R58920 VINN.n312 VINN.n144 4.5005
R58921 VINN.n259 VINN.n144 4.5005
R58922 VINN.n314 VINN.n144 4.5005
R58923 VINN.n258 VINN.n144 4.5005
R58924 VINN.n316 VINN.n144 4.5005
R58925 VINN.n257 VINN.n144 4.5005
R58926 VINN.n318 VINN.n144 4.5005
R58927 VINN.n256 VINN.n144 4.5005
R58928 VINN.n320 VINN.n144 4.5005
R58929 VINN.n255 VINN.n144 4.5005
R58930 VINN.n322 VINN.n144 4.5005
R58931 VINN.n254 VINN.n144 4.5005
R58932 VINN.n324 VINN.n144 4.5005
R58933 VINN.n253 VINN.n144 4.5005
R58934 VINN.n326 VINN.n144 4.5005
R58935 VINN.n252 VINN.n144 4.5005
R58936 VINN.n328 VINN.n144 4.5005
R58937 VINN.n251 VINN.n144 4.5005
R58938 VINN.n330 VINN.n144 4.5005
R58939 VINN.n250 VINN.n144 4.5005
R58940 VINN.n332 VINN.n144 4.5005
R58941 VINN.n249 VINN.n144 4.5005
R58942 VINN.n334 VINN.n144 4.5005
R58943 VINN.n248 VINN.n144 4.5005
R58944 VINN.n336 VINN.n144 4.5005
R58945 VINN.n247 VINN.n144 4.5005
R58946 VINN.n338 VINN.n144 4.5005
R58947 VINN.n246 VINN.n144 4.5005
R58948 VINN.n340 VINN.n144 4.5005
R58949 VINN.n245 VINN.n144 4.5005
R58950 VINN.n342 VINN.n144 4.5005
R58951 VINN.n244 VINN.n144 4.5005
R58952 VINN.n344 VINN.n144 4.5005
R58953 VINN.n243 VINN.n144 4.5005
R58954 VINN.n346 VINN.n144 4.5005
R58955 VINN.n242 VINN.n144 4.5005
R58956 VINN.n348 VINN.n144 4.5005
R58957 VINN.n241 VINN.n144 4.5005
R58958 VINN.n350 VINN.n144 4.5005
R58959 VINN.n240 VINN.n144 4.5005
R58960 VINN.n352 VINN.n144 4.5005
R58961 VINN.n239 VINN.n144 4.5005
R58962 VINN.n354 VINN.n144 4.5005
R58963 VINN.n238 VINN.n144 4.5005
R58964 VINN.n356 VINN.n144 4.5005
R58965 VINN.n237 VINN.n144 4.5005
R58966 VINN.n358 VINN.n144 4.5005
R58967 VINN.n236 VINN.n144 4.5005
R58968 VINN.n360 VINN.n144 4.5005
R58969 VINN.n235 VINN.n144 4.5005
R58970 VINN.n362 VINN.n144 4.5005
R58971 VINN.n234 VINN.n144 4.5005
R58972 VINN.n364 VINN.n144 4.5005
R58973 VINN.n233 VINN.n144 4.5005
R58974 VINN.n366 VINN.n144 4.5005
R58975 VINN.n232 VINN.n144 4.5005
R58976 VINN.n368 VINN.n144 4.5005
R58977 VINN.n231 VINN.n144 4.5005
R58978 VINN.n370 VINN.n144 4.5005
R58979 VINN.n230 VINN.n144 4.5005
R58980 VINN.n372 VINN.n144 4.5005
R58981 VINN.n229 VINN.n144 4.5005
R58982 VINN.n374 VINN.n144 4.5005
R58983 VINN.n228 VINN.n144 4.5005
R58984 VINN.n376 VINN.n144 4.5005
R58985 VINN.n227 VINN.n144 4.5005
R58986 VINN.n378 VINN.n144 4.5005
R58987 VINN.n226 VINN.n144 4.5005
R58988 VINN.n380 VINN.n144 4.5005
R58989 VINN.n225 VINN.n144 4.5005
R58990 VINN.n382 VINN.n144 4.5005
R58991 VINN.n224 VINN.n144 4.5005
R58992 VINN.n384 VINN.n144 4.5005
R58993 VINN.n223 VINN.n144 4.5005
R58994 VINN.n386 VINN.n144 4.5005
R58995 VINN.n222 VINN.n144 4.5005
R58996 VINN.n388 VINN.n144 4.5005
R58997 VINN.n221 VINN.n144 4.5005
R58998 VINN.n390 VINN.n144 4.5005
R58999 VINN.n220 VINN.n144 4.5005
R59000 VINN.n392 VINN.n144 4.5005
R59001 VINN.n219 VINN.n144 4.5005
R59002 VINN.n394 VINN.n144 4.5005
R59003 VINN.n218 VINN.n144 4.5005
R59004 VINN.n396 VINN.n144 4.5005
R59005 VINN.n217 VINN.n144 4.5005
R59006 VINN.n398 VINN.n144 4.5005
R59007 VINN.n216 VINN.n144 4.5005
R59008 VINN.n400 VINN.n144 4.5005
R59009 VINN.n215 VINN.n144 4.5005
R59010 VINN.n654 VINN.n144 4.5005
R59011 VINN.n656 VINN.n144 4.5005
R59012 VINN.n144 VINN.n0 4.5005
R59013 VINN.n278 VINN.n157 4.5005
R59014 VINN.n276 VINN.n157 4.5005
R59015 VINN.n280 VINN.n157 4.5005
R59016 VINN.n275 VINN.n157 4.5005
R59017 VINN.n282 VINN.n157 4.5005
R59018 VINN.n274 VINN.n157 4.5005
R59019 VINN.n284 VINN.n157 4.5005
R59020 VINN.n273 VINN.n157 4.5005
R59021 VINN.n286 VINN.n157 4.5005
R59022 VINN.n272 VINN.n157 4.5005
R59023 VINN.n288 VINN.n157 4.5005
R59024 VINN.n271 VINN.n157 4.5005
R59025 VINN.n290 VINN.n157 4.5005
R59026 VINN.n270 VINN.n157 4.5005
R59027 VINN.n292 VINN.n157 4.5005
R59028 VINN.n269 VINN.n157 4.5005
R59029 VINN.n294 VINN.n157 4.5005
R59030 VINN.n268 VINN.n157 4.5005
R59031 VINN.n296 VINN.n157 4.5005
R59032 VINN.n267 VINN.n157 4.5005
R59033 VINN.n298 VINN.n157 4.5005
R59034 VINN.n266 VINN.n157 4.5005
R59035 VINN.n300 VINN.n157 4.5005
R59036 VINN.n265 VINN.n157 4.5005
R59037 VINN.n302 VINN.n157 4.5005
R59038 VINN.n264 VINN.n157 4.5005
R59039 VINN.n304 VINN.n157 4.5005
R59040 VINN.n263 VINN.n157 4.5005
R59041 VINN.n306 VINN.n157 4.5005
R59042 VINN.n262 VINN.n157 4.5005
R59043 VINN.n308 VINN.n157 4.5005
R59044 VINN.n261 VINN.n157 4.5005
R59045 VINN.n310 VINN.n157 4.5005
R59046 VINN.n260 VINN.n157 4.5005
R59047 VINN.n312 VINN.n157 4.5005
R59048 VINN.n259 VINN.n157 4.5005
R59049 VINN.n314 VINN.n157 4.5005
R59050 VINN.n258 VINN.n157 4.5005
R59051 VINN.n316 VINN.n157 4.5005
R59052 VINN.n257 VINN.n157 4.5005
R59053 VINN.n318 VINN.n157 4.5005
R59054 VINN.n256 VINN.n157 4.5005
R59055 VINN.n320 VINN.n157 4.5005
R59056 VINN.n255 VINN.n157 4.5005
R59057 VINN.n322 VINN.n157 4.5005
R59058 VINN.n254 VINN.n157 4.5005
R59059 VINN.n324 VINN.n157 4.5005
R59060 VINN.n253 VINN.n157 4.5005
R59061 VINN.n326 VINN.n157 4.5005
R59062 VINN.n252 VINN.n157 4.5005
R59063 VINN.n328 VINN.n157 4.5005
R59064 VINN.n251 VINN.n157 4.5005
R59065 VINN.n330 VINN.n157 4.5005
R59066 VINN.n250 VINN.n157 4.5005
R59067 VINN.n332 VINN.n157 4.5005
R59068 VINN.n249 VINN.n157 4.5005
R59069 VINN.n334 VINN.n157 4.5005
R59070 VINN.n248 VINN.n157 4.5005
R59071 VINN.n336 VINN.n157 4.5005
R59072 VINN.n247 VINN.n157 4.5005
R59073 VINN.n338 VINN.n157 4.5005
R59074 VINN.n246 VINN.n157 4.5005
R59075 VINN.n340 VINN.n157 4.5005
R59076 VINN.n245 VINN.n157 4.5005
R59077 VINN.n342 VINN.n157 4.5005
R59078 VINN.n244 VINN.n157 4.5005
R59079 VINN.n344 VINN.n157 4.5005
R59080 VINN.n243 VINN.n157 4.5005
R59081 VINN.n346 VINN.n157 4.5005
R59082 VINN.n242 VINN.n157 4.5005
R59083 VINN.n348 VINN.n157 4.5005
R59084 VINN.n241 VINN.n157 4.5005
R59085 VINN.n350 VINN.n157 4.5005
R59086 VINN.n240 VINN.n157 4.5005
R59087 VINN.n352 VINN.n157 4.5005
R59088 VINN.n239 VINN.n157 4.5005
R59089 VINN.n354 VINN.n157 4.5005
R59090 VINN.n238 VINN.n157 4.5005
R59091 VINN.n356 VINN.n157 4.5005
R59092 VINN.n237 VINN.n157 4.5005
R59093 VINN.n358 VINN.n157 4.5005
R59094 VINN.n236 VINN.n157 4.5005
R59095 VINN.n360 VINN.n157 4.5005
R59096 VINN.n235 VINN.n157 4.5005
R59097 VINN.n362 VINN.n157 4.5005
R59098 VINN.n234 VINN.n157 4.5005
R59099 VINN.n364 VINN.n157 4.5005
R59100 VINN.n233 VINN.n157 4.5005
R59101 VINN.n366 VINN.n157 4.5005
R59102 VINN.n232 VINN.n157 4.5005
R59103 VINN.n368 VINN.n157 4.5005
R59104 VINN.n231 VINN.n157 4.5005
R59105 VINN.n370 VINN.n157 4.5005
R59106 VINN.n230 VINN.n157 4.5005
R59107 VINN.n372 VINN.n157 4.5005
R59108 VINN.n229 VINN.n157 4.5005
R59109 VINN.n374 VINN.n157 4.5005
R59110 VINN.n228 VINN.n157 4.5005
R59111 VINN.n376 VINN.n157 4.5005
R59112 VINN.n227 VINN.n157 4.5005
R59113 VINN.n378 VINN.n157 4.5005
R59114 VINN.n226 VINN.n157 4.5005
R59115 VINN.n380 VINN.n157 4.5005
R59116 VINN.n225 VINN.n157 4.5005
R59117 VINN.n382 VINN.n157 4.5005
R59118 VINN.n224 VINN.n157 4.5005
R59119 VINN.n384 VINN.n157 4.5005
R59120 VINN.n223 VINN.n157 4.5005
R59121 VINN.n386 VINN.n157 4.5005
R59122 VINN.n222 VINN.n157 4.5005
R59123 VINN.n388 VINN.n157 4.5005
R59124 VINN.n221 VINN.n157 4.5005
R59125 VINN.n390 VINN.n157 4.5005
R59126 VINN.n220 VINN.n157 4.5005
R59127 VINN.n392 VINN.n157 4.5005
R59128 VINN.n219 VINN.n157 4.5005
R59129 VINN.n394 VINN.n157 4.5005
R59130 VINN.n218 VINN.n157 4.5005
R59131 VINN.n396 VINN.n157 4.5005
R59132 VINN.n217 VINN.n157 4.5005
R59133 VINN.n398 VINN.n157 4.5005
R59134 VINN.n216 VINN.n157 4.5005
R59135 VINN.n400 VINN.n157 4.5005
R59136 VINN.n215 VINN.n157 4.5005
R59137 VINN.n654 VINN.n157 4.5005
R59138 VINN.n656 VINN.n157 4.5005
R59139 VINN.n157 VINN.n0 4.5005
R59140 VINN.n278 VINN.n143 4.5005
R59141 VINN.n276 VINN.n143 4.5005
R59142 VINN.n280 VINN.n143 4.5005
R59143 VINN.n275 VINN.n143 4.5005
R59144 VINN.n282 VINN.n143 4.5005
R59145 VINN.n274 VINN.n143 4.5005
R59146 VINN.n284 VINN.n143 4.5005
R59147 VINN.n273 VINN.n143 4.5005
R59148 VINN.n286 VINN.n143 4.5005
R59149 VINN.n272 VINN.n143 4.5005
R59150 VINN.n288 VINN.n143 4.5005
R59151 VINN.n271 VINN.n143 4.5005
R59152 VINN.n290 VINN.n143 4.5005
R59153 VINN.n270 VINN.n143 4.5005
R59154 VINN.n292 VINN.n143 4.5005
R59155 VINN.n269 VINN.n143 4.5005
R59156 VINN.n294 VINN.n143 4.5005
R59157 VINN.n268 VINN.n143 4.5005
R59158 VINN.n296 VINN.n143 4.5005
R59159 VINN.n267 VINN.n143 4.5005
R59160 VINN.n298 VINN.n143 4.5005
R59161 VINN.n266 VINN.n143 4.5005
R59162 VINN.n300 VINN.n143 4.5005
R59163 VINN.n265 VINN.n143 4.5005
R59164 VINN.n302 VINN.n143 4.5005
R59165 VINN.n264 VINN.n143 4.5005
R59166 VINN.n304 VINN.n143 4.5005
R59167 VINN.n263 VINN.n143 4.5005
R59168 VINN.n306 VINN.n143 4.5005
R59169 VINN.n262 VINN.n143 4.5005
R59170 VINN.n308 VINN.n143 4.5005
R59171 VINN.n261 VINN.n143 4.5005
R59172 VINN.n310 VINN.n143 4.5005
R59173 VINN.n260 VINN.n143 4.5005
R59174 VINN.n312 VINN.n143 4.5005
R59175 VINN.n259 VINN.n143 4.5005
R59176 VINN.n314 VINN.n143 4.5005
R59177 VINN.n258 VINN.n143 4.5005
R59178 VINN.n316 VINN.n143 4.5005
R59179 VINN.n257 VINN.n143 4.5005
R59180 VINN.n318 VINN.n143 4.5005
R59181 VINN.n256 VINN.n143 4.5005
R59182 VINN.n320 VINN.n143 4.5005
R59183 VINN.n255 VINN.n143 4.5005
R59184 VINN.n322 VINN.n143 4.5005
R59185 VINN.n254 VINN.n143 4.5005
R59186 VINN.n324 VINN.n143 4.5005
R59187 VINN.n253 VINN.n143 4.5005
R59188 VINN.n326 VINN.n143 4.5005
R59189 VINN.n252 VINN.n143 4.5005
R59190 VINN.n328 VINN.n143 4.5005
R59191 VINN.n251 VINN.n143 4.5005
R59192 VINN.n330 VINN.n143 4.5005
R59193 VINN.n250 VINN.n143 4.5005
R59194 VINN.n332 VINN.n143 4.5005
R59195 VINN.n249 VINN.n143 4.5005
R59196 VINN.n334 VINN.n143 4.5005
R59197 VINN.n248 VINN.n143 4.5005
R59198 VINN.n336 VINN.n143 4.5005
R59199 VINN.n247 VINN.n143 4.5005
R59200 VINN.n338 VINN.n143 4.5005
R59201 VINN.n246 VINN.n143 4.5005
R59202 VINN.n340 VINN.n143 4.5005
R59203 VINN.n245 VINN.n143 4.5005
R59204 VINN.n342 VINN.n143 4.5005
R59205 VINN.n244 VINN.n143 4.5005
R59206 VINN.n344 VINN.n143 4.5005
R59207 VINN.n243 VINN.n143 4.5005
R59208 VINN.n346 VINN.n143 4.5005
R59209 VINN.n242 VINN.n143 4.5005
R59210 VINN.n348 VINN.n143 4.5005
R59211 VINN.n241 VINN.n143 4.5005
R59212 VINN.n350 VINN.n143 4.5005
R59213 VINN.n240 VINN.n143 4.5005
R59214 VINN.n352 VINN.n143 4.5005
R59215 VINN.n239 VINN.n143 4.5005
R59216 VINN.n354 VINN.n143 4.5005
R59217 VINN.n238 VINN.n143 4.5005
R59218 VINN.n356 VINN.n143 4.5005
R59219 VINN.n237 VINN.n143 4.5005
R59220 VINN.n358 VINN.n143 4.5005
R59221 VINN.n236 VINN.n143 4.5005
R59222 VINN.n360 VINN.n143 4.5005
R59223 VINN.n235 VINN.n143 4.5005
R59224 VINN.n362 VINN.n143 4.5005
R59225 VINN.n234 VINN.n143 4.5005
R59226 VINN.n364 VINN.n143 4.5005
R59227 VINN.n233 VINN.n143 4.5005
R59228 VINN.n366 VINN.n143 4.5005
R59229 VINN.n232 VINN.n143 4.5005
R59230 VINN.n368 VINN.n143 4.5005
R59231 VINN.n231 VINN.n143 4.5005
R59232 VINN.n370 VINN.n143 4.5005
R59233 VINN.n230 VINN.n143 4.5005
R59234 VINN.n372 VINN.n143 4.5005
R59235 VINN.n229 VINN.n143 4.5005
R59236 VINN.n374 VINN.n143 4.5005
R59237 VINN.n228 VINN.n143 4.5005
R59238 VINN.n376 VINN.n143 4.5005
R59239 VINN.n227 VINN.n143 4.5005
R59240 VINN.n378 VINN.n143 4.5005
R59241 VINN.n226 VINN.n143 4.5005
R59242 VINN.n380 VINN.n143 4.5005
R59243 VINN.n225 VINN.n143 4.5005
R59244 VINN.n382 VINN.n143 4.5005
R59245 VINN.n224 VINN.n143 4.5005
R59246 VINN.n384 VINN.n143 4.5005
R59247 VINN.n223 VINN.n143 4.5005
R59248 VINN.n386 VINN.n143 4.5005
R59249 VINN.n222 VINN.n143 4.5005
R59250 VINN.n388 VINN.n143 4.5005
R59251 VINN.n221 VINN.n143 4.5005
R59252 VINN.n390 VINN.n143 4.5005
R59253 VINN.n220 VINN.n143 4.5005
R59254 VINN.n392 VINN.n143 4.5005
R59255 VINN.n219 VINN.n143 4.5005
R59256 VINN.n394 VINN.n143 4.5005
R59257 VINN.n218 VINN.n143 4.5005
R59258 VINN.n396 VINN.n143 4.5005
R59259 VINN.n217 VINN.n143 4.5005
R59260 VINN.n398 VINN.n143 4.5005
R59261 VINN.n216 VINN.n143 4.5005
R59262 VINN.n400 VINN.n143 4.5005
R59263 VINN.n215 VINN.n143 4.5005
R59264 VINN.n654 VINN.n143 4.5005
R59265 VINN.n656 VINN.n143 4.5005
R59266 VINN.n143 VINN.n0 4.5005
R59267 VINN.n278 VINN.n158 4.5005
R59268 VINN.n276 VINN.n158 4.5005
R59269 VINN.n280 VINN.n158 4.5005
R59270 VINN.n275 VINN.n158 4.5005
R59271 VINN.n282 VINN.n158 4.5005
R59272 VINN.n274 VINN.n158 4.5005
R59273 VINN.n284 VINN.n158 4.5005
R59274 VINN.n273 VINN.n158 4.5005
R59275 VINN.n286 VINN.n158 4.5005
R59276 VINN.n272 VINN.n158 4.5005
R59277 VINN.n288 VINN.n158 4.5005
R59278 VINN.n271 VINN.n158 4.5005
R59279 VINN.n290 VINN.n158 4.5005
R59280 VINN.n270 VINN.n158 4.5005
R59281 VINN.n292 VINN.n158 4.5005
R59282 VINN.n269 VINN.n158 4.5005
R59283 VINN.n294 VINN.n158 4.5005
R59284 VINN.n268 VINN.n158 4.5005
R59285 VINN.n296 VINN.n158 4.5005
R59286 VINN.n267 VINN.n158 4.5005
R59287 VINN.n298 VINN.n158 4.5005
R59288 VINN.n266 VINN.n158 4.5005
R59289 VINN.n300 VINN.n158 4.5005
R59290 VINN.n265 VINN.n158 4.5005
R59291 VINN.n302 VINN.n158 4.5005
R59292 VINN.n264 VINN.n158 4.5005
R59293 VINN.n304 VINN.n158 4.5005
R59294 VINN.n263 VINN.n158 4.5005
R59295 VINN.n306 VINN.n158 4.5005
R59296 VINN.n262 VINN.n158 4.5005
R59297 VINN.n308 VINN.n158 4.5005
R59298 VINN.n261 VINN.n158 4.5005
R59299 VINN.n310 VINN.n158 4.5005
R59300 VINN.n260 VINN.n158 4.5005
R59301 VINN.n312 VINN.n158 4.5005
R59302 VINN.n259 VINN.n158 4.5005
R59303 VINN.n314 VINN.n158 4.5005
R59304 VINN.n258 VINN.n158 4.5005
R59305 VINN.n316 VINN.n158 4.5005
R59306 VINN.n257 VINN.n158 4.5005
R59307 VINN.n318 VINN.n158 4.5005
R59308 VINN.n256 VINN.n158 4.5005
R59309 VINN.n320 VINN.n158 4.5005
R59310 VINN.n255 VINN.n158 4.5005
R59311 VINN.n322 VINN.n158 4.5005
R59312 VINN.n254 VINN.n158 4.5005
R59313 VINN.n324 VINN.n158 4.5005
R59314 VINN.n253 VINN.n158 4.5005
R59315 VINN.n326 VINN.n158 4.5005
R59316 VINN.n252 VINN.n158 4.5005
R59317 VINN.n328 VINN.n158 4.5005
R59318 VINN.n251 VINN.n158 4.5005
R59319 VINN.n330 VINN.n158 4.5005
R59320 VINN.n250 VINN.n158 4.5005
R59321 VINN.n332 VINN.n158 4.5005
R59322 VINN.n249 VINN.n158 4.5005
R59323 VINN.n334 VINN.n158 4.5005
R59324 VINN.n248 VINN.n158 4.5005
R59325 VINN.n336 VINN.n158 4.5005
R59326 VINN.n247 VINN.n158 4.5005
R59327 VINN.n338 VINN.n158 4.5005
R59328 VINN.n246 VINN.n158 4.5005
R59329 VINN.n340 VINN.n158 4.5005
R59330 VINN.n245 VINN.n158 4.5005
R59331 VINN.n342 VINN.n158 4.5005
R59332 VINN.n244 VINN.n158 4.5005
R59333 VINN.n344 VINN.n158 4.5005
R59334 VINN.n243 VINN.n158 4.5005
R59335 VINN.n346 VINN.n158 4.5005
R59336 VINN.n242 VINN.n158 4.5005
R59337 VINN.n348 VINN.n158 4.5005
R59338 VINN.n241 VINN.n158 4.5005
R59339 VINN.n350 VINN.n158 4.5005
R59340 VINN.n240 VINN.n158 4.5005
R59341 VINN.n352 VINN.n158 4.5005
R59342 VINN.n239 VINN.n158 4.5005
R59343 VINN.n354 VINN.n158 4.5005
R59344 VINN.n238 VINN.n158 4.5005
R59345 VINN.n356 VINN.n158 4.5005
R59346 VINN.n237 VINN.n158 4.5005
R59347 VINN.n358 VINN.n158 4.5005
R59348 VINN.n236 VINN.n158 4.5005
R59349 VINN.n360 VINN.n158 4.5005
R59350 VINN.n235 VINN.n158 4.5005
R59351 VINN.n362 VINN.n158 4.5005
R59352 VINN.n234 VINN.n158 4.5005
R59353 VINN.n364 VINN.n158 4.5005
R59354 VINN.n233 VINN.n158 4.5005
R59355 VINN.n366 VINN.n158 4.5005
R59356 VINN.n232 VINN.n158 4.5005
R59357 VINN.n368 VINN.n158 4.5005
R59358 VINN.n231 VINN.n158 4.5005
R59359 VINN.n370 VINN.n158 4.5005
R59360 VINN.n230 VINN.n158 4.5005
R59361 VINN.n372 VINN.n158 4.5005
R59362 VINN.n229 VINN.n158 4.5005
R59363 VINN.n374 VINN.n158 4.5005
R59364 VINN.n228 VINN.n158 4.5005
R59365 VINN.n376 VINN.n158 4.5005
R59366 VINN.n227 VINN.n158 4.5005
R59367 VINN.n378 VINN.n158 4.5005
R59368 VINN.n226 VINN.n158 4.5005
R59369 VINN.n380 VINN.n158 4.5005
R59370 VINN.n225 VINN.n158 4.5005
R59371 VINN.n382 VINN.n158 4.5005
R59372 VINN.n224 VINN.n158 4.5005
R59373 VINN.n384 VINN.n158 4.5005
R59374 VINN.n223 VINN.n158 4.5005
R59375 VINN.n386 VINN.n158 4.5005
R59376 VINN.n222 VINN.n158 4.5005
R59377 VINN.n388 VINN.n158 4.5005
R59378 VINN.n221 VINN.n158 4.5005
R59379 VINN.n390 VINN.n158 4.5005
R59380 VINN.n220 VINN.n158 4.5005
R59381 VINN.n392 VINN.n158 4.5005
R59382 VINN.n219 VINN.n158 4.5005
R59383 VINN.n394 VINN.n158 4.5005
R59384 VINN.n218 VINN.n158 4.5005
R59385 VINN.n396 VINN.n158 4.5005
R59386 VINN.n217 VINN.n158 4.5005
R59387 VINN.n398 VINN.n158 4.5005
R59388 VINN.n216 VINN.n158 4.5005
R59389 VINN.n400 VINN.n158 4.5005
R59390 VINN.n215 VINN.n158 4.5005
R59391 VINN.n654 VINN.n158 4.5005
R59392 VINN.n656 VINN.n158 4.5005
R59393 VINN.n158 VINN.n0 4.5005
R59394 VINN.n278 VINN.n142 4.5005
R59395 VINN.n276 VINN.n142 4.5005
R59396 VINN.n280 VINN.n142 4.5005
R59397 VINN.n275 VINN.n142 4.5005
R59398 VINN.n282 VINN.n142 4.5005
R59399 VINN.n274 VINN.n142 4.5005
R59400 VINN.n284 VINN.n142 4.5005
R59401 VINN.n273 VINN.n142 4.5005
R59402 VINN.n286 VINN.n142 4.5005
R59403 VINN.n272 VINN.n142 4.5005
R59404 VINN.n288 VINN.n142 4.5005
R59405 VINN.n271 VINN.n142 4.5005
R59406 VINN.n290 VINN.n142 4.5005
R59407 VINN.n270 VINN.n142 4.5005
R59408 VINN.n292 VINN.n142 4.5005
R59409 VINN.n269 VINN.n142 4.5005
R59410 VINN.n294 VINN.n142 4.5005
R59411 VINN.n268 VINN.n142 4.5005
R59412 VINN.n296 VINN.n142 4.5005
R59413 VINN.n267 VINN.n142 4.5005
R59414 VINN.n298 VINN.n142 4.5005
R59415 VINN.n266 VINN.n142 4.5005
R59416 VINN.n300 VINN.n142 4.5005
R59417 VINN.n265 VINN.n142 4.5005
R59418 VINN.n302 VINN.n142 4.5005
R59419 VINN.n264 VINN.n142 4.5005
R59420 VINN.n304 VINN.n142 4.5005
R59421 VINN.n263 VINN.n142 4.5005
R59422 VINN.n306 VINN.n142 4.5005
R59423 VINN.n262 VINN.n142 4.5005
R59424 VINN.n308 VINN.n142 4.5005
R59425 VINN.n261 VINN.n142 4.5005
R59426 VINN.n310 VINN.n142 4.5005
R59427 VINN.n260 VINN.n142 4.5005
R59428 VINN.n312 VINN.n142 4.5005
R59429 VINN.n259 VINN.n142 4.5005
R59430 VINN.n314 VINN.n142 4.5005
R59431 VINN.n258 VINN.n142 4.5005
R59432 VINN.n316 VINN.n142 4.5005
R59433 VINN.n257 VINN.n142 4.5005
R59434 VINN.n318 VINN.n142 4.5005
R59435 VINN.n256 VINN.n142 4.5005
R59436 VINN.n320 VINN.n142 4.5005
R59437 VINN.n255 VINN.n142 4.5005
R59438 VINN.n322 VINN.n142 4.5005
R59439 VINN.n254 VINN.n142 4.5005
R59440 VINN.n324 VINN.n142 4.5005
R59441 VINN.n253 VINN.n142 4.5005
R59442 VINN.n326 VINN.n142 4.5005
R59443 VINN.n252 VINN.n142 4.5005
R59444 VINN.n328 VINN.n142 4.5005
R59445 VINN.n251 VINN.n142 4.5005
R59446 VINN.n330 VINN.n142 4.5005
R59447 VINN.n250 VINN.n142 4.5005
R59448 VINN.n332 VINN.n142 4.5005
R59449 VINN.n249 VINN.n142 4.5005
R59450 VINN.n334 VINN.n142 4.5005
R59451 VINN.n248 VINN.n142 4.5005
R59452 VINN.n336 VINN.n142 4.5005
R59453 VINN.n247 VINN.n142 4.5005
R59454 VINN.n338 VINN.n142 4.5005
R59455 VINN.n246 VINN.n142 4.5005
R59456 VINN.n340 VINN.n142 4.5005
R59457 VINN.n245 VINN.n142 4.5005
R59458 VINN.n342 VINN.n142 4.5005
R59459 VINN.n244 VINN.n142 4.5005
R59460 VINN.n344 VINN.n142 4.5005
R59461 VINN.n243 VINN.n142 4.5005
R59462 VINN.n346 VINN.n142 4.5005
R59463 VINN.n242 VINN.n142 4.5005
R59464 VINN.n348 VINN.n142 4.5005
R59465 VINN.n241 VINN.n142 4.5005
R59466 VINN.n350 VINN.n142 4.5005
R59467 VINN.n240 VINN.n142 4.5005
R59468 VINN.n352 VINN.n142 4.5005
R59469 VINN.n239 VINN.n142 4.5005
R59470 VINN.n354 VINN.n142 4.5005
R59471 VINN.n238 VINN.n142 4.5005
R59472 VINN.n356 VINN.n142 4.5005
R59473 VINN.n237 VINN.n142 4.5005
R59474 VINN.n358 VINN.n142 4.5005
R59475 VINN.n236 VINN.n142 4.5005
R59476 VINN.n360 VINN.n142 4.5005
R59477 VINN.n235 VINN.n142 4.5005
R59478 VINN.n362 VINN.n142 4.5005
R59479 VINN.n234 VINN.n142 4.5005
R59480 VINN.n364 VINN.n142 4.5005
R59481 VINN.n233 VINN.n142 4.5005
R59482 VINN.n366 VINN.n142 4.5005
R59483 VINN.n232 VINN.n142 4.5005
R59484 VINN.n368 VINN.n142 4.5005
R59485 VINN.n231 VINN.n142 4.5005
R59486 VINN.n370 VINN.n142 4.5005
R59487 VINN.n230 VINN.n142 4.5005
R59488 VINN.n372 VINN.n142 4.5005
R59489 VINN.n229 VINN.n142 4.5005
R59490 VINN.n374 VINN.n142 4.5005
R59491 VINN.n228 VINN.n142 4.5005
R59492 VINN.n376 VINN.n142 4.5005
R59493 VINN.n227 VINN.n142 4.5005
R59494 VINN.n378 VINN.n142 4.5005
R59495 VINN.n226 VINN.n142 4.5005
R59496 VINN.n380 VINN.n142 4.5005
R59497 VINN.n225 VINN.n142 4.5005
R59498 VINN.n382 VINN.n142 4.5005
R59499 VINN.n224 VINN.n142 4.5005
R59500 VINN.n384 VINN.n142 4.5005
R59501 VINN.n223 VINN.n142 4.5005
R59502 VINN.n386 VINN.n142 4.5005
R59503 VINN.n222 VINN.n142 4.5005
R59504 VINN.n388 VINN.n142 4.5005
R59505 VINN.n221 VINN.n142 4.5005
R59506 VINN.n390 VINN.n142 4.5005
R59507 VINN.n220 VINN.n142 4.5005
R59508 VINN.n392 VINN.n142 4.5005
R59509 VINN.n219 VINN.n142 4.5005
R59510 VINN.n394 VINN.n142 4.5005
R59511 VINN.n218 VINN.n142 4.5005
R59512 VINN.n396 VINN.n142 4.5005
R59513 VINN.n217 VINN.n142 4.5005
R59514 VINN.n398 VINN.n142 4.5005
R59515 VINN.n216 VINN.n142 4.5005
R59516 VINN.n400 VINN.n142 4.5005
R59517 VINN.n215 VINN.n142 4.5005
R59518 VINN.n654 VINN.n142 4.5005
R59519 VINN.n656 VINN.n142 4.5005
R59520 VINN.n142 VINN.n0 4.5005
R59521 VINN.n278 VINN.n159 4.5005
R59522 VINN.n276 VINN.n159 4.5005
R59523 VINN.n280 VINN.n159 4.5005
R59524 VINN.n275 VINN.n159 4.5005
R59525 VINN.n282 VINN.n159 4.5005
R59526 VINN.n274 VINN.n159 4.5005
R59527 VINN.n284 VINN.n159 4.5005
R59528 VINN.n273 VINN.n159 4.5005
R59529 VINN.n286 VINN.n159 4.5005
R59530 VINN.n272 VINN.n159 4.5005
R59531 VINN.n288 VINN.n159 4.5005
R59532 VINN.n271 VINN.n159 4.5005
R59533 VINN.n290 VINN.n159 4.5005
R59534 VINN.n270 VINN.n159 4.5005
R59535 VINN.n292 VINN.n159 4.5005
R59536 VINN.n269 VINN.n159 4.5005
R59537 VINN.n294 VINN.n159 4.5005
R59538 VINN.n268 VINN.n159 4.5005
R59539 VINN.n296 VINN.n159 4.5005
R59540 VINN.n267 VINN.n159 4.5005
R59541 VINN.n298 VINN.n159 4.5005
R59542 VINN.n266 VINN.n159 4.5005
R59543 VINN.n300 VINN.n159 4.5005
R59544 VINN.n265 VINN.n159 4.5005
R59545 VINN.n302 VINN.n159 4.5005
R59546 VINN.n264 VINN.n159 4.5005
R59547 VINN.n304 VINN.n159 4.5005
R59548 VINN.n263 VINN.n159 4.5005
R59549 VINN.n306 VINN.n159 4.5005
R59550 VINN.n262 VINN.n159 4.5005
R59551 VINN.n308 VINN.n159 4.5005
R59552 VINN.n261 VINN.n159 4.5005
R59553 VINN.n310 VINN.n159 4.5005
R59554 VINN.n260 VINN.n159 4.5005
R59555 VINN.n312 VINN.n159 4.5005
R59556 VINN.n259 VINN.n159 4.5005
R59557 VINN.n314 VINN.n159 4.5005
R59558 VINN.n258 VINN.n159 4.5005
R59559 VINN.n316 VINN.n159 4.5005
R59560 VINN.n257 VINN.n159 4.5005
R59561 VINN.n318 VINN.n159 4.5005
R59562 VINN.n256 VINN.n159 4.5005
R59563 VINN.n320 VINN.n159 4.5005
R59564 VINN.n255 VINN.n159 4.5005
R59565 VINN.n322 VINN.n159 4.5005
R59566 VINN.n254 VINN.n159 4.5005
R59567 VINN.n324 VINN.n159 4.5005
R59568 VINN.n253 VINN.n159 4.5005
R59569 VINN.n326 VINN.n159 4.5005
R59570 VINN.n252 VINN.n159 4.5005
R59571 VINN.n328 VINN.n159 4.5005
R59572 VINN.n251 VINN.n159 4.5005
R59573 VINN.n330 VINN.n159 4.5005
R59574 VINN.n250 VINN.n159 4.5005
R59575 VINN.n332 VINN.n159 4.5005
R59576 VINN.n249 VINN.n159 4.5005
R59577 VINN.n334 VINN.n159 4.5005
R59578 VINN.n248 VINN.n159 4.5005
R59579 VINN.n336 VINN.n159 4.5005
R59580 VINN.n247 VINN.n159 4.5005
R59581 VINN.n338 VINN.n159 4.5005
R59582 VINN.n246 VINN.n159 4.5005
R59583 VINN.n340 VINN.n159 4.5005
R59584 VINN.n245 VINN.n159 4.5005
R59585 VINN.n342 VINN.n159 4.5005
R59586 VINN.n244 VINN.n159 4.5005
R59587 VINN.n344 VINN.n159 4.5005
R59588 VINN.n243 VINN.n159 4.5005
R59589 VINN.n346 VINN.n159 4.5005
R59590 VINN.n242 VINN.n159 4.5005
R59591 VINN.n348 VINN.n159 4.5005
R59592 VINN.n241 VINN.n159 4.5005
R59593 VINN.n350 VINN.n159 4.5005
R59594 VINN.n240 VINN.n159 4.5005
R59595 VINN.n352 VINN.n159 4.5005
R59596 VINN.n239 VINN.n159 4.5005
R59597 VINN.n354 VINN.n159 4.5005
R59598 VINN.n238 VINN.n159 4.5005
R59599 VINN.n356 VINN.n159 4.5005
R59600 VINN.n237 VINN.n159 4.5005
R59601 VINN.n358 VINN.n159 4.5005
R59602 VINN.n236 VINN.n159 4.5005
R59603 VINN.n360 VINN.n159 4.5005
R59604 VINN.n235 VINN.n159 4.5005
R59605 VINN.n362 VINN.n159 4.5005
R59606 VINN.n234 VINN.n159 4.5005
R59607 VINN.n364 VINN.n159 4.5005
R59608 VINN.n233 VINN.n159 4.5005
R59609 VINN.n366 VINN.n159 4.5005
R59610 VINN.n232 VINN.n159 4.5005
R59611 VINN.n368 VINN.n159 4.5005
R59612 VINN.n231 VINN.n159 4.5005
R59613 VINN.n370 VINN.n159 4.5005
R59614 VINN.n230 VINN.n159 4.5005
R59615 VINN.n372 VINN.n159 4.5005
R59616 VINN.n229 VINN.n159 4.5005
R59617 VINN.n374 VINN.n159 4.5005
R59618 VINN.n228 VINN.n159 4.5005
R59619 VINN.n376 VINN.n159 4.5005
R59620 VINN.n227 VINN.n159 4.5005
R59621 VINN.n378 VINN.n159 4.5005
R59622 VINN.n226 VINN.n159 4.5005
R59623 VINN.n380 VINN.n159 4.5005
R59624 VINN.n225 VINN.n159 4.5005
R59625 VINN.n382 VINN.n159 4.5005
R59626 VINN.n224 VINN.n159 4.5005
R59627 VINN.n384 VINN.n159 4.5005
R59628 VINN.n223 VINN.n159 4.5005
R59629 VINN.n386 VINN.n159 4.5005
R59630 VINN.n222 VINN.n159 4.5005
R59631 VINN.n388 VINN.n159 4.5005
R59632 VINN.n221 VINN.n159 4.5005
R59633 VINN.n390 VINN.n159 4.5005
R59634 VINN.n220 VINN.n159 4.5005
R59635 VINN.n392 VINN.n159 4.5005
R59636 VINN.n219 VINN.n159 4.5005
R59637 VINN.n394 VINN.n159 4.5005
R59638 VINN.n218 VINN.n159 4.5005
R59639 VINN.n396 VINN.n159 4.5005
R59640 VINN.n217 VINN.n159 4.5005
R59641 VINN.n398 VINN.n159 4.5005
R59642 VINN.n216 VINN.n159 4.5005
R59643 VINN.n400 VINN.n159 4.5005
R59644 VINN.n215 VINN.n159 4.5005
R59645 VINN.n654 VINN.n159 4.5005
R59646 VINN.n656 VINN.n159 4.5005
R59647 VINN.n159 VINN.n0 4.5005
R59648 VINN.n278 VINN.n141 4.5005
R59649 VINN.n276 VINN.n141 4.5005
R59650 VINN.n280 VINN.n141 4.5005
R59651 VINN.n275 VINN.n141 4.5005
R59652 VINN.n282 VINN.n141 4.5005
R59653 VINN.n274 VINN.n141 4.5005
R59654 VINN.n284 VINN.n141 4.5005
R59655 VINN.n273 VINN.n141 4.5005
R59656 VINN.n286 VINN.n141 4.5005
R59657 VINN.n272 VINN.n141 4.5005
R59658 VINN.n288 VINN.n141 4.5005
R59659 VINN.n271 VINN.n141 4.5005
R59660 VINN.n290 VINN.n141 4.5005
R59661 VINN.n270 VINN.n141 4.5005
R59662 VINN.n292 VINN.n141 4.5005
R59663 VINN.n269 VINN.n141 4.5005
R59664 VINN.n294 VINN.n141 4.5005
R59665 VINN.n268 VINN.n141 4.5005
R59666 VINN.n296 VINN.n141 4.5005
R59667 VINN.n267 VINN.n141 4.5005
R59668 VINN.n298 VINN.n141 4.5005
R59669 VINN.n266 VINN.n141 4.5005
R59670 VINN.n300 VINN.n141 4.5005
R59671 VINN.n265 VINN.n141 4.5005
R59672 VINN.n302 VINN.n141 4.5005
R59673 VINN.n264 VINN.n141 4.5005
R59674 VINN.n304 VINN.n141 4.5005
R59675 VINN.n263 VINN.n141 4.5005
R59676 VINN.n306 VINN.n141 4.5005
R59677 VINN.n262 VINN.n141 4.5005
R59678 VINN.n308 VINN.n141 4.5005
R59679 VINN.n261 VINN.n141 4.5005
R59680 VINN.n310 VINN.n141 4.5005
R59681 VINN.n260 VINN.n141 4.5005
R59682 VINN.n312 VINN.n141 4.5005
R59683 VINN.n259 VINN.n141 4.5005
R59684 VINN.n314 VINN.n141 4.5005
R59685 VINN.n258 VINN.n141 4.5005
R59686 VINN.n316 VINN.n141 4.5005
R59687 VINN.n257 VINN.n141 4.5005
R59688 VINN.n318 VINN.n141 4.5005
R59689 VINN.n256 VINN.n141 4.5005
R59690 VINN.n320 VINN.n141 4.5005
R59691 VINN.n255 VINN.n141 4.5005
R59692 VINN.n322 VINN.n141 4.5005
R59693 VINN.n254 VINN.n141 4.5005
R59694 VINN.n324 VINN.n141 4.5005
R59695 VINN.n253 VINN.n141 4.5005
R59696 VINN.n326 VINN.n141 4.5005
R59697 VINN.n252 VINN.n141 4.5005
R59698 VINN.n328 VINN.n141 4.5005
R59699 VINN.n251 VINN.n141 4.5005
R59700 VINN.n330 VINN.n141 4.5005
R59701 VINN.n250 VINN.n141 4.5005
R59702 VINN.n332 VINN.n141 4.5005
R59703 VINN.n249 VINN.n141 4.5005
R59704 VINN.n334 VINN.n141 4.5005
R59705 VINN.n248 VINN.n141 4.5005
R59706 VINN.n336 VINN.n141 4.5005
R59707 VINN.n247 VINN.n141 4.5005
R59708 VINN.n338 VINN.n141 4.5005
R59709 VINN.n246 VINN.n141 4.5005
R59710 VINN.n340 VINN.n141 4.5005
R59711 VINN.n245 VINN.n141 4.5005
R59712 VINN.n342 VINN.n141 4.5005
R59713 VINN.n244 VINN.n141 4.5005
R59714 VINN.n344 VINN.n141 4.5005
R59715 VINN.n243 VINN.n141 4.5005
R59716 VINN.n346 VINN.n141 4.5005
R59717 VINN.n242 VINN.n141 4.5005
R59718 VINN.n348 VINN.n141 4.5005
R59719 VINN.n241 VINN.n141 4.5005
R59720 VINN.n350 VINN.n141 4.5005
R59721 VINN.n240 VINN.n141 4.5005
R59722 VINN.n352 VINN.n141 4.5005
R59723 VINN.n239 VINN.n141 4.5005
R59724 VINN.n354 VINN.n141 4.5005
R59725 VINN.n238 VINN.n141 4.5005
R59726 VINN.n356 VINN.n141 4.5005
R59727 VINN.n237 VINN.n141 4.5005
R59728 VINN.n358 VINN.n141 4.5005
R59729 VINN.n236 VINN.n141 4.5005
R59730 VINN.n360 VINN.n141 4.5005
R59731 VINN.n235 VINN.n141 4.5005
R59732 VINN.n362 VINN.n141 4.5005
R59733 VINN.n234 VINN.n141 4.5005
R59734 VINN.n364 VINN.n141 4.5005
R59735 VINN.n233 VINN.n141 4.5005
R59736 VINN.n366 VINN.n141 4.5005
R59737 VINN.n232 VINN.n141 4.5005
R59738 VINN.n368 VINN.n141 4.5005
R59739 VINN.n231 VINN.n141 4.5005
R59740 VINN.n370 VINN.n141 4.5005
R59741 VINN.n230 VINN.n141 4.5005
R59742 VINN.n372 VINN.n141 4.5005
R59743 VINN.n229 VINN.n141 4.5005
R59744 VINN.n374 VINN.n141 4.5005
R59745 VINN.n228 VINN.n141 4.5005
R59746 VINN.n376 VINN.n141 4.5005
R59747 VINN.n227 VINN.n141 4.5005
R59748 VINN.n378 VINN.n141 4.5005
R59749 VINN.n226 VINN.n141 4.5005
R59750 VINN.n380 VINN.n141 4.5005
R59751 VINN.n225 VINN.n141 4.5005
R59752 VINN.n382 VINN.n141 4.5005
R59753 VINN.n224 VINN.n141 4.5005
R59754 VINN.n384 VINN.n141 4.5005
R59755 VINN.n223 VINN.n141 4.5005
R59756 VINN.n386 VINN.n141 4.5005
R59757 VINN.n222 VINN.n141 4.5005
R59758 VINN.n388 VINN.n141 4.5005
R59759 VINN.n221 VINN.n141 4.5005
R59760 VINN.n390 VINN.n141 4.5005
R59761 VINN.n220 VINN.n141 4.5005
R59762 VINN.n392 VINN.n141 4.5005
R59763 VINN.n219 VINN.n141 4.5005
R59764 VINN.n394 VINN.n141 4.5005
R59765 VINN.n218 VINN.n141 4.5005
R59766 VINN.n396 VINN.n141 4.5005
R59767 VINN.n217 VINN.n141 4.5005
R59768 VINN.n398 VINN.n141 4.5005
R59769 VINN.n216 VINN.n141 4.5005
R59770 VINN.n400 VINN.n141 4.5005
R59771 VINN.n215 VINN.n141 4.5005
R59772 VINN.n654 VINN.n141 4.5005
R59773 VINN.n656 VINN.n141 4.5005
R59774 VINN.n141 VINN.n0 4.5005
R59775 VINN.n278 VINN.n160 4.5005
R59776 VINN.n276 VINN.n160 4.5005
R59777 VINN.n280 VINN.n160 4.5005
R59778 VINN.n275 VINN.n160 4.5005
R59779 VINN.n282 VINN.n160 4.5005
R59780 VINN.n274 VINN.n160 4.5005
R59781 VINN.n284 VINN.n160 4.5005
R59782 VINN.n273 VINN.n160 4.5005
R59783 VINN.n286 VINN.n160 4.5005
R59784 VINN.n272 VINN.n160 4.5005
R59785 VINN.n288 VINN.n160 4.5005
R59786 VINN.n271 VINN.n160 4.5005
R59787 VINN.n290 VINN.n160 4.5005
R59788 VINN.n270 VINN.n160 4.5005
R59789 VINN.n292 VINN.n160 4.5005
R59790 VINN.n269 VINN.n160 4.5005
R59791 VINN.n294 VINN.n160 4.5005
R59792 VINN.n268 VINN.n160 4.5005
R59793 VINN.n296 VINN.n160 4.5005
R59794 VINN.n267 VINN.n160 4.5005
R59795 VINN.n298 VINN.n160 4.5005
R59796 VINN.n266 VINN.n160 4.5005
R59797 VINN.n300 VINN.n160 4.5005
R59798 VINN.n265 VINN.n160 4.5005
R59799 VINN.n302 VINN.n160 4.5005
R59800 VINN.n264 VINN.n160 4.5005
R59801 VINN.n304 VINN.n160 4.5005
R59802 VINN.n263 VINN.n160 4.5005
R59803 VINN.n306 VINN.n160 4.5005
R59804 VINN.n262 VINN.n160 4.5005
R59805 VINN.n308 VINN.n160 4.5005
R59806 VINN.n261 VINN.n160 4.5005
R59807 VINN.n310 VINN.n160 4.5005
R59808 VINN.n260 VINN.n160 4.5005
R59809 VINN.n312 VINN.n160 4.5005
R59810 VINN.n259 VINN.n160 4.5005
R59811 VINN.n314 VINN.n160 4.5005
R59812 VINN.n258 VINN.n160 4.5005
R59813 VINN.n316 VINN.n160 4.5005
R59814 VINN.n257 VINN.n160 4.5005
R59815 VINN.n318 VINN.n160 4.5005
R59816 VINN.n256 VINN.n160 4.5005
R59817 VINN.n320 VINN.n160 4.5005
R59818 VINN.n255 VINN.n160 4.5005
R59819 VINN.n322 VINN.n160 4.5005
R59820 VINN.n254 VINN.n160 4.5005
R59821 VINN.n324 VINN.n160 4.5005
R59822 VINN.n253 VINN.n160 4.5005
R59823 VINN.n326 VINN.n160 4.5005
R59824 VINN.n252 VINN.n160 4.5005
R59825 VINN.n328 VINN.n160 4.5005
R59826 VINN.n251 VINN.n160 4.5005
R59827 VINN.n330 VINN.n160 4.5005
R59828 VINN.n250 VINN.n160 4.5005
R59829 VINN.n332 VINN.n160 4.5005
R59830 VINN.n249 VINN.n160 4.5005
R59831 VINN.n334 VINN.n160 4.5005
R59832 VINN.n248 VINN.n160 4.5005
R59833 VINN.n336 VINN.n160 4.5005
R59834 VINN.n247 VINN.n160 4.5005
R59835 VINN.n338 VINN.n160 4.5005
R59836 VINN.n246 VINN.n160 4.5005
R59837 VINN.n340 VINN.n160 4.5005
R59838 VINN.n245 VINN.n160 4.5005
R59839 VINN.n342 VINN.n160 4.5005
R59840 VINN.n244 VINN.n160 4.5005
R59841 VINN.n344 VINN.n160 4.5005
R59842 VINN.n243 VINN.n160 4.5005
R59843 VINN.n346 VINN.n160 4.5005
R59844 VINN.n242 VINN.n160 4.5005
R59845 VINN.n348 VINN.n160 4.5005
R59846 VINN.n241 VINN.n160 4.5005
R59847 VINN.n350 VINN.n160 4.5005
R59848 VINN.n240 VINN.n160 4.5005
R59849 VINN.n352 VINN.n160 4.5005
R59850 VINN.n239 VINN.n160 4.5005
R59851 VINN.n354 VINN.n160 4.5005
R59852 VINN.n238 VINN.n160 4.5005
R59853 VINN.n356 VINN.n160 4.5005
R59854 VINN.n237 VINN.n160 4.5005
R59855 VINN.n358 VINN.n160 4.5005
R59856 VINN.n236 VINN.n160 4.5005
R59857 VINN.n360 VINN.n160 4.5005
R59858 VINN.n235 VINN.n160 4.5005
R59859 VINN.n362 VINN.n160 4.5005
R59860 VINN.n234 VINN.n160 4.5005
R59861 VINN.n364 VINN.n160 4.5005
R59862 VINN.n233 VINN.n160 4.5005
R59863 VINN.n366 VINN.n160 4.5005
R59864 VINN.n232 VINN.n160 4.5005
R59865 VINN.n368 VINN.n160 4.5005
R59866 VINN.n231 VINN.n160 4.5005
R59867 VINN.n370 VINN.n160 4.5005
R59868 VINN.n230 VINN.n160 4.5005
R59869 VINN.n372 VINN.n160 4.5005
R59870 VINN.n229 VINN.n160 4.5005
R59871 VINN.n374 VINN.n160 4.5005
R59872 VINN.n228 VINN.n160 4.5005
R59873 VINN.n376 VINN.n160 4.5005
R59874 VINN.n227 VINN.n160 4.5005
R59875 VINN.n378 VINN.n160 4.5005
R59876 VINN.n226 VINN.n160 4.5005
R59877 VINN.n380 VINN.n160 4.5005
R59878 VINN.n225 VINN.n160 4.5005
R59879 VINN.n382 VINN.n160 4.5005
R59880 VINN.n224 VINN.n160 4.5005
R59881 VINN.n384 VINN.n160 4.5005
R59882 VINN.n223 VINN.n160 4.5005
R59883 VINN.n386 VINN.n160 4.5005
R59884 VINN.n222 VINN.n160 4.5005
R59885 VINN.n388 VINN.n160 4.5005
R59886 VINN.n221 VINN.n160 4.5005
R59887 VINN.n390 VINN.n160 4.5005
R59888 VINN.n220 VINN.n160 4.5005
R59889 VINN.n392 VINN.n160 4.5005
R59890 VINN.n219 VINN.n160 4.5005
R59891 VINN.n394 VINN.n160 4.5005
R59892 VINN.n218 VINN.n160 4.5005
R59893 VINN.n396 VINN.n160 4.5005
R59894 VINN.n217 VINN.n160 4.5005
R59895 VINN.n398 VINN.n160 4.5005
R59896 VINN.n216 VINN.n160 4.5005
R59897 VINN.n400 VINN.n160 4.5005
R59898 VINN.n215 VINN.n160 4.5005
R59899 VINN.n654 VINN.n160 4.5005
R59900 VINN.n656 VINN.n160 4.5005
R59901 VINN.n160 VINN.n0 4.5005
R59902 VINN.n278 VINN.n140 4.5005
R59903 VINN.n276 VINN.n140 4.5005
R59904 VINN.n280 VINN.n140 4.5005
R59905 VINN.n275 VINN.n140 4.5005
R59906 VINN.n282 VINN.n140 4.5005
R59907 VINN.n274 VINN.n140 4.5005
R59908 VINN.n284 VINN.n140 4.5005
R59909 VINN.n273 VINN.n140 4.5005
R59910 VINN.n286 VINN.n140 4.5005
R59911 VINN.n272 VINN.n140 4.5005
R59912 VINN.n288 VINN.n140 4.5005
R59913 VINN.n271 VINN.n140 4.5005
R59914 VINN.n290 VINN.n140 4.5005
R59915 VINN.n270 VINN.n140 4.5005
R59916 VINN.n292 VINN.n140 4.5005
R59917 VINN.n269 VINN.n140 4.5005
R59918 VINN.n294 VINN.n140 4.5005
R59919 VINN.n268 VINN.n140 4.5005
R59920 VINN.n296 VINN.n140 4.5005
R59921 VINN.n267 VINN.n140 4.5005
R59922 VINN.n298 VINN.n140 4.5005
R59923 VINN.n266 VINN.n140 4.5005
R59924 VINN.n300 VINN.n140 4.5005
R59925 VINN.n265 VINN.n140 4.5005
R59926 VINN.n302 VINN.n140 4.5005
R59927 VINN.n264 VINN.n140 4.5005
R59928 VINN.n304 VINN.n140 4.5005
R59929 VINN.n263 VINN.n140 4.5005
R59930 VINN.n306 VINN.n140 4.5005
R59931 VINN.n262 VINN.n140 4.5005
R59932 VINN.n308 VINN.n140 4.5005
R59933 VINN.n261 VINN.n140 4.5005
R59934 VINN.n310 VINN.n140 4.5005
R59935 VINN.n260 VINN.n140 4.5005
R59936 VINN.n312 VINN.n140 4.5005
R59937 VINN.n259 VINN.n140 4.5005
R59938 VINN.n314 VINN.n140 4.5005
R59939 VINN.n258 VINN.n140 4.5005
R59940 VINN.n316 VINN.n140 4.5005
R59941 VINN.n257 VINN.n140 4.5005
R59942 VINN.n318 VINN.n140 4.5005
R59943 VINN.n256 VINN.n140 4.5005
R59944 VINN.n320 VINN.n140 4.5005
R59945 VINN.n255 VINN.n140 4.5005
R59946 VINN.n322 VINN.n140 4.5005
R59947 VINN.n254 VINN.n140 4.5005
R59948 VINN.n324 VINN.n140 4.5005
R59949 VINN.n253 VINN.n140 4.5005
R59950 VINN.n326 VINN.n140 4.5005
R59951 VINN.n252 VINN.n140 4.5005
R59952 VINN.n328 VINN.n140 4.5005
R59953 VINN.n251 VINN.n140 4.5005
R59954 VINN.n330 VINN.n140 4.5005
R59955 VINN.n250 VINN.n140 4.5005
R59956 VINN.n332 VINN.n140 4.5005
R59957 VINN.n249 VINN.n140 4.5005
R59958 VINN.n334 VINN.n140 4.5005
R59959 VINN.n248 VINN.n140 4.5005
R59960 VINN.n336 VINN.n140 4.5005
R59961 VINN.n247 VINN.n140 4.5005
R59962 VINN.n338 VINN.n140 4.5005
R59963 VINN.n246 VINN.n140 4.5005
R59964 VINN.n340 VINN.n140 4.5005
R59965 VINN.n245 VINN.n140 4.5005
R59966 VINN.n342 VINN.n140 4.5005
R59967 VINN.n244 VINN.n140 4.5005
R59968 VINN.n344 VINN.n140 4.5005
R59969 VINN.n243 VINN.n140 4.5005
R59970 VINN.n346 VINN.n140 4.5005
R59971 VINN.n242 VINN.n140 4.5005
R59972 VINN.n348 VINN.n140 4.5005
R59973 VINN.n241 VINN.n140 4.5005
R59974 VINN.n350 VINN.n140 4.5005
R59975 VINN.n240 VINN.n140 4.5005
R59976 VINN.n352 VINN.n140 4.5005
R59977 VINN.n239 VINN.n140 4.5005
R59978 VINN.n354 VINN.n140 4.5005
R59979 VINN.n238 VINN.n140 4.5005
R59980 VINN.n356 VINN.n140 4.5005
R59981 VINN.n237 VINN.n140 4.5005
R59982 VINN.n358 VINN.n140 4.5005
R59983 VINN.n236 VINN.n140 4.5005
R59984 VINN.n360 VINN.n140 4.5005
R59985 VINN.n235 VINN.n140 4.5005
R59986 VINN.n362 VINN.n140 4.5005
R59987 VINN.n234 VINN.n140 4.5005
R59988 VINN.n364 VINN.n140 4.5005
R59989 VINN.n233 VINN.n140 4.5005
R59990 VINN.n366 VINN.n140 4.5005
R59991 VINN.n232 VINN.n140 4.5005
R59992 VINN.n368 VINN.n140 4.5005
R59993 VINN.n231 VINN.n140 4.5005
R59994 VINN.n370 VINN.n140 4.5005
R59995 VINN.n230 VINN.n140 4.5005
R59996 VINN.n372 VINN.n140 4.5005
R59997 VINN.n229 VINN.n140 4.5005
R59998 VINN.n374 VINN.n140 4.5005
R59999 VINN.n228 VINN.n140 4.5005
R60000 VINN.n376 VINN.n140 4.5005
R60001 VINN.n227 VINN.n140 4.5005
R60002 VINN.n378 VINN.n140 4.5005
R60003 VINN.n226 VINN.n140 4.5005
R60004 VINN.n380 VINN.n140 4.5005
R60005 VINN.n225 VINN.n140 4.5005
R60006 VINN.n382 VINN.n140 4.5005
R60007 VINN.n224 VINN.n140 4.5005
R60008 VINN.n384 VINN.n140 4.5005
R60009 VINN.n223 VINN.n140 4.5005
R60010 VINN.n386 VINN.n140 4.5005
R60011 VINN.n222 VINN.n140 4.5005
R60012 VINN.n388 VINN.n140 4.5005
R60013 VINN.n221 VINN.n140 4.5005
R60014 VINN.n390 VINN.n140 4.5005
R60015 VINN.n220 VINN.n140 4.5005
R60016 VINN.n392 VINN.n140 4.5005
R60017 VINN.n219 VINN.n140 4.5005
R60018 VINN.n394 VINN.n140 4.5005
R60019 VINN.n218 VINN.n140 4.5005
R60020 VINN.n396 VINN.n140 4.5005
R60021 VINN.n217 VINN.n140 4.5005
R60022 VINN.n398 VINN.n140 4.5005
R60023 VINN.n216 VINN.n140 4.5005
R60024 VINN.n400 VINN.n140 4.5005
R60025 VINN.n215 VINN.n140 4.5005
R60026 VINN.n654 VINN.n140 4.5005
R60027 VINN.n656 VINN.n140 4.5005
R60028 VINN.n140 VINN.n0 4.5005
R60029 VINN.n278 VINN.n161 4.5005
R60030 VINN.n276 VINN.n161 4.5005
R60031 VINN.n280 VINN.n161 4.5005
R60032 VINN.n275 VINN.n161 4.5005
R60033 VINN.n282 VINN.n161 4.5005
R60034 VINN.n274 VINN.n161 4.5005
R60035 VINN.n284 VINN.n161 4.5005
R60036 VINN.n273 VINN.n161 4.5005
R60037 VINN.n286 VINN.n161 4.5005
R60038 VINN.n272 VINN.n161 4.5005
R60039 VINN.n288 VINN.n161 4.5005
R60040 VINN.n271 VINN.n161 4.5005
R60041 VINN.n290 VINN.n161 4.5005
R60042 VINN.n270 VINN.n161 4.5005
R60043 VINN.n292 VINN.n161 4.5005
R60044 VINN.n269 VINN.n161 4.5005
R60045 VINN.n294 VINN.n161 4.5005
R60046 VINN.n268 VINN.n161 4.5005
R60047 VINN.n296 VINN.n161 4.5005
R60048 VINN.n267 VINN.n161 4.5005
R60049 VINN.n298 VINN.n161 4.5005
R60050 VINN.n266 VINN.n161 4.5005
R60051 VINN.n300 VINN.n161 4.5005
R60052 VINN.n265 VINN.n161 4.5005
R60053 VINN.n302 VINN.n161 4.5005
R60054 VINN.n264 VINN.n161 4.5005
R60055 VINN.n304 VINN.n161 4.5005
R60056 VINN.n263 VINN.n161 4.5005
R60057 VINN.n306 VINN.n161 4.5005
R60058 VINN.n262 VINN.n161 4.5005
R60059 VINN.n308 VINN.n161 4.5005
R60060 VINN.n261 VINN.n161 4.5005
R60061 VINN.n310 VINN.n161 4.5005
R60062 VINN.n260 VINN.n161 4.5005
R60063 VINN.n312 VINN.n161 4.5005
R60064 VINN.n259 VINN.n161 4.5005
R60065 VINN.n314 VINN.n161 4.5005
R60066 VINN.n258 VINN.n161 4.5005
R60067 VINN.n316 VINN.n161 4.5005
R60068 VINN.n257 VINN.n161 4.5005
R60069 VINN.n318 VINN.n161 4.5005
R60070 VINN.n256 VINN.n161 4.5005
R60071 VINN.n320 VINN.n161 4.5005
R60072 VINN.n255 VINN.n161 4.5005
R60073 VINN.n322 VINN.n161 4.5005
R60074 VINN.n254 VINN.n161 4.5005
R60075 VINN.n324 VINN.n161 4.5005
R60076 VINN.n253 VINN.n161 4.5005
R60077 VINN.n326 VINN.n161 4.5005
R60078 VINN.n252 VINN.n161 4.5005
R60079 VINN.n328 VINN.n161 4.5005
R60080 VINN.n251 VINN.n161 4.5005
R60081 VINN.n330 VINN.n161 4.5005
R60082 VINN.n250 VINN.n161 4.5005
R60083 VINN.n332 VINN.n161 4.5005
R60084 VINN.n249 VINN.n161 4.5005
R60085 VINN.n334 VINN.n161 4.5005
R60086 VINN.n248 VINN.n161 4.5005
R60087 VINN.n336 VINN.n161 4.5005
R60088 VINN.n247 VINN.n161 4.5005
R60089 VINN.n338 VINN.n161 4.5005
R60090 VINN.n246 VINN.n161 4.5005
R60091 VINN.n340 VINN.n161 4.5005
R60092 VINN.n245 VINN.n161 4.5005
R60093 VINN.n342 VINN.n161 4.5005
R60094 VINN.n244 VINN.n161 4.5005
R60095 VINN.n344 VINN.n161 4.5005
R60096 VINN.n243 VINN.n161 4.5005
R60097 VINN.n346 VINN.n161 4.5005
R60098 VINN.n242 VINN.n161 4.5005
R60099 VINN.n348 VINN.n161 4.5005
R60100 VINN.n241 VINN.n161 4.5005
R60101 VINN.n350 VINN.n161 4.5005
R60102 VINN.n240 VINN.n161 4.5005
R60103 VINN.n352 VINN.n161 4.5005
R60104 VINN.n239 VINN.n161 4.5005
R60105 VINN.n354 VINN.n161 4.5005
R60106 VINN.n238 VINN.n161 4.5005
R60107 VINN.n356 VINN.n161 4.5005
R60108 VINN.n237 VINN.n161 4.5005
R60109 VINN.n358 VINN.n161 4.5005
R60110 VINN.n236 VINN.n161 4.5005
R60111 VINN.n360 VINN.n161 4.5005
R60112 VINN.n235 VINN.n161 4.5005
R60113 VINN.n362 VINN.n161 4.5005
R60114 VINN.n234 VINN.n161 4.5005
R60115 VINN.n364 VINN.n161 4.5005
R60116 VINN.n233 VINN.n161 4.5005
R60117 VINN.n366 VINN.n161 4.5005
R60118 VINN.n232 VINN.n161 4.5005
R60119 VINN.n368 VINN.n161 4.5005
R60120 VINN.n231 VINN.n161 4.5005
R60121 VINN.n370 VINN.n161 4.5005
R60122 VINN.n230 VINN.n161 4.5005
R60123 VINN.n372 VINN.n161 4.5005
R60124 VINN.n229 VINN.n161 4.5005
R60125 VINN.n374 VINN.n161 4.5005
R60126 VINN.n228 VINN.n161 4.5005
R60127 VINN.n376 VINN.n161 4.5005
R60128 VINN.n227 VINN.n161 4.5005
R60129 VINN.n378 VINN.n161 4.5005
R60130 VINN.n226 VINN.n161 4.5005
R60131 VINN.n380 VINN.n161 4.5005
R60132 VINN.n225 VINN.n161 4.5005
R60133 VINN.n382 VINN.n161 4.5005
R60134 VINN.n224 VINN.n161 4.5005
R60135 VINN.n384 VINN.n161 4.5005
R60136 VINN.n223 VINN.n161 4.5005
R60137 VINN.n386 VINN.n161 4.5005
R60138 VINN.n222 VINN.n161 4.5005
R60139 VINN.n388 VINN.n161 4.5005
R60140 VINN.n221 VINN.n161 4.5005
R60141 VINN.n390 VINN.n161 4.5005
R60142 VINN.n220 VINN.n161 4.5005
R60143 VINN.n392 VINN.n161 4.5005
R60144 VINN.n219 VINN.n161 4.5005
R60145 VINN.n394 VINN.n161 4.5005
R60146 VINN.n218 VINN.n161 4.5005
R60147 VINN.n396 VINN.n161 4.5005
R60148 VINN.n217 VINN.n161 4.5005
R60149 VINN.n398 VINN.n161 4.5005
R60150 VINN.n216 VINN.n161 4.5005
R60151 VINN.n400 VINN.n161 4.5005
R60152 VINN.n215 VINN.n161 4.5005
R60153 VINN.n654 VINN.n161 4.5005
R60154 VINN.n656 VINN.n161 4.5005
R60155 VINN.n161 VINN.n0 4.5005
R60156 VINN.n278 VINN.n139 4.5005
R60157 VINN.n276 VINN.n139 4.5005
R60158 VINN.n280 VINN.n139 4.5005
R60159 VINN.n275 VINN.n139 4.5005
R60160 VINN.n282 VINN.n139 4.5005
R60161 VINN.n274 VINN.n139 4.5005
R60162 VINN.n284 VINN.n139 4.5005
R60163 VINN.n273 VINN.n139 4.5005
R60164 VINN.n286 VINN.n139 4.5005
R60165 VINN.n272 VINN.n139 4.5005
R60166 VINN.n288 VINN.n139 4.5005
R60167 VINN.n271 VINN.n139 4.5005
R60168 VINN.n290 VINN.n139 4.5005
R60169 VINN.n270 VINN.n139 4.5005
R60170 VINN.n292 VINN.n139 4.5005
R60171 VINN.n269 VINN.n139 4.5005
R60172 VINN.n294 VINN.n139 4.5005
R60173 VINN.n268 VINN.n139 4.5005
R60174 VINN.n296 VINN.n139 4.5005
R60175 VINN.n267 VINN.n139 4.5005
R60176 VINN.n298 VINN.n139 4.5005
R60177 VINN.n266 VINN.n139 4.5005
R60178 VINN.n300 VINN.n139 4.5005
R60179 VINN.n265 VINN.n139 4.5005
R60180 VINN.n302 VINN.n139 4.5005
R60181 VINN.n264 VINN.n139 4.5005
R60182 VINN.n304 VINN.n139 4.5005
R60183 VINN.n263 VINN.n139 4.5005
R60184 VINN.n306 VINN.n139 4.5005
R60185 VINN.n262 VINN.n139 4.5005
R60186 VINN.n308 VINN.n139 4.5005
R60187 VINN.n261 VINN.n139 4.5005
R60188 VINN.n310 VINN.n139 4.5005
R60189 VINN.n260 VINN.n139 4.5005
R60190 VINN.n312 VINN.n139 4.5005
R60191 VINN.n259 VINN.n139 4.5005
R60192 VINN.n314 VINN.n139 4.5005
R60193 VINN.n258 VINN.n139 4.5005
R60194 VINN.n316 VINN.n139 4.5005
R60195 VINN.n257 VINN.n139 4.5005
R60196 VINN.n318 VINN.n139 4.5005
R60197 VINN.n256 VINN.n139 4.5005
R60198 VINN.n320 VINN.n139 4.5005
R60199 VINN.n255 VINN.n139 4.5005
R60200 VINN.n322 VINN.n139 4.5005
R60201 VINN.n254 VINN.n139 4.5005
R60202 VINN.n324 VINN.n139 4.5005
R60203 VINN.n253 VINN.n139 4.5005
R60204 VINN.n326 VINN.n139 4.5005
R60205 VINN.n252 VINN.n139 4.5005
R60206 VINN.n328 VINN.n139 4.5005
R60207 VINN.n251 VINN.n139 4.5005
R60208 VINN.n330 VINN.n139 4.5005
R60209 VINN.n250 VINN.n139 4.5005
R60210 VINN.n332 VINN.n139 4.5005
R60211 VINN.n249 VINN.n139 4.5005
R60212 VINN.n334 VINN.n139 4.5005
R60213 VINN.n248 VINN.n139 4.5005
R60214 VINN.n336 VINN.n139 4.5005
R60215 VINN.n247 VINN.n139 4.5005
R60216 VINN.n338 VINN.n139 4.5005
R60217 VINN.n246 VINN.n139 4.5005
R60218 VINN.n340 VINN.n139 4.5005
R60219 VINN.n245 VINN.n139 4.5005
R60220 VINN.n342 VINN.n139 4.5005
R60221 VINN.n244 VINN.n139 4.5005
R60222 VINN.n344 VINN.n139 4.5005
R60223 VINN.n243 VINN.n139 4.5005
R60224 VINN.n346 VINN.n139 4.5005
R60225 VINN.n242 VINN.n139 4.5005
R60226 VINN.n348 VINN.n139 4.5005
R60227 VINN.n241 VINN.n139 4.5005
R60228 VINN.n350 VINN.n139 4.5005
R60229 VINN.n240 VINN.n139 4.5005
R60230 VINN.n352 VINN.n139 4.5005
R60231 VINN.n239 VINN.n139 4.5005
R60232 VINN.n354 VINN.n139 4.5005
R60233 VINN.n238 VINN.n139 4.5005
R60234 VINN.n356 VINN.n139 4.5005
R60235 VINN.n237 VINN.n139 4.5005
R60236 VINN.n358 VINN.n139 4.5005
R60237 VINN.n236 VINN.n139 4.5005
R60238 VINN.n360 VINN.n139 4.5005
R60239 VINN.n235 VINN.n139 4.5005
R60240 VINN.n362 VINN.n139 4.5005
R60241 VINN.n234 VINN.n139 4.5005
R60242 VINN.n364 VINN.n139 4.5005
R60243 VINN.n233 VINN.n139 4.5005
R60244 VINN.n366 VINN.n139 4.5005
R60245 VINN.n232 VINN.n139 4.5005
R60246 VINN.n368 VINN.n139 4.5005
R60247 VINN.n231 VINN.n139 4.5005
R60248 VINN.n370 VINN.n139 4.5005
R60249 VINN.n230 VINN.n139 4.5005
R60250 VINN.n372 VINN.n139 4.5005
R60251 VINN.n229 VINN.n139 4.5005
R60252 VINN.n374 VINN.n139 4.5005
R60253 VINN.n228 VINN.n139 4.5005
R60254 VINN.n376 VINN.n139 4.5005
R60255 VINN.n227 VINN.n139 4.5005
R60256 VINN.n378 VINN.n139 4.5005
R60257 VINN.n226 VINN.n139 4.5005
R60258 VINN.n380 VINN.n139 4.5005
R60259 VINN.n225 VINN.n139 4.5005
R60260 VINN.n382 VINN.n139 4.5005
R60261 VINN.n224 VINN.n139 4.5005
R60262 VINN.n384 VINN.n139 4.5005
R60263 VINN.n223 VINN.n139 4.5005
R60264 VINN.n386 VINN.n139 4.5005
R60265 VINN.n222 VINN.n139 4.5005
R60266 VINN.n388 VINN.n139 4.5005
R60267 VINN.n221 VINN.n139 4.5005
R60268 VINN.n390 VINN.n139 4.5005
R60269 VINN.n220 VINN.n139 4.5005
R60270 VINN.n392 VINN.n139 4.5005
R60271 VINN.n219 VINN.n139 4.5005
R60272 VINN.n394 VINN.n139 4.5005
R60273 VINN.n218 VINN.n139 4.5005
R60274 VINN.n396 VINN.n139 4.5005
R60275 VINN.n217 VINN.n139 4.5005
R60276 VINN.n398 VINN.n139 4.5005
R60277 VINN.n216 VINN.n139 4.5005
R60278 VINN.n400 VINN.n139 4.5005
R60279 VINN.n215 VINN.n139 4.5005
R60280 VINN.n654 VINN.n139 4.5005
R60281 VINN.n656 VINN.n139 4.5005
R60282 VINN.n139 VINN.n0 4.5005
R60283 VINN.n278 VINN.n162 4.5005
R60284 VINN.n276 VINN.n162 4.5005
R60285 VINN.n280 VINN.n162 4.5005
R60286 VINN.n275 VINN.n162 4.5005
R60287 VINN.n282 VINN.n162 4.5005
R60288 VINN.n274 VINN.n162 4.5005
R60289 VINN.n284 VINN.n162 4.5005
R60290 VINN.n273 VINN.n162 4.5005
R60291 VINN.n286 VINN.n162 4.5005
R60292 VINN.n272 VINN.n162 4.5005
R60293 VINN.n288 VINN.n162 4.5005
R60294 VINN.n271 VINN.n162 4.5005
R60295 VINN.n290 VINN.n162 4.5005
R60296 VINN.n270 VINN.n162 4.5005
R60297 VINN.n292 VINN.n162 4.5005
R60298 VINN.n269 VINN.n162 4.5005
R60299 VINN.n294 VINN.n162 4.5005
R60300 VINN.n268 VINN.n162 4.5005
R60301 VINN.n296 VINN.n162 4.5005
R60302 VINN.n267 VINN.n162 4.5005
R60303 VINN.n298 VINN.n162 4.5005
R60304 VINN.n266 VINN.n162 4.5005
R60305 VINN.n300 VINN.n162 4.5005
R60306 VINN.n265 VINN.n162 4.5005
R60307 VINN.n302 VINN.n162 4.5005
R60308 VINN.n264 VINN.n162 4.5005
R60309 VINN.n304 VINN.n162 4.5005
R60310 VINN.n263 VINN.n162 4.5005
R60311 VINN.n306 VINN.n162 4.5005
R60312 VINN.n262 VINN.n162 4.5005
R60313 VINN.n308 VINN.n162 4.5005
R60314 VINN.n261 VINN.n162 4.5005
R60315 VINN.n310 VINN.n162 4.5005
R60316 VINN.n260 VINN.n162 4.5005
R60317 VINN.n312 VINN.n162 4.5005
R60318 VINN.n259 VINN.n162 4.5005
R60319 VINN.n314 VINN.n162 4.5005
R60320 VINN.n258 VINN.n162 4.5005
R60321 VINN.n316 VINN.n162 4.5005
R60322 VINN.n257 VINN.n162 4.5005
R60323 VINN.n318 VINN.n162 4.5005
R60324 VINN.n256 VINN.n162 4.5005
R60325 VINN.n320 VINN.n162 4.5005
R60326 VINN.n255 VINN.n162 4.5005
R60327 VINN.n322 VINN.n162 4.5005
R60328 VINN.n254 VINN.n162 4.5005
R60329 VINN.n324 VINN.n162 4.5005
R60330 VINN.n253 VINN.n162 4.5005
R60331 VINN.n326 VINN.n162 4.5005
R60332 VINN.n252 VINN.n162 4.5005
R60333 VINN.n328 VINN.n162 4.5005
R60334 VINN.n251 VINN.n162 4.5005
R60335 VINN.n330 VINN.n162 4.5005
R60336 VINN.n250 VINN.n162 4.5005
R60337 VINN.n332 VINN.n162 4.5005
R60338 VINN.n249 VINN.n162 4.5005
R60339 VINN.n334 VINN.n162 4.5005
R60340 VINN.n248 VINN.n162 4.5005
R60341 VINN.n336 VINN.n162 4.5005
R60342 VINN.n247 VINN.n162 4.5005
R60343 VINN.n338 VINN.n162 4.5005
R60344 VINN.n246 VINN.n162 4.5005
R60345 VINN.n340 VINN.n162 4.5005
R60346 VINN.n245 VINN.n162 4.5005
R60347 VINN.n342 VINN.n162 4.5005
R60348 VINN.n244 VINN.n162 4.5005
R60349 VINN.n344 VINN.n162 4.5005
R60350 VINN.n243 VINN.n162 4.5005
R60351 VINN.n346 VINN.n162 4.5005
R60352 VINN.n242 VINN.n162 4.5005
R60353 VINN.n348 VINN.n162 4.5005
R60354 VINN.n241 VINN.n162 4.5005
R60355 VINN.n350 VINN.n162 4.5005
R60356 VINN.n240 VINN.n162 4.5005
R60357 VINN.n352 VINN.n162 4.5005
R60358 VINN.n239 VINN.n162 4.5005
R60359 VINN.n354 VINN.n162 4.5005
R60360 VINN.n238 VINN.n162 4.5005
R60361 VINN.n356 VINN.n162 4.5005
R60362 VINN.n237 VINN.n162 4.5005
R60363 VINN.n358 VINN.n162 4.5005
R60364 VINN.n236 VINN.n162 4.5005
R60365 VINN.n360 VINN.n162 4.5005
R60366 VINN.n235 VINN.n162 4.5005
R60367 VINN.n362 VINN.n162 4.5005
R60368 VINN.n234 VINN.n162 4.5005
R60369 VINN.n364 VINN.n162 4.5005
R60370 VINN.n233 VINN.n162 4.5005
R60371 VINN.n366 VINN.n162 4.5005
R60372 VINN.n232 VINN.n162 4.5005
R60373 VINN.n368 VINN.n162 4.5005
R60374 VINN.n231 VINN.n162 4.5005
R60375 VINN.n370 VINN.n162 4.5005
R60376 VINN.n230 VINN.n162 4.5005
R60377 VINN.n372 VINN.n162 4.5005
R60378 VINN.n229 VINN.n162 4.5005
R60379 VINN.n374 VINN.n162 4.5005
R60380 VINN.n228 VINN.n162 4.5005
R60381 VINN.n376 VINN.n162 4.5005
R60382 VINN.n227 VINN.n162 4.5005
R60383 VINN.n378 VINN.n162 4.5005
R60384 VINN.n226 VINN.n162 4.5005
R60385 VINN.n380 VINN.n162 4.5005
R60386 VINN.n225 VINN.n162 4.5005
R60387 VINN.n382 VINN.n162 4.5005
R60388 VINN.n224 VINN.n162 4.5005
R60389 VINN.n384 VINN.n162 4.5005
R60390 VINN.n223 VINN.n162 4.5005
R60391 VINN.n386 VINN.n162 4.5005
R60392 VINN.n222 VINN.n162 4.5005
R60393 VINN.n388 VINN.n162 4.5005
R60394 VINN.n221 VINN.n162 4.5005
R60395 VINN.n390 VINN.n162 4.5005
R60396 VINN.n220 VINN.n162 4.5005
R60397 VINN.n392 VINN.n162 4.5005
R60398 VINN.n219 VINN.n162 4.5005
R60399 VINN.n394 VINN.n162 4.5005
R60400 VINN.n218 VINN.n162 4.5005
R60401 VINN.n396 VINN.n162 4.5005
R60402 VINN.n217 VINN.n162 4.5005
R60403 VINN.n398 VINN.n162 4.5005
R60404 VINN.n216 VINN.n162 4.5005
R60405 VINN.n400 VINN.n162 4.5005
R60406 VINN.n215 VINN.n162 4.5005
R60407 VINN.n654 VINN.n162 4.5005
R60408 VINN.n656 VINN.n162 4.5005
R60409 VINN.n162 VINN.n0 4.5005
R60410 VINN.n278 VINN.n138 4.5005
R60411 VINN.n276 VINN.n138 4.5005
R60412 VINN.n280 VINN.n138 4.5005
R60413 VINN.n275 VINN.n138 4.5005
R60414 VINN.n282 VINN.n138 4.5005
R60415 VINN.n274 VINN.n138 4.5005
R60416 VINN.n284 VINN.n138 4.5005
R60417 VINN.n273 VINN.n138 4.5005
R60418 VINN.n286 VINN.n138 4.5005
R60419 VINN.n272 VINN.n138 4.5005
R60420 VINN.n288 VINN.n138 4.5005
R60421 VINN.n271 VINN.n138 4.5005
R60422 VINN.n290 VINN.n138 4.5005
R60423 VINN.n270 VINN.n138 4.5005
R60424 VINN.n292 VINN.n138 4.5005
R60425 VINN.n269 VINN.n138 4.5005
R60426 VINN.n294 VINN.n138 4.5005
R60427 VINN.n268 VINN.n138 4.5005
R60428 VINN.n296 VINN.n138 4.5005
R60429 VINN.n267 VINN.n138 4.5005
R60430 VINN.n298 VINN.n138 4.5005
R60431 VINN.n266 VINN.n138 4.5005
R60432 VINN.n300 VINN.n138 4.5005
R60433 VINN.n265 VINN.n138 4.5005
R60434 VINN.n302 VINN.n138 4.5005
R60435 VINN.n264 VINN.n138 4.5005
R60436 VINN.n304 VINN.n138 4.5005
R60437 VINN.n263 VINN.n138 4.5005
R60438 VINN.n306 VINN.n138 4.5005
R60439 VINN.n262 VINN.n138 4.5005
R60440 VINN.n308 VINN.n138 4.5005
R60441 VINN.n261 VINN.n138 4.5005
R60442 VINN.n310 VINN.n138 4.5005
R60443 VINN.n260 VINN.n138 4.5005
R60444 VINN.n312 VINN.n138 4.5005
R60445 VINN.n259 VINN.n138 4.5005
R60446 VINN.n314 VINN.n138 4.5005
R60447 VINN.n258 VINN.n138 4.5005
R60448 VINN.n316 VINN.n138 4.5005
R60449 VINN.n257 VINN.n138 4.5005
R60450 VINN.n318 VINN.n138 4.5005
R60451 VINN.n256 VINN.n138 4.5005
R60452 VINN.n320 VINN.n138 4.5005
R60453 VINN.n255 VINN.n138 4.5005
R60454 VINN.n322 VINN.n138 4.5005
R60455 VINN.n254 VINN.n138 4.5005
R60456 VINN.n324 VINN.n138 4.5005
R60457 VINN.n253 VINN.n138 4.5005
R60458 VINN.n326 VINN.n138 4.5005
R60459 VINN.n252 VINN.n138 4.5005
R60460 VINN.n328 VINN.n138 4.5005
R60461 VINN.n251 VINN.n138 4.5005
R60462 VINN.n330 VINN.n138 4.5005
R60463 VINN.n250 VINN.n138 4.5005
R60464 VINN.n332 VINN.n138 4.5005
R60465 VINN.n249 VINN.n138 4.5005
R60466 VINN.n334 VINN.n138 4.5005
R60467 VINN.n248 VINN.n138 4.5005
R60468 VINN.n336 VINN.n138 4.5005
R60469 VINN.n247 VINN.n138 4.5005
R60470 VINN.n338 VINN.n138 4.5005
R60471 VINN.n246 VINN.n138 4.5005
R60472 VINN.n340 VINN.n138 4.5005
R60473 VINN.n245 VINN.n138 4.5005
R60474 VINN.n342 VINN.n138 4.5005
R60475 VINN.n244 VINN.n138 4.5005
R60476 VINN.n344 VINN.n138 4.5005
R60477 VINN.n243 VINN.n138 4.5005
R60478 VINN.n346 VINN.n138 4.5005
R60479 VINN.n242 VINN.n138 4.5005
R60480 VINN.n348 VINN.n138 4.5005
R60481 VINN.n241 VINN.n138 4.5005
R60482 VINN.n350 VINN.n138 4.5005
R60483 VINN.n240 VINN.n138 4.5005
R60484 VINN.n352 VINN.n138 4.5005
R60485 VINN.n239 VINN.n138 4.5005
R60486 VINN.n354 VINN.n138 4.5005
R60487 VINN.n238 VINN.n138 4.5005
R60488 VINN.n356 VINN.n138 4.5005
R60489 VINN.n237 VINN.n138 4.5005
R60490 VINN.n358 VINN.n138 4.5005
R60491 VINN.n236 VINN.n138 4.5005
R60492 VINN.n360 VINN.n138 4.5005
R60493 VINN.n235 VINN.n138 4.5005
R60494 VINN.n362 VINN.n138 4.5005
R60495 VINN.n234 VINN.n138 4.5005
R60496 VINN.n364 VINN.n138 4.5005
R60497 VINN.n233 VINN.n138 4.5005
R60498 VINN.n366 VINN.n138 4.5005
R60499 VINN.n232 VINN.n138 4.5005
R60500 VINN.n368 VINN.n138 4.5005
R60501 VINN.n231 VINN.n138 4.5005
R60502 VINN.n370 VINN.n138 4.5005
R60503 VINN.n230 VINN.n138 4.5005
R60504 VINN.n372 VINN.n138 4.5005
R60505 VINN.n229 VINN.n138 4.5005
R60506 VINN.n374 VINN.n138 4.5005
R60507 VINN.n228 VINN.n138 4.5005
R60508 VINN.n376 VINN.n138 4.5005
R60509 VINN.n227 VINN.n138 4.5005
R60510 VINN.n378 VINN.n138 4.5005
R60511 VINN.n226 VINN.n138 4.5005
R60512 VINN.n380 VINN.n138 4.5005
R60513 VINN.n225 VINN.n138 4.5005
R60514 VINN.n382 VINN.n138 4.5005
R60515 VINN.n224 VINN.n138 4.5005
R60516 VINN.n384 VINN.n138 4.5005
R60517 VINN.n223 VINN.n138 4.5005
R60518 VINN.n386 VINN.n138 4.5005
R60519 VINN.n222 VINN.n138 4.5005
R60520 VINN.n388 VINN.n138 4.5005
R60521 VINN.n221 VINN.n138 4.5005
R60522 VINN.n390 VINN.n138 4.5005
R60523 VINN.n220 VINN.n138 4.5005
R60524 VINN.n392 VINN.n138 4.5005
R60525 VINN.n219 VINN.n138 4.5005
R60526 VINN.n394 VINN.n138 4.5005
R60527 VINN.n218 VINN.n138 4.5005
R60528 VINN.n396 VINN.n138 4.5005
R60529 VINN.n217 VINN.n138 4.5005
R60530 VINN.n398 VINN.n138 4.5005
R60531 VINN.n216 VINN.n138 4.5005
R60532 VINN.n400 VINN.n138 4.5005
R60533 VINN.n215 VINN.n138 4.5005
R60534 VINN.n654 VINN.n138 4.5005
R60535 VINN.n656 VINN.n138 4.5005
R60536 VINN.n138 VINN.n0 4.5005
R60537 VINN.n278 VINN.n163 4.5005
R60538 VINN.n276 VINN.n163 4.5005
R60539 VINN.n280 VINN.n163 4.5005
R60540 VINN.n275 VINN.n163 4.5005
R60541 VINN.n282 VINN.n163 4.5005
R60542 VINN.n274 VINN.n163 4.5005
R60543 VINN.n284 VINN.n163 4.5005
R60544 VINN.n273 VINN.n163 4.5005
R60545 VINN.n286 VINN.n163 4.5005
R60546 VINN.n272 VINN.n163 4.5005
R60547 VINN.n288 VINN.n163 4.5005
R60548 VINN.n271 VINN.n163 4.5005
R60549 VINN.n290 VINN.n163 4.5005
R60550 VINN.n270 VINN.n163 4.5005
R60551 VINN.n292 VINN.n163 4.5005
R60552 VINN.n269 VINN.n163 4.5005
R60553 VINN.n294 VINN.n163 4.5005
R60554 VINN.n268 VINN.n163 4.5005
R60555 VINN.n296 VINN.n163 4.5005
R60556 VINN.n267 VINN.n163 4.5005
R60557 VINN.n298 VINN.n163 4.5005
R60558 VINN.n266 VINN.n163 4.5005
R60559 VINN.n300 VINN.n163 4.5005
R60560 VINN.n265 VINN.n163 4.5005
R60561 VINN.n302 VINN.n163 4.5005
R60562 VINN.n264 VINN.n163 4.5005
R60563 VINN.n304 VINN.n163 4.5005
R60564 VINN.n263 VINN.n163 4.5005
R60565 VINN.n306 VINN.n163 4.5005
R60566 VINN.n262 VINN.n163 4.5005
R60567 VINN.n308 VINN.n163 4.5005
R60568 VINN.n261 VINN.n163 4.5005
R60569 VINN.n310 VINN.n163 4.5005
R60570 VINN.n260 VINN.n163 4.5005
R60571 VINN.n312 VINN.n163 4.5005
R60572 VINN.n259 VINN.n163 4.5005
R60573 VINN.n314 VINN.n163 4.5005
R60574 VINN.n258 VINN.n163 4.5005
R60575 VINN.n316 VINN.n163 4.5005
R60576 VINN.n257 VINN.n163 4.5005
R60577 VINN.n318 VINN.n163 4.5005
R60578 VINN.n256 VINN.n163 4.5005
R60579 VINN.n320 VINN.n163 4.5005
R60580 VINN.n255 VINN.n163 4.5005
R60581 VINN.n322 VINN.n163 4.5005
R60582 VINN.n254 VINN.n163 4.5005
R60583 VINN.n324 VINN.n163 4.5005
R60584 VINN.n253 VINN.n163 4.5005
R60585 VINN.n326 VINN.n163 4.5005
R60586 VINN.n252 VINN.n163 4.5005
R60587 VINN.n328 VINN.n163 4.5005
R60588 VINN.n251 VINN.n163 4.5005
R60589 VINN.n330 VINN.n163 4.5005
R60590 VINN.n250 VINN.n163 4.5005
R60591 VINN.n332 VINN.n163 4.5005
R60592 VINN.n249 VINN.n163 4.5005
R60593 VINN.n334 VINN.n163 4.5005
R60594 VINN.n248 VINN.n163 4.5005
R60595 VINN.n336 VINN.n163 4.5005
R60596 VINN.n247 VINN.n163 4.5005
R60597 VINN.n338 VINN.n163 4.5005
R60598 VINN.n246 VINN.n163 4.5005
R60599 VINN.n340 VINN.n163 4.5005
R60600 VINN.n245 VINN.n163 4.5005
R60601 VINN.n342 VINN.n163 4.5005
R60602 VINN.n244 VINN.n163 4.5005
R60603 VINN.n344 VINN.n163 4.5005
R60604 VINN.n243 VINN.n163 4.5005
R60605 VINN.n346 VINN.n163 4.5005
R60606 VINN.n242 VINN.n163 4.5005
R60607 VINN.n348 VINN.n163 4.5005
R60608 VINN.n241 VINN.n163 4.5005
R60609 VINN.n350 VINN.n163 4.5005
R60610 VINN.n240 VINN.n163 4.5005
R60611 VINN.n352 VINN.n163 4.5005
R60612 VINN.n239 VINN.n163 4.5005
R60613 VINN.n354 VINN.n163 4.5005
R60614 VINN.n238 VINN.n163 4.5005
R60615 VINN.n356 VINN.n163 4.5005
R60616 VINN.n237 VINN.n163 4.5005
R60617 VINN.n358 VINN.n163 4.5005
R60618 VINN.n236 VINN.n163 4.5005
R60619 VINN.n360 VINN.n163 4.5005
R60620 VINN.n235 VINN.n163 4.5005
R60621 VINN.n362 VINN.n163 4.5005
R60622 VINN.n234 VINN.n163 4.5005
R60623 VINN.n364 VINN.n163 4.5005
R60624 VINN.n233 VINN.n163 4.5005
R60625 VINN.n366 VINN.n163 4.5005
R60626 VINN.n232 VINN.n163 4.5005
R60627 VINN.n368 VINN.n163 4.5005
R60628 VINN.n231 VINN.n163 4.5005
R60629 VINN.n370 VINN.n163 4.5005
R60630 VINN.n230 VINN.n163 4.5005
R60631 VINN.n372 VINN.n163 4.5005
R60632 VINN.n229 VINN.n163 4.5005
R60633 VINN.n374 VINN.n163 4.5005
R60634 VINN.n228 VINN.n163 4.5005
R60635 VINN.n376 VINN.n163 4.5005
R60636 VINN.n227 VINN.n163 4.5005
R60637 VINN.n378 VINN.n163 4.5005
R60638 VINN.n226 VINN.n163 4.5005
R60639 VINN.n380 VINN.n163 4.5005
R60640 VINN.n225 VINN.n163 4.5005
R60641 VINN.n382 VINN.n163 4.5005
R60642 VINN.n224 VINN.n163 4.5005
R60643 VINN.n384 VINN.n163 4.5005
R60644 VINN.n223 VINN.n163 4.5005
R60645 VINN.n386 VINN.n163 4.5005
R60646 VINN.n222 VINN.n163 4.5005
R60647 VINN.n388 VINN.n163 4.5005
R60648 VINN.n221 VINN.n163 4.5005
R60649 VINN.n390 VINN.n163 4.5005
R60650 VINN.n220 VINN.n163 4.5005
R60651 VINN.n392 VINN.n163 4.5005
R60652 VINN.n219 VINN.n163 4.5005
R60653 VINN.n394 VINN.n163 4.5005
R60654 VINN.n218 VINN.n163 4.5005
R60655 VINN.n396 VINN.n163 4.5005
R60656 VINN.n217 VINN.n163 4.5005
R60657 VINN.n398 VINN.n163 4.5005
R60658 VINN.n216 VINN.n163 4.5005
R60659 VINN.n400 VINN.n163 4.5005
R60660 VINN.n215 VINN.n163 4.5005
R60661 VINN.n654 VINN.n163 4.5005
R60662 VINN.n656 VINN.n163 4.5005
R60663 VINN.n163 VINN.n0 4.5005
R60664 VINN.n278 VINN.n137 4.5005
R60665 VINN.n276 VINN.n137 4.5005
R60666 VINN.n280 VINN.n137 4.5005
R60667 VINN.n275 VINN.n137 4.5005
R60668 VINN.n282 VINN.n137 4.5005
R60669 VINN.n274 VINN.n137 4.5005
R60670 VINN.n284 VINN.n137 4.5005
R60671 VINN.n273 VINN.n137 4.5005
R60672 VINN.n286 VINN.n137 4.5005
R60673 VINN.n272 VINN.n137 4.5005
R60674 VINN.n288 VINN.n137 4.5005
R60675 VINN.n271 VINN.n137 4.5005
R60676 VINN.n290 VINN.n137 4.5005
R60677 VINN.n270 VINN.n137 4.5005
R60678 VINN.n292 VINN.n137 4.5005
R60679 VINN.n269 VINN.n137 4.5005
R60680 VINN.n294 VINN.n137 4.5005
R60681 VINN.n268 VINN.n137 4.5005
R60682 VINN.n296 VINN.n137 4.5005
R60683 VINN.n267 VINN.n137 4.5005
R60684 VINN.n298 VINN.n137 4.5005
R60685 VINN.n266 VINN.n137 4.5005
R60686 VINN.n300 VINN.n137 4.5005
R60687 VINN.n265 VINN.n137 4.5005
R60688 VINN.n302 VINN.n137 4.5005
R60689 VINN.n264 VINN.n137 4.5005
R60690 VINN.n304 VINN.n137 4.5005
R60691 VINN.n263 VINN.n137 4.5005
R60692 VINN.n306 VINN.n137 4.5005
R60693 VINN.n262 VINN.n137 4.5005
R60694 VINN.n308 VINN.n137 4.5005
R60695 VINN.n261 VINN.n137 4.5005
R60696 VINN.n310 VINN.n137 4.5005
R60697 VINN.n260 VINN.n137 4.5005
R60698 VINN.n312 VINN.n137 4.5005
R60699 VINN.n259 VINN.n137 4.5005
R60700 VINN.n314 VINN.n137 4.5005
R60701 VINN.n258 VINN.n137 4.5005
R60702 VINN.n316 VINN.n137 4.5005
R60703 VINN.n257 VINN.n137 4.5005
R60704 VINN.n318 VINN.n137 4.5005
R60705 VINN.n256 VINN.n137 4.5005
R60706 VINN.n320 VINN.n137 4.5005
R60707 VINN.n255 VINN.n137 4.5005
R60708 VINN.n322 VINN.n137 4.5005
R60709 VINN.n254 VINN.n137 4.5005
R60710 VINN.n324 VINN.n137 4.5005
R60711 VINN.n253 VINN.n137 4.5005
R60712 VINN.n326 VINN.n137 4.5005
R60713 VINN.n252 VINN.n137 4.5005
R60714 VINN.n328 VINN.n137 4.5005
R60715 VINN.n251 VINN.n137 4.5005
R60716 VINN.n330 VINN.n137 4.5005
R60717 VINN.n250 VINN.n137 4.5005
R60718 VINN.n332 VINN.n137 4.5005
R60719 VINN.n249 VINN.n137 4.5005
R60720 VINN.n334 VINN.n137 4.5005
R60721 VINN.n248 VINN.n137 4.5005
R60722 VINN.n336 VINN.n137 4.5005
R60723 VINN.n247 VINN.n137 4.5005
R60724 VINN.n338 VINN.n137 4.5005
R60725 VINN.n246 VINN.n137 4.5005
R60726 VINN.n340 VINN.n137 4.5005
R60727 VINN.n245 VINN.n137 4.5005
R60728 VINN.n342 VINN.n137 4.5005
R60729 VINN.n244 VINN.n137 4.5005
R60730 VINN.n344 VINN.n137 4.5005
R60731 VINN.n243 VINN.n137 4.5005
R60732 VINN.n346 VINN.n137 4.5005
R60733 VINN.n242 VINN.n137 4.5005
R60734 VINN.n348 VINN.n137 4.5005
R60735 VINN.n241 VINN.n137 4.5005
R60736 VINN.n350 VINN.n137 4.5005
R60737 VINN.n240 VINN.n137 4.5005
R60738 VINN.n352 VINN.n137 4.5005
R60739 VINN.n239 VINN.n137 4.5005
R60740 VINN.n354 VINN.n137 4.5005
R60741 VINN.n238 VINN.n137 4.5005
R60742 VINN.n356 VINN.n137 4.5005
R60743 VINN.n237 VINN.n137 4.5005
R60744 VINN.n358 VINN.n137 4.5005
R60745 VINN.n236 VINN.n137 4.5005
R60746 VINN.n360 VINN.n137 4.5005
R60747 VINN.n235 VINN.n137 4.5005
R60748 VINN.n362 VINN.n137 4.5005
R60749 VINN.n234 VINN.n137 4.5005
R60750 VINN.n364 VINN.n137 4.5005
R60751 VINN.n233 VINN.n137 4.5005
R60752 VINN.n366 VINN.n137 4.5005
R60753 VINN.n232 VINN.n137 4.5005
R60754 VINN.n368 VINN.n137 4.5005
R60755 VINN.n231 VINN.n137 4.5005
R60756 VINN.n370 VINN.n137 4.5005
R60757 VINN.n230 VINN.n137 4.5005
R60758 VINN.n372 VINN.n137 4.5005
R60759 VINN.n229 VINN.n137 4.5005
R60760 VINN.n374 VINN.n137 4.5005
R60761 VINN.n228 VINN.n137 4.5005
R60762 VINN.n376 VINN.n137 4.5005
R60763 VINN.n227 VINN.n137 4.5005
R60764 VINN.n378 VINN.n137 4.5005
R60765 VINN.n226 VINN.n137 4.5005
R60766 VINN.n380 VINN.n137 4.5005
R60767 VINN.n225 VINN.n137 4.5005
R60768 VINN.n382 VINN.n137 4.5005
R60769 VINN.n224 VINN.n137 4.5005
R60770 VINN.n384 VINN.n137 4.5005
R60771 VINN.n223 VINN.n137 4.5005
R60772 VINN.n386 VINN.n137 4.5005
R60773 VINN.n222 VINN.n137 4.5005
R60774 VINN.n388 VINN.n137 4.5005
R60775 VINN.n221 VINN.n137 4.5005
R60776 VINN.n390 VINN.n137 4.5005
R60777 VINN.n220 VINN.n137 4.5005
R60778 VINN.n392 VINN.n137 4.5005
R60779 VINN.n219 VINN.n137 4.5005
R60780 VINN.n394 VINN.n137 4.5005
R60781 VINN.n218 VINN.n137 4.5005
R60782 VINN.n396 VINN.n137 4.5005
R60783 VINN.n217 VINN.n137 4.5005
R60784 VINN.n398 VINN.n137 4.5005
R60785 VINN.n216 VINN.n137 4.5005
R60786 VINN.n400 VINN.n137 4.5005
R60787 VINN.n215 VINN.n137 4.5005
R60788 VINN.n654 VINN.n137 4.5005
R60789 VINN.n656 VINN.n137 4.5005
R60790 VINN.n137 VINN.n0 4.5005
R60791 VINN.n278 VINN.n164 4.5005
R60792 VINN.n276 VINN.n164 4.5005
R60793 VINN.n280 VINN.n164 4.5005
R60794 VINN.n275 VINN.n164 4.5005
R60795 VINN.n282 VINN.n164 4.5005
R60796 VINN.n274 VINN.n164 4.5005
R60797 VINN.n284 VINN.n164 4.5005
R60798 VINN.n273 VINN.n164 4.5005
R60799 VINN.n286 VINN.n164 4.5005
R60800 VINN.n272 VINN.n164 4.5005
R60801 VINN.n288 VINN.n164 4.5005
R60802 VINN.n271 VINN.n164 4.5005
R60803 VINN.n290 VINN.n164 4.5005
R60804 VINN.n270 VINN.n164 4.5005
R60805 VINN.n292 VINN.n164 4.5005
R60806 VINN.n269 VINN.n164 4.5005
R60807 VINN.n294 VINN.n164 4.5005
R60808 VINN.n268 VINN.n164 4.5005
R60809 VINN.n296 VINN.n164 4.5005
R60810 VINN.n267 VINN.n164 4.5005
R60811 VINN.n298 VINN.n164 4.5005
R60812 VINN.n266 VINN.n164 4.5005
R60813 VINN.n300 VINN.n164 4.5005
R60814 VINN.n265 VINN.n164 4.5005
R60815 VINN.n302 VINN.n164 4.5005
R60816 VINN.n264 VINN.n164 4.5005
R60817 VINN.n304 VINN.n164 4.5005
R60818 VINN.n263 VINN.n164 4.5005
R60819 VINN.n306 VINN.n164 4.5005
R60820 VINN.n262 VINN.n164 4.5005
R60821 VINN.n308 VINN.n164 4.5005
R60822 VINN.n261 VINN.n164 4.5005
R60823 VINN.n310 VINN.n164 4.5005
R60824 VINN.n260 VINN.n164 4.5005
R60825 VINN.n312 VINN.n164 4.5005
R60826 VINN.n259 VINN.n164 4.5005
R60827 VINN.n314 VINN.n164 4.5005
R60828 VINN.n258 VINN.n164 4.5005
R60829 VINN.n316 VINN.n164 4.5005
R60830 VINN.n257 VINN.n164 4.5005
R60831 VINN.n318 VINN.n164 4.5005
R60832 VINN.n256 VINN.n164 4.5005
R60833 VINN.n320 VINN.n164 4.5005
R60834 VINN.n255 VINN.n164 4.5005
R60835 VINN.n322 VINN.n164 4.5005
R60836 VINN.n254 VINN.n164 4.5005
R60837 VINN.n324 VINN.n164 4.5005
R60838 VINN.n253 VINN.n164 4.5005
R60839 VINN.n326 VINN.n164 4.5005
R60840 VINN.n252 VINN.n164 4.5005
R60841 VINN.n328 VINN.n164 4.5005
R60842 VINN.n251 VINN.n164 4.5005
R60843 VINN.n330 VINN.n164 4.5005
R60844 VINN.n250 VINN.n164 4.5005
R60845 VINN.n332 VINN.n164 4.5005
R60846 VINN.n249 VINN.n164 4.5005
R60847 VINN.n334 VINN.n164 4.5005
R60848 VINN.n248 VINN.n164 4.5005
R60849 VINN.n336 VINN.n164 4.5005
R60850 VINN.n247 VINN.n164 4.5005
R60851 VINN.n338 VINN.n164 4.5005
R60852 VINN.n246 VINN.n164 4.5005
R60853 VINN.n340 VINN.n164 4.5005
R60854 VINN.n245 VINN.n164 4.5005
R60855 VINN.n342 VINN.n164 4.5005
R60856 VINN.n244 VINN.n164 4.5005
R60857 VINN.n344 VINN.n164 4.5005
R60858 VINN.n243 VINN.n164 4.5005
R60859 VINN.n346 VINN.n164 4.5005
R60860 VINN.n242 VINN.n164 4.5005
R60861 VINN.n348 VINN.n164 4.5005
R60862 VINN.n241 VINN.n164 4.5005
R60863 VINN.n350 VINN.n164 4.5005
R60864 VINN.n240 VINN.n164 4.5005
R60865 VINN.n352 VINN.n164 4.5005
R60866 VINN.n239 VINN.n164 4.5005
R60867 VINN.n354 VINN.n164 4.5005
R60868 VINN.n238 VINN.n164 4.5005
R60869 VINN.n356 VINN.n164 4.5005
R60870 VINN.n237 VINN.n164 4.5005
R60871 VINN.n358 VINN.n164 4.5005
R60872 VINN.n236 VINN.n164 4.5005
R60873 VINN.n360 VINN.n164 4.5005
R60874 VINN.n235 VINN.n164 4.5005
R60875 VINN.n362 VINN.n164 4.5005
R60876 VINN.n234 VINN.n164 4.5005
R60877 VINN.n364 VINN.n164 4.5005
R60878 VINN.n233 VINN.n164 4.5005
R60879 VINN.n366 VINN.n164 4.5005
R60880 VINN.n232 VINN.n164 4.5005
R60881 VINN.n368 VINN.n164 4.5005
R60882 VINN.n231 VINN.n164 4.5005
R60883 VINN.n370 VINN.n164 4.5005
R60884 VINN.n230 VINN.n164 4.5005
R60885 VINN.n372 VINN.n164 4.5005
R60886 VINN.n229 VINN.n164 4.5005
R60887 VINN.n374 VINN.n164 4.5005
R60888 VINN.n228 VINN.n164 4.5005
R60889 VINN.n376 VINN.n164 4.5005
R60890 VINN.n227 VINN.n164 4.5005
R60891 VINN.n378 VINN.n164 4.5005
R60892 VINN.n226 VINN.n164 4.5005
R60893 VINN.n380 VINN.n164 4.5005
R60894 VINN.n225 VINN.n164 4.5005
R60895 VINN.n382 VINN.n164 4.5005
R60896 VINN.n224 VINN.n164 4.5005
R60897 VINN.n384 VINN.n164 4.5005
R60898 VINN.n223 VINN.n164 4.5005
R60899 VINN.n386 VINN.n164 4.5005
R60900 VINN.n222 VINN.n164 4.5005
R60901 VINN.n388 VINN.n164 4.5005
R60902 VINN.n221 VINN.n164 4.5005
R60903 VINN.n390 VINN.n164 4.5005
R60904 VINN.n220 VINN.n164 4.5005
R60905 VINN.n392 VINN.n164 4.5005
R60906 VINN.n219 VINN.n164 4.5005
R60907 VINN.n394 VINN.n164 4.5005
R60908 VINN.n218 VINN.n164 4.5005
R60909 VINN.n396 VINN.n164 4.5005
R60910 VINN.n217 VINN.n164 4.5005
R60911 VINN.n398 VINN.n164 4.5005
R60912 VINN.n216 VINN.n164 4.5005
R60913 VINN.n400 VINN.n164 4.5005
R60914 VINN.n215 VINN.n164 4.5005
R60915 VINN.n654 VINN.n164 4.5005
R60916 VINN.n656 VINN.n164 4.5005
R60917 VINN.n164 VINN.n0 4.5005
R60918 VINN.n278 VINN.n136 4.5005
R60919 VINN.n276 VINN.n136 4.5005
R60920 VINN.n280 VINN.n136 4.5005
R60921 VINN.n275 VINN.n136 4.5005
R60922 VINN.n282 VINN.n136 4.5005
R60923 VINN.n274 VINN.n136 4.5005
R60924 VINN.n284 VINN.n136 4.5005
R60925 VINN.n273 VINN.n136 4.5005
R60926 VINN.n286 VINN.n136 4.5005
R60927 VINN.n272 VINN.n136 4.5005
R60928 VINN.n288 VINN.n136 4.5005
R60929 VINN.n271 VINN.n136 4.5005
R60930 VINN.n290 VINN.n136 4.5005
R60931 VINN.n270 VINN.n136 4.5005
R60932 VINN.n292 VINN.n136 4.5005
R60933 VINN.n269 VINN.n136 4.5005
R60934 VINN.n294 VINN.n136 4.5005
R60935 VINN.n268 VINN.n136 4.5005
R60936 VINN.n296 VINN.n136 4.5005
R60937 VINN.n267 VINN.n136 4.5005
R60938 VINN.n298 VINN.n136 4.5005
R60939 VINN.n266 VINN.n136 4.5005
R60940 VINN.n300 VINN.n136 4.5005
R60941 VINN.n265 VINN.n136 4.5005
R60942 VINN.n302 VINN.n136 4.5005
R60943 VINN.n264 VINN.n136 4.5005
R60944 VINN.n304 VINN.n136 4.5005
R60945 VINN.n263 VINN.n136 4.5005
R60946 VINN.n306 VINN.n136 4.5005
R60947 VINN.n262 VINN.n136 4.5005
R60948 VINN.n308 VINN.n136 4.5005
R60949 VINN.n261 VINN.n136 4.5005
R60950 VINN.n310 VINN.n136 4.5005
R60951 VINN.n260 VINN.n136 4.5005
R60952 VINN.n312 VINN.n136 4.5005
R60953 VINN.n259 VINN.n136 4.5005
R60954 VINN.n314 VINN.n136 4.5005
R60955 VINN.n258 VINN.n136 4.5005
R60956 VINN.n316 VINN.n136 4.5005
R60957 VINN.n257 VINN.n136 4.5005
R60958 VINN.n318 VINN.n136 4.5005
R60959 VINN.n256 VINN.n136 4.5005
R60960 VINN.n320 VINN.n136 4.5005
R60961 VINN.n255 VINN.n136 4.5005
R60962 VINN.n322 VINN.n136 4.5005
R60963 VINN.n254 VINN.n136 4.5005
R60964 VINN.n324 VINN.n136 4.5005
R60965 VINN.n253 VINN.n136 4.5005
R60966 VINN.n326 VINN.n136 4.5005
R60967 VINN.n252 VINN.n136 4.5005
R60968 VINN.n328 VINN.n136 4.5005
R60969 VINN.n251 VINN.n136 4.5005
R60970 VINN.n330 VINN.n136 4.5005
R60971 VINN.n250 VINN.n136 4.5005
R60972 VINN.n332 VINN.n136 4.5005
R60973 VINN.n249 VINN.n136 4.5005
R60974 VINN.n334 VINN.n136 4.5005
R60975 VINN.n248 VINN.n136 4.5005
R60976 VINN.n336 VINN.n136 4.5005
R60977 VINN.n247 VINN.n136 4.5005
R60978 VINN.n338 VINN.n136 4.5005
R60979 VINN.n246 VINN.n136 4.5005
R60980 VINN.n340 VINN.n136 4.5005
R60981 VINN.n245 VINN.n136 4.5005
R60982 VINN.n342 VINN.n136 4.5005
R60983 VINN.n244 VINN.n136 4.5005
R60984 VINN.n344 VINN.n136 4.5005
R60985 VINN.n243 VINN.n136 4.5005
R60986 VINN.n346 VINN.n136 4.5005
R60987 VINN.n242 VINN.n136 4.5005
R60988 VINN.n348 VINN.n136 4.5005
R60989 VINN.n241 VINN.n136 4.5005
R60990 VINN.n350 VINN.n136 4.5005
R60991 VINN.n240 VINN.n136 4.5005
R60992 VINN.n352 VINN.n136 4.5005
R60993 VINN.n239 VINN.n136 4.5005
R60994 VINN.n354 VINN.n136 4.5005
R60995 VINN.n238 VINN.n136 4.5005
R60996 VINN.n356 VINN.n136 4.5005
R60997 VINN.n237 VINN.n136 4.5005
R60998 VINN.n358 VINN.n136 4.5005
R60999 VINN.n236 VINN.n136 4.5005
R61000 VINN.n360 VINN.n136 4.5005
R61001 VINN.n235 VINN.n136 4.5005
R61002 VINN.n362 VINN.n136 4.5005
R61003 VINN.n234 VINN.n136 4.5005
R61004 VINN.n364 VINN.n136 4.5005
R61005 VINN.n233 VINN.n136 4.5005
R61006 VINN.n366 VINN.n136 4.5005
R61007 VINN.n232 VINN.n136 4.5005
R61008 VINN.n368 VINN.n136 4.5005
R61009 VINN.n231 VINN.n136 4.5005
R61010 VINN.n370 VINN.n136 4.5005
R61011 VINN.n230 VINN.n136 4.5005
R61012 VINN.n372 VINN.n136 4.5005
R61013 VINN.n229 VINN.n136 4.5005
R61014 VINN.n374 VINN.n136 4.5005
R61015 VINN.n228 VINN.n136 4.5005
R61016 VINN.n376 VINN.n136 4.5005
R61017 VINN.n227 VINN.n136 4.5005
R61018 VINN.n378 VINN.n136 4.5005
R61019 VINN.n226 VINN.n136 4.5005
R61020 VINN.n380 VINN.n136 4.5005
R61021 VINN.n225 VINN.n136 4.5005
R61022 VINN.n382 VINN.n136 4.5005
R61023 VINN.n224 VINN.n136 4.5005
R61024 VINN.n384 VINN.n136 4.5005
R61025 VINN.n223 VINN.n136 4.5005
R61026 VINN.n386 VINN.n136 4.5005
R61027 VINN.n222 VINN.n136 4.5005
R61028 VINN.n388 VINN.n136 4.5005
R61029 VINN.n221 VINN.n136 4.5005
R61030 VINN.n390 VINN.n136 4.5005
R61031 VINN.n220 VINN.n136 4.5005
R61032 VINN.n392 VINN.n136 4.5005
R61033 VINN.n219 VINN.n136 4.5005
R61034 VINN.n394 VINN.n136 4.5005
R61035 VINN.n218 VINN.n136 4.5005
R61036 VINN.n396 VINN.n136 4.5005
R61037 VINN.n217 VINN.n136 4.5005
R61038 VINN.n398 VINN.n136 4.5005
R61039 VINN.n216 VINN.n136 4.5005
R61040 VINN.n400 VINN.n136 4.5005
R61041 VINN.n215 VINN.n136 4.5005
R61042 VINN.n654 VINN.n136 4.5005
R61043 VINN.n656 VINN.n136 4.5005
R61044 VINN.n136 VINN.n0 4.5005
R61045 VINN.n278 VINN.n165 4.5005
R61046 VINN.n276 VINN.n165 4.5005
R61047 VINN.n280 VINN.n165 4.5005
R61048 VINN.n275 VINN.n165 4.5005
R61049 VINN.n282 VINN.n165 4.5005
R61050 VINN.n274 VINN.n165 4.5005
R61051 VINN.n284 VINN.n165 4.5005
R61052 VINN.n273 VINN.n165 4.5005
R61053 VINN.n286 VINN.n165 4.5005
R61054 VINN.n272 VINN.n165 4.5005
R61055 VINN.n288 VINN.n165 4.5005
R61056 VINN.n271 VINN.n165 4.5005
R61057 VINN.n290 VINN.n165 4.5005
R61058 VINN.n270 VINN.n165 4.5005
R61059 VINN.n292 VINN.n165 4.5005
R61060 VINN.n269 VINN.n165 4.5005
R61061 VINN.n294 VINN.n165 4.5005
R61062 VINN.n268 VINN.n165 4.5005
R61063 VINN.n296 VINN.n165 4.5005
R61064 VINN.n267 VINN.n165 4.5005
R61065 VINN.n298 VINN.n165 4.5005
R61066 VINN.n266 VINN.n165 4.5005
R61067 VINN.n300 VINN.n165 4.5005
R61068 VINN.n265 VINN.n165 4.5005
R61069 VINN.n302 VINN.n165 4.5005
R61070 VINN.n264 VINN.n165 4.5005
R61071 VINN.n304 VINN.n165 4.5005
R61072 VINN.n263 VINN.n165 4.5005
R61073 VINN.n306 VINN.n165 4.5005
R61074 VINN.n262 VINN.n165 4.5005
R61075 VINN.n308 VINN.n165 4.5005
R61076 VINN.n261 VINN.n165 4.5005
R61077 VINN.n310 VINN.n165 4.5005
R61078 VINN.n260 VINN.n165 4.5005
R61079 VINN.n312 VINN.n165 4.5005
R61080 VINN.n259 VINN.n165 4.5005
R61081 VINN.n314 VINN.n165 4.5005
R61082 VINN.n258 VINN.n165 4.5005
R61083 VINN.n316 VINN.n165 4.5005
R61084 VINN.n257 VINN.n165 4.5005
R61085 VINN.n318 VINN.n165 4.5005
R61086 VINN.n256 VINN.n165 4.5005
R61087 VINN.n320 VINN.n165 4.5005
R61088 VINN.n255 VINN.n165 4.5005
R61089 VINN.n322 VINN.n165 4.5005
R61090 VINN.n254 VINN.n165 4.5005
R61091 VINN.n324 VINN.n165 4.5005
R61092 VINN.n253 VINN.n165 4.5005
R61093 VINN.n326 VINN.n165 4.5005
R61094 VINN.n252 VINN.n165 4.5005
R61095 VINN.n328 VINN.n165 4.5005
R61096 VINN.n251 VINN.n165 4.5005
R61097 VINN.n330 VINN.n165 4.5005
R61098 VINN.n250 VINN.n165 4.5005
R61099 VINN.n332 VINN.n165 4.5005
R61100 VINN.n249 VINN.n165 4.5005
R61101 VINN.n334 VINN.n165 4.5005
R61102 VINN.n248 VINN.n165 4.5005
R61103 VINN.n336 VINN.n165 4.5005
R61104 VINN.n247 VINN.n165 4.5005
R61105 VINN.n338 VINN.n165 4.5005
R61106 VINN.n246 VINN.n165 4.5005
R61107 VINN.n340 VINN.n165 4.5005
R61108 VINN.n245 VINN.n165 4.5005
R61109 VINN.n342 VINN.n165 4.5005
R61110 VINN.n244 VINN.n165 4.5005
R61111 VINN.n344 VINN.n165 4.5005
R61112 VINN.n243 VINN.n165 4.5005
R61113 VINN.n346 VINN.n165 4.5005
R61114 VINN.n242 VINN.n165 4.5005
R61115 VINN.n348 VINN.n165 4.5005
R61116 VINN.n241 VINN.n165 4.5005
R61117 VINN.n350 VINN.n165 4.5005
R61118 VINN.n240 VINN.n165 4.5005
R61119 VINN.n352 VINN.n165 4.5005
R61120 VINN.n239 VINN.n165 4.5005
R61121 VINN.n354 VINN.n165 4.5005
R61122 VINN.n238 VINN.n165 4.5005
R61123 VINN.n356 VINN.n165 4.5005
R61124 VINN.n237 VINN.n165 4.5005
R61125 VINN.n358 VINN.n165 4.5005
R61126 VINN.n236 VINN.n165 4.5005
R61127 VINN.n360 VINN.n165 4.5005
R61128 VINN.n235 VINN.n165 4.5005
R61129 VINN.n362 VINN.n165 4.5005
R61130 VINN.n234 VINN.n165 4.5005
R61131 VINN.n364 VINN.n165 4.5005
R61132 VINN.n233 VINN.n165 4.5005
R61133 VINN.n366 VINN.n165 4.5005
R61134 VINN.n232 VINN.n165 4.5005
R61135 VINN.n368 VINN.n165 4.5005
R61136 VINN.n231 VINN.n165 4.5005
R61137 VINN.n370 VINN.n165 4.5005
R61138 VINN.n230 VINN.n165 4.5005
R61139 VINN.n372 VINN.n165 4.5005
R61140 VINN.n229 VINN.n165 4.5005
R61141 VINN.n374 VINN.n165 4.5005
R61142 VINN.n228 VINN.n165 4.5005
R61143 VINN.n376 VINN.n165 4.5005
R61144 VINN.n227 VINN.n165 4.5005
R61145 VINN.n378 VINN.n165 4.5005
R61146 VINN.n226 VINN.n165 4.5005
R61147 VINN.n380 VINN.n165 4.5005
R61148 VINN.n225 VINN.n165 4.5005
R61149 VINN.n382 VINN.n165 4.5005
R61150 VINN.n224 VINN.n165 4.5005
R61151 VINN.n384 VINN.n165 4.5005
R61152 VINN.n223 VINN.n165 4.5005
R61153 VINN.n386 VINN.n165 4.5005
R61154 VINN.n222 VINN.n165 4.5005
R61155 VINN.n388 VINN.n165 4.5005
R61156 VINN.n221 VINN.n165 4.5005
R61157 VINN.n390 VINN.n165 4.5005
R61158 VINN.n220 VINN.n165 4.5005
R61159 VINN.n392 VINN.n165 4.5005
R61160 VINN.n219 VINN.n165 4.5005
R61161 VINN.n394 VINN.n165 4.5005
R61162 VINN.n218 VINN.n165 4.5005
R61163 VINN.n396 VINN.n165 4.5005
R61164 VINN.n217 VINN.n165 4.5005
R61165 VINN.n398 VINN.n165 4.5005
R61166 VINN.n216 VINN.n165 4.5005
R61167 VINN.n400 VINN.n165 4.5005
R61168 VINN.n215 VINN.n165 4.5005
R61169 VINN.n654 VINN.n165 4.5005
R61170 VINN.n656 VINN.n165 4.5005
R61171 VINN.n165 VINN.n0 4.5005
R61172 VINN.n278 VINN.n135 4.5005
R61173 VINN.n276 VINN.n135 4.5005
R61174 VINN.n280 VINN.n135 4.5005
R61175 VINN.n275 VINN.n135 4.5005
R61176 VINN.n282 VINN.n135 4.5005
R61177 VINN.n274 VINN.n135 4.5005
R61178 VINN.n284 VINN.n135 4.5005
R61179 VINN.n273 VINN.n135 4.5005
R61180 VINN.n286 VINN.n135 4.5005
R61181 VINN.n272 VINN.n135 4.5005
R61182 VINN.n288 VINN.n135 4.5005
R61183 VINN.n271 VINN.n135 4.5005
R61184 VINN.n290 VINN.n135 4.5005
R61185 VINN.n270 VINN.n135 4.5005
R61186 VINN.n292 VINN.n135 4.5005
R61187 VINN.n269 VINN.n135 4.5005
R61188 VINN.n294 VINN.n135 4.5005
R61189 VINN.n268 VINN.n135 4.5005
R61190 VINN.n296 VINN.n135 4.5005
R61191 VINN.n267 VINN.n135 4.5005
R61192 VINN.n298 VINN.n135 4.5005
R61193 VINN.n266 VINN.n135 4.5005
R61194 VINN.n300 VINN.n135 4.5005
R61195 VINN.n265 VINN.n135 4.5005
R61196 VINN.n302 VINN.n135 4.5005
R61197 VINN.n264 VINN.n135 4.5005
R61198 VINN.n304 VINN.n135 4.5005
R61199 VINN.n263 VINN.n135 4.5005
R61200 VINN.n306 VINN.n135 4.5005
R61201 VINN.n262 VINN.n135 4.5005
R61202 VINN.n308 VINN.n135 4.5005
R61203 VINN.n261 VINN.n135 4.5005
R61204 VINN.n310 VINN.n135 4.5005
R61205 VINN.n260 VINN.n135 4.5005
R61206 VINN.n312 VINN.n135 4.5005
R61207 VINN.n259 VINN.n135 4.5005
R61208 VINN.n314 VINN.n135 4.5005
R61209 VINN.n258 VINN.n135 4.5005
R61210 VINN.n316 VINN.n135 4.5005
R61211 VINN.n257 VINN.n135 4.5005
R61212 VINN.n318 VINN.n135 4.5005
R61213 VINN.n256 VINN.n135 4.5005
R61214 VINN.n320 VINN.n135 4.5005
R61215 VINN.n255 VINN.n135 4.5005
R61216 VINN.n322 VINN.n135 4.5005
R61217 VINN.n254 VINN.n135 4.5005
R61218 VINN.n324 VINN.n135 4.5005
R61219 VINN.n253 VINN.n135 4.5005
R61220 VINN.n326 VINN.n135 4.5005
R61221 VINN.n252 VINN.n135 4.5005
R61222 VINN.n328 VINN.n135 4.5005
R61223 VINN.n251 VINN.n135 4.5005
R61224 VINN.n330 VINN.n135 4.5005
R61225 VINN.n250 VINN.n135 4.5005
R61226 VINN.n332 VINN.n135 4.5005
R61227 VINN.n249 VINN.n135 4.5005
R61228 VINN.n334 VINN.n135 4.5005
R61229 VINN.n248 VINN.n135 4.5005
R61230 VINN.n336 VINN.n135 4.5005
R61231 VINN.n247 VINN.n135 4.5005
R61232 VINN.n338 VINN.n135 4.5005
R61233 VINN.n246 VINN.n135 4.5005
R61234 VINN.n340 VINN.n135 4.5005
R61235 VINN.n245 VINN.n135 4.5005
R61236 VINN.n342 VINN.n135 4.5005
R61237 VINN.n244 VINN.n135 4.5005
R61238 VINN.n344 VINN.n135 4.5005
R61239 VINN.n243 VINN.n135 4.5005
R61240 VINN.n346 VINN.n135 4.5005
R61241 VINN.n242 VINN.n135 4.5005
R61242 VINN.n348 VINN.n135 4.5005
R61243 VINN.n241 VINN.n135 4.5005
R61244 VINN.n350 VINN.n135 4.5005
R61245 VINN.n240 VINN.n135 4.5005
R61246 VINN.n352 VINN.n135 4.5005
R61247 VINN.n239 VINN.n135 4.5005
R61248 VINN.n354 VINN.n135 4.5005
R61249 VINN.n238 VINN.n135 4.5005
R61250 VINN.n356 VINN.n135 4.5005
R61251 VINN.n237 VINN.n135 4.5005
R61252 VINN.n358 VINN.n135 4.5005
R61253 VINN.n236 VINN.n135 4.5005
R61254 VINN.n360 VINN.n135 4.5005
R61255 VINN.n235 VINN.n135 4.5005
R61256 VINN.n362 VINN.n135 4.5005
R61257 VINN.n234 VINN.n135 4.5005
R61258 VINN.n364 VINN.n135 4.5005
R61259 VINN.n233 VINN.n135 4.5005
R61260 VINN.n366 VINN.n135 4.5005
R61261 VINN.n232 VINN.n135 4.5005
R61262 VINN.n368 VINN.n135 4.5005
R61263 VINN.n231 VINN.n135 4.5005
R61264 VINN.n370 VINN.n135 4.5005
R61265 VINN.n230 VINN.n135 4.5005
R61266 VINN.n372 VINN.n135 4.5005
R61267 VINN.n229 VINN.n135 4.5005
R61268 VINN.n374 VINN.n135 4.5005
R61269 VINN.n228 VINN.n135 4.5005
R61270 VINN.n376 VINN.n135 4.5005
R61271 VINN.n227 VINN.n135 4.5005
R61272 VINN.n378 VINN.n135 4.5005
R61273 VINN.n226 VINN.n135 4.5005
R61274 VINN.n380 VINN.n135 4.5005
R61275 VINN.n225 VINN.n135 4.5005
R61276 VINN.n382 VINN.n135 4.5005
R61277 VINN.n224 VINN.n135 4.5005
R61278 VINN.n384 VINN.n135 4.5005
R61279 VINN.n223 VINN.n135 4.5005
R61280 VINN.n386 VINN.n135 4.5005
R61281 VINN.n222 VINN.n135 4.5005
R61282 VINN.n388 VINN.n135 4.5005
R61283 VINN.n221 VINN.n135 4.5005
R61284 VINN.n390 VINN.n135 4.5005
R61285 VINN.n220 VINN.n135 4.5005
R61286 VINN.n392 VINN.n135 4.5005
R61287 VINN.n219 VINN.n135 4.5005
R61288 VINN.n394 VINN.n135 4.5005
R61289 VINN.n218 VINN.n135 4.5005
R61290 VINN.n396 VINN.n135 4.5005
R61291 VINN.n217 VINN.n135 4.5005
R61292 VINN.n398 VINN.n135 4.5005
R61293 VINN.n216 VINN.n135 4.5005
R61294 VINN.n400 VINN.n135 4.5005
R61295 VINN.n215 VINN.n135 4.5005
R61296 VINN.n654 VINN.n135 4.5005
R61297 VINN.n656 VINN.n135 4.5005
R61298 VINN.n135 VINN.n0 4.5005
R61299 VINN.n278 VINN.n166 4.5005
R61300 VINN.n276 VINN.n166 4.5005
R61301 VINN.n280 VINN.n166 4.5005
R61302 VINN.n275 VINN.n166 4.5005
R61303 VINN.n282 VINN.n166 4.5005
R61304 VINN.n274 VINN.n166 4.5005
R61305 VINN.n284 VINN.n166 4.5005
R61306 VINN.n273 VINN.n166 4.5005
R61307 VINN.n286 VINN.n166 4.5005
R61308 VINN.n272 VINN.n166 4.5005
R61309 VINN.n288 VINN.n166 4.5005
R61310 VINN.n271 VINN.n166 4.5005
R61311 VINN.n290 VINN.n166 4.5005
R61312 VINN.n270 VINN.n166 4.5005
R61313 VINN.n292 VINN.n166 4.5005
R61314 VINN.n269 VINN.n166 4.5005
R61315 VINN.n294 VINN.n166 4.5005
R61316 VINN.n268 VINN.n166 4.5005
R61317 VINN.n296 VINN.n166 4.5005
R61318 VINN.n267 VINN.n166 4.5005
R61319 VINN.n298 VINN.n166 4.5005
R61320 VINN.n266 VINN.n166 4.5005
R61321 VINN.n300 VINN.n166 4.5005
R61322 VINN.n265 VINN.n166 4.5005
R61323 VINN.n302 VINN.n166 4.5005
R61324 VINN.n264 VINN.n166 4.5005
R61325 VINN.n304 VINN.n166 4.5005
R61326 VINN.n263 VINN.n166 4.5005
R61327 VINN.n306 VINN.n166 4.5005
R61328 VINN.n262 VINN.n166 4.5005
R61329 VINN.n308 VINN.n166 4.5005
R61330 VINN.n261 VINN.n166 4.5005
R61331 VINN.n310 VINN.n166 4.5005
R61332 VINN.n260 VINN.n166 4.5005
R61333 VINN.n312 VINN.n166 4.5005
R61334 VINN.n259 VINN.n166 4.5005
R61335 VINN.n314 VINN.n166 4.5005
R61336 VINN.n258 VINN.n166 4.5005
R61337 VINN.n316 VINN.n166 4.5005
R61338 VINN.n257 VINN.n166 4.5005
R61339 VINN.n318 VINN.n166 4.5005
R61340 VINN.n256 VINN.n166 4.5005
R61341 VINN.n320 VINN.n166 4.5005
R61342 VINN.n255 VINN.n166 4.5005
R61343 VINN.n322 VINN.n166 4.5005
R61344 VINN.n254 VINN.n166 4.5005
R61345 VINN.n324 VINN.n166 4.5005
R61346 VINN.n253 VINN.n166 4.5005
R61347 VINN.n326 VINN.n166 4.5005
R61348 VINN.n252 VINN.n166 4.5005
R61349 VINN.n328 VINN.n166 4.5005
R61350 VINN.n251 VINN.n166 4.5005
R61351 VINN.n330 VINN.n166 4.5005
R61352 VINN.n250 VINN.n166 4.5005
R61353 VINN.n332 VINN.n166 4.5005
R61354 VINN.n249 VINN.n166 4.5005
R61355 VINN.n334 VINN.n166 4.5005
R61356 VINN.n248 VINN.n166 4.5005
R61357 VINN.n336 VINN.n166 4.5005
R61358 VINN.n247 VINN.n166 4.5005
R61359 VINN.n338 VINN.n166 4.5005
R61360 VINN.n246 VINN.n166 4.5005
R61361 VINN.n340 VINN.n166 4.5005
R61362 VINN.n245 VINN.n166 4.5005
R61363 VINN.n342 VINN.n166 4.5005
R61364 VINN.n244 VINN.n166 4.5005
R61365 VINN.n344 VINN.n166 4.5005
R61366 VINN.n243 VINN.n166 4.5005
R61367 VINN.n346 VINN.n166 4.5005
R61368 VINN.n242 VINN.n166 4.5005
R61369 VINN.n348 VINN.n166 4.5005
R61370 VINN.n241 VINN.n166 4.5005
R61371 VINN.n350 VINN.n166 4.5005
R61372 VINN.n240 VINN.n166 4.5005
R61373 VINN.n352 VINN.n166 4.5005
R61374 VINN.n239 VINN.n166 4.5005
R61375 VINN.n354 VINN.n166 4.5005
R61376 VINN.n238 VINN.n166 4.5005
R61377 VINN.n356 VINN.n166 4.5005
R61378 VINN.n237 VINN.n166 4.5005
R61379 VINN.n358 VINN.n166 4.5005
R61380 VINN.n236 VINN.n166 4.5005
R61381 VINN.n360 VINN.n166 4.5005
R61382 VINN.n235 VINN.n166 4.5005
R61383 VINN.n362 VINN.n166 4.5005
R61384 VINN.n234 VINN.n166 4.5005
R61385 VINN.n364 VINN.n166 4.5005
R61386 VINN.n233 VINN.n166 4.5005
R61387 VINN.n366 VINN.n166 4.5005
R61388 VINN.n232 VINN.n166 4.5005
R61389 VINN.n368 VINN.n166 4.5005
R61390 VINN.n231 VINN.n166 4.5005
R61391 VINN.n370 VINN.n166 4.5005
R61392 VINN.n230 VINN.n166 4.5005
R61393 VINN.n372 VINN.n166 4.5005
R61394 VINN.n229 VINN.n166 4.5005
R61395 VINN.n374 VINN.n166 4.5005
R61396 VINN.n228 VINN.n166 4.5005
R61397 VINN.n376 VINN.n166 4.5005
R61398 VINN.n227 VINN.n166 4.5005
R61399 VINN.n378 VINN.n166 4.5005
R61400 VINN.n226 VINN.n166 4.5005
R61401 VINN.n380 VINN.n166 4.5005
R61402 VINN.n225 VINN.n166 4.5005
R61403 VINN.n382 VINN.n166 4.5005
R61404 VINN.n224 VINN.n166 4.5005
R61405 VINN.n384 VINN.n166 4.5005
R61406 VINN.n223 VINN.n166 4.5005
R61407 VINN.n386 VINN.n166 4.5005
R61408 VINN.n222 VINN.n166 4.5005
R61409 VINN.n388 VINN.n166 4.5005
R61410 VINN.n221 VINN.n166 4.5005
R61411 VINN.n390 VINN.n166 4.5005
R61412 VINN.n220 VINN.n166 4.5005
R61413 VINN.n392 VINN.n166 4.5005
R61414 VINN.n219 VINN.n166 4.5005
R61415 VINN.n394 VINN.n166 4.5005
R61416 VINN.n218 VINN.n166 4.5005
R61417 VINN.n396 VINN.n166 4.5005
R61418 VINN.n217 VINN.n166 4.5005
R61419 VINN.n398 VINN.n166 4.5005
R61420 VINN.n216 VINN.n166 4.5005
R61421 VINN.n400 VINN.n166 4.5005
R61422 VINN.n215 VINN.n166 4.5005
R61423 VINN.n654 VINN.n166 4.5005
R61424 VINN.n656 VINN.n166 4.5005
R61425 VINN.n166 VINN.n0 4.5005
R61426 VINN.n278 VINN.n134 4.5005
R61427 VINN.n276 VINN.n134 4.5005
R61428 VINN.n280 VINN.n134 4.5005
R61429 VINN.n275 VINN.n134 4.5005
R61430 VINN.n282 VINN.n134 4.5005
R61431 VINN.n274 VINN.n134 4.5005
R61432 VINN.n284 VINN.n134 4.5005
R61433 VINN.n273 VINN.n134 4.5005
R61434 VINN.n286 VINN.n134 4.5005
R61435 VINN.n272 VINN.n134 4.5005
R61436 VINN.n288 VINN.n134 4.5005
R61437 VINN.n271 VINN.n134 4.5005
R61438 VINN.n290 VINN.n134 4.5005
R61439 VINN.n270 VINN.n134 4.5005
R61440 VINN.n292 VINN.n134 4.5005
R61441 VINN.n269 VINN.n134 4.5005
R61442 VINN.n294 VINN.n134 4.5005
R61443 VINN.n268 VINN.n134 4.5005
R61444 VINN.n296 VINN.n134 4.5005
R61445 VINN.n267 VINN.n134 4.5005
R61446 VINN.n298 VINN.n134 4.5005
R61447 VINN.n266 VINN.n134 4.5005
R61448 VINN.n300 VINN.n134 4.5005
R61449 VINN.n265 VINN.n134 4.5005
R61450 VINN.n302 VINN.n134 4.5005
R61451 VINN.n264 VINN.n134 4.5005
R61452 VINN.n304 VINN.n134 4.5005
R61453 VINN.n263 VINN.n134 4.5005
R61454 VINN.n306 VINN.n134 4.5005
R61455 VINN.n262 VINN.n134 4.5005
R61456 VINN.n308 VINN.n134 4.5005
R61457 VINN.n261 VINN.n134 4.5005
R61458 VINN.n310 VINN.n134 4.5005
R61459 VINN.n260 VINN.n134 4.5005
R61460 VINN.n312 VINN.n134 4.5005
R61461 VINN.n259 VINN.n134 4.5005
R61462 VINN.n314 VINN.n134 4.5005
R61463 VINN.n258 VINN.n134 4.5005
R61464 VINN.n316 VINN.n134 4.5005
R61465 VINN.n257 VINN.n134 4.5005
R61466 VINN.n318 VINN.n134 4.5005
R61467 VINN.n256 VINN.n134 4.5005
R61468 VINN.n320 VINN.n134 4.5005
R61469 VINN.n255 VINN.n134 4.5005
R61470 VINN.n322 VINN.n134 4.5005
R61471 VINN.n254 VINN.n134 4.5005
R61472 VINN.n324 VINN.n134 4.5005
R61473 VINN.n253 VINN.n134 4.5005
R61474 VINN.n326 VINN.n134 4.5005
R61475 VINN.n252 VINN.n134 4.5005
R61476 VINN.n328 VINN.n134 4.5005
R61477 VINN.n251 VINN.n134 4.5005
R61478 VINN.n330 VINN.n134 4.5005
R61479 VINN.n250 VINN.n134 4.5005
R61480 VINN.n332 VINN.n134 4.5005
R61481 VINN.n249 VINN.n134 4.5005
R61482 VINN.n334 VINN.n134 4.5005
R61483 VINN.n248 VINN.n134 4.5005
R61484 VINN.n336 VINN.n134 4.5005
R61485 VINN.n247 VINN.n134 4.5005
R61486 VINN.n338 VINN.n134 4.5005
R61487 VINN.n246 VINN.n134 4.5005
R61488 VINN.n340 VINN.n134 4.5005
R61489 VINN.n245 VINN.n134 4.5005
R61490 VINN.n342 VINN.n134 4.5005
R61491 VINN.n244 VINN.n134 4.5005
R61492 VINN.n344 VINN.n134 4.5005
R61493 VINN.n243 VINN.n134 4.5005
R61494 VINN.n346 VINN.n134 4.5005
R61495 VINN.n242 VINN.n134 4.5005
R61496 VINN.n348 VINN.n134 4.5005
R61497 VINN.n241 VINN.n134 4.5005
R61498 VINN.n350 VINN.n134 4.5005
R61499 VINN.n240 VINN.n134 4.5005
R61500 VINN.n352 VINN.n134 4.5005
R61501 VINN.n239 VINN.n134 4.5005
R61502 VINN.n354 VINN.n134 4.5005
R61503 VINN.n238 VINN.n134 4.5005
R61504 VINN.n356 VINN.n134 4.5005
R61505 VINN.n237 VINN.n134 4.5005
R61506 VINN.n358 VINN.n134 4.5005
R61507 VINN.n236 VINN.n134 4.5005
R61508 VINN.n360 VINN.n134 4.5005
R61509 VINN.n235 VINN.n134 4.5005
R61510 VINN.n362 VINN.n134 4.5005
R61511 VINN.n234 VINN.n134 4.5005
R61512 VINN.n364 VINN.n134 4.5005
R61513 VINN.n233 VINN.n134 4.5005
R61514 VINN.n366 VINN.n134 4.5005
R61515 VINN.n232 VINN.n134 4.5005
R61516 VINN.n368 VINN.n134 4.5005
R61517 VINN.n231 VINN.n134 4.5005
R61518 VINN.n370 VINN.n134 4.5005
R61519 VINN.n230 VINN.n134 4.5005
R61520 VINN.n372 VINN.n134 4.5005
R61521 VINN.n229 VINN.n134 4.5005
R61522 VINN.n374 VINN.n134 4.5005
R61523 VINN.n228 VINN.n134 4.5005
R61524 VINN.n376 VINN.n134 4.5005
R61525 VINN.n227 VINN.n134 4.5005
R61526 VINN.n378 VINN.n134 4.5005
R61527 VINN.n226 VINN.n134 4.5005
R61528 VINN.n380 VINN.n134 4.5005
R61529 VINN.n225 VINN.n134 4.5005
R61530 VINN.n382 VINN.n134 4.5005
R61531 VINN.n224 VINN.n134 4.5005
R61532 VINN.n384 VINN.n134 4.5005
R61533 VINN.n223 VINN.n134 4.5005
R61534 VINN.n386 VINN.n134 4.5005
R61535 VINN.n222 VINN.n134 4.5005
R61536 VINN.n388 VINN.n134 4.5005
R61537 VINN.n221 VINN.n134 4.5005
R61538 VINN.n390 VINN.n134 4.5005
R61539 VINN.n220 VINN.n134 4.5005
R61540 VINN.n392 VINN.n134 4.5005
R61541 VINN.n219 VINN.n134 4.5005
R61542 VINN.n394 VINN.n134 4.5005
R61543 VINN.n218 VINN.n134 4.5005
R61544 VINN.n396 VINN.n134 4.5005
R61545 VINN.n217 VINN.n134 4.5005
R61546 VINN.n398 VINN.n134 4.5005
R61547 VINN.n216 VINN.n134 4.5005
R61548 VINN.n400 VINN.n134 4.5005
R61549 VINN.n215 VINN.n134 4.5005
R61550 VINN.n654 VINN.n134 4.5005
R61551 VINN.n656 VINN.n134 4.5005
R61552 VINN.n134 VINN.n0 4.5005
R61553 VINN.n278 VINN.n167 4.5005
R61554 VINN.n276 VINN.n167 4.5005
R61555 VINN.n280 VINN.n167 4.5005
R61556 VINN.n275 VINN.n167 4.5005
R61557 VINN.n282 VINN.n167 4.5005
R61558 VINN.n274 VINN.n167 4.5005
R61559 VINN.n284 VINN.n167 4.5005
R61560 VINN.n273 VINN.n167 4.5005
R61561 VINN.n286 VINN.n167 4.5005
R61562 VINN.n272 VINN.n167 4.5005
R61563 VINN.n288 VINN.n167 4.5005
R61564 VINN.n271 VINN.n167 4.5005
R61565 VINN.n290 VINN.n167 4.5005
R61566 VINN.n270 VINN.n167 4.5005
R61567 VINN.n292 VINN.n167 4.5005
R61568 VINN.n269 VINN.n167 4.5005
R61569 VINN.n294 VINN.n167 4.5005
R61570 VINN.n268 VINN.n167 4.5005
R61571 VINN.n296 VINN.n167 4.5005
R61572 VINN.n267 VINN.n167 4.5005
R61573 VINN.n298 VINN.n167 4.5005
R61574 VINN.n266 VINN.n167 4.5005
R61575 VINN.n300 VINN.n167 4.5005
R61576 VINN.n265 VINN.n167 4.5005
R61577 VINN.n302 VINN.n167 4.5005
R61578 VINN.n264 VINN.n167 4.5005
R61579 VINN.n304 VINN.n167 4.5005
R61580 VINN.n263 VINN.n167 4.5005
R61581 VINN.n306 VINN.n167 4.5005
R61582 VINN.n262 VINN.n167 4.5005
R61583 VINN.n308 VINN.n167 4.5005
R61584 VINN.n261 VINN.n167 4.5005
R61585 VINN.n310 VINN.n167 4.5005
R61586 VINN.n260 VINN.n167 4.5005
R61587 VINN.n312 VINN.n167 4.5005
R61588 VINN.n259 VINN.n167 4.5005
R61589 VINN.n314 VINN.n167 4.5005
R61590 VINN.n258 VINN.n167 4.5005
R61591 VINN.n316 VINN.n167 4.5005
R61592 VINN.n257 VINN.n167 4.5005
R61593 VINN.n318 VINN.n167 4.5005
R61594 VINN.n256 VINN.n167 4.5005
R61595 VINN.n320 VINN.n167 4.5005
R61596 VINN.n255 VINN.n167 4.5005
R61597 VINN.n322 VINN.n167 4.5005
R61598 VINN.n254 VINN.n167 4.5005
R61599 VINN.n324 VINN.n167 4.5005
R61600 VINN.n253 VINN.n167 4.5005
R61601 VINN.n326 VINN.n167 4.5005
R61602 VINN.n252 VINN.n167 4.5005
R61603 VINN.n328 VINN.n167 4.5005
R61604 VINN.n251 VINN.n167 4.5005
R61605 VINN.n330 VINN.n167 4.5005
R61606 VINN.n250 VINN.n167 4.5005
R61607 VINN.n332 VINN.n167 4.5005
R61608 VINN.n249 VINN.n167 4.5005
R61609 VINN.n334 VINN.n167 4.5005
R61610 VINN.n248 VINN.n167 4.5005
R61611 VINN.n336 VINN.n167 4.5005
R61612 VINN.n247 VINN.n167 4.5005
R61613 VINN.n338 VINN.n167 4.5005
R61614 VINN.n246 VINN.n167 4.5005
R61615 VINN.n340 VINN.n167 4.5005
R61616 VINN.n245 VINN.n167 4.5005
R61617 VINN.n342 VINN.n167 4.5005
R61618 VINN.n244 VINN.n167 4.5005
R61619 VINN.n344 VINN.n167 4.5005
R61620 VINN.n243 VINN.n167 4.5005
R61621 VINN.n346 VINN.n167 4.5005
R61622 VINN.n242 VINN.n167 4.5005
R61623 VINN.n348 VINN.n167 4.5005
R61624 VINN.n241 VINN.n167 4.5005
R61625 VINN.n350 VINN.n167 4.5005
R61626 VINN.n240 VINN.n167 4.5005
R61627 VINN.n352 VINN.n167 4.5005
R61628 VINN.n239 VINN.n167 4.5005
R61629 VINN.n354 VINN.n167 4.5005
R61630 VINN.n238 VINN.n167 4.5005
R61631 VINN.n356 VINN.n167 4.5005
R61632 VINN.n237 VINN.n167 4.5005
R61633 VINN.n358 VINN.n167 4.5005
R61634 VINN.n236 VINN.n167 4.5005
R61635 VINN.n360 VINN.n167 4.5005
R61636 VINN.n235 VINN.n167 4.5005
R61637 VINN.n362 VINN.n167 4.5005
R61638 VINN.n234 VINN.n167 4.5005
R61639 VINN.n364 VINN.n167 4.5005
R61640 VINN.n233 VINN.n167 4.5005
R61641 VINN.n366 VINN.n167 4.5005
R61642 VINN.n232 VINN.n167 4.5005
R61643 VINN.n368 VINN.n167 4.5005
R61644 VINN.n231 VINN.n167 4.5005
R61645 VINN.n370 VINN.n167 4.5005
R61646 VINN.n230 VINN.n167 4.5005
R61647 VINN.n372 VINN.n167 4.5005
R61648 VINN.n229 VINN.n167 4.5005
R61649 VINN.n374 VINN.n167 4.5005
R61650 VINN.n228 VINN.n167 4.5005
R61651 VINN.n376 VINN.n167 4.5005
R61652 VINN.n227 VINN.n167 4.5005
R61653 VINN.n378 VINN.n167 4.5005
R61654 VINN.n226 VINN.n167 4.5005
R61655 VINN.n380 VINN.n167 4.5005
R61656 VINN.n225 VINN.n167 4.5005
R61657 VINN.n382 VINN.n167 4.5005
R61658 VINN.n224 VINN.n167 4.5005
R61659 VINN.n384 VINN.n167 4.5005
R61660 VINN.n223 VINN.n167 4.5005
R61661 VINN.n386 VINN.n167 4.5005
R61662 VINN.n222 VINN.n167 4.5005
R61663 VINN.n388 VINN.n167 4.5005
R61664 VINN.n221 VINN.n167 4.5005
R61665 VINN.n390 VINN.n167 4.5005
R61666 VINN.n220 VINN.n167 4.5005
R61667 VINN.n392 VINN.n167 4.5005
R61668 VINN.n219 VINN.n167 4.5005
R61669 VINN.n394 VINN.n167 4.5005
R61670 VINN.n218 VINN.n167 4.5005
R61671 VINN.n396 VINN.n167 4.5005
R61672 VINN.n217 VINN.n167 4.5005
R61673 VINN.n398 VINN.n167 4.5005
R61674 VINN.n216 VINN.n167 4.5005
R61675 VINN.n400 VINN.n167 4.5005
R61676 VINN.n215 VINN.n167 4.5005
R61677 VINN.n654 VINN.n167 4.5005
R61678 VINN.n656 VINN.n167 4.5005
R61679 VINN.n167 VINN.n0 4.5005
R61680 VINN.n278 VINN.n133 4.5005
R61681 VINN.n276 VINN.n133 4.5005
R61682 VINN.n280 VINN.n133 4.5005
R61683 VINN.n275 VINN.n133 4.5005
R61684 VINN.n282 VINN.n133 4.5005
R61685 VINN.n274 VINN.n133 4.5005
R61686 VINN.n284 VINN.n133 4.5005
R61687 VINN.n273 VINN.n133 4.5005
R61688 VINN.n286 VINN.n133 4.5005
R61689 VINN.n272 VINN.n133 4.5005
R61690 VINN.n288 VINN.n133 4.5005
R61691 VINN.n271 VINN.n133 4.5005
R61692 VINN.n290 VINN.n133 4.5005
R61693 VINN.n270 VINN.n133 4.5005
R61694 VINN.n292 VINN.n133 4.5005
R61695 VINN.n269 VINN.n133 4.5005
R61696 VINN.n294 VINN.n133 4.5005
R61697 VINN.n268 VINN.n133 4.5005
R61698 VINN.n296 VINN.n133 4.5005
R61699 VINN.n267 VINN.n133 4.5005
R61700 VINN.n298 VINN.n133 4.5005
R61701 VINN.n266 VINN.n133 4.5005
R61702 VINN.n300 VINN.n133 4.5005
R61703 VINN.n265 VINN.n133 4.5005
R61704 VINN.n302 VINN.n133 4.5005
R61705 VINN.n264 VINN.n133 4.5005
R61706 VINN.n304 VINN.n133 4.5005
R61707 VINN.n263 VINN.n133 4.5005
R61708 VINN.n306 VINN.n133 4.5005
R61709 VINN.n262 VINN.n133 4.5005
R61710 VINN.n308 VINN.n133 4.5005
R61711 VINN.n261 VINN.n133 4.5005
R61712 VINN.n310 VINN.n133 4.5005
R61713 VINN.n260 VINN.n133 4.5005
R61714 VINN.n312 VINN.n133 4.5005
R61715 VINN.n259 VINN.n133 4.5005
R61716 VINN.n314 VINN.n133 4.5005
R61717 VINN.n258 VINN.n133 4.5005
R61718 VINN.n316 VINN.n133 4.5005
R61719 VINN.n257 VINN.n133 4.5005
R61720 VINN.n318 VINN.n133 4.5005
R61721 VINN.n256 VINN.n133 4.5005
R61722 VINN.n320 VINN.n133 4.5005
R61723 VINN.n255 VINN.n133 4.5005
R61724 VINN.n322 VINN.n133 4.5005
R61725 VINN.n254 VINN.n133 4.5005
R61726 VINN.n324 VINN.n133 4.5005
R61727 VINN.n253 VINN.n133 4.5005
R61728 VINN.n326 VINN.n133 4.5005
R61729 VINN.n252 VINN.n133 4.5005
R61730 VINN.n328 VINN.n133 4.5005
R61731 VINN.n251 VINN.n133 4.5005
R61732 VINN.n330 VINN.n133 4.5005
R61733 VINN.n250 VINN.n133 4.5005
R61734 VINN.n332 VINN.n133 4.5005
R61735 VINN.n249 VINN.n133 4.5005
R61736 VINN.n334 VINN.n133 4.5005
R61737 VINN.n248 VINN.n133 4.5005
R61738 VINN.n336 VINN.n133 4.5005
R61739 VINN.n247 VINN.n133 4.5005
R61740 VINN.n338 VINN.n133 4.5005
R61741 VINN.n246 VINN.n133 4.5005
R61742 VINN.n340 VINN.n133 4.5005
R61743 VINN.n245 VINN.n133 4.5005
R61744 VINN.n342 VINN.n133 4.5005
R61745 VINN.n244 VINN.n133 4.5005
R61746 VINN.n344 VINN.n133 4.5005
R61747 VINN.n243 VINN.n133 4.5005
R61748 VINN.n346 VINN.n133 4.5005
R61749 VINN.n242 VINN.n133 4.5005
R61750 VINN.n348 VINN.n133 4.5005
R61751 VINN.n241 VINN.n133 4.5005
R61752 VINN.n350 VINN.n133 4.5005
R61753 VINN.n240 VINN.n133 4.5005
R61754 VINN.n352 VINN.n133 4.5005
R61755 VINN.n239 VINN.n133 4.5005
R61756 VINN.n354 VINN.n133 4.5005
R61757 VINN.n238 VINN.n133 4.5005
R61758 VINN.n356 VINN.n133 4.5005
R61759 VINN.n237 VINN.n133 4.5005
R61760 VINN.n358 VINN.n133 4.5005
R61761 VINN.n236 VINN.n133 4.5005
R61762 VINN.n360 VINN.n133 4.5005
R61763 VINN.n235 VINN.n133 4.5005
R61764 VINN.n362 VINN.n133 4.5005
R61765 VINN.n234 VINN.n133 4.5005
R61766 VINN.n364 VINN.n133 4.5005
R61767 VINN.n233 VINN.n133 4.5005
R61768 VINN.n366 VINN.n133 4.5005
R61769 VINN.n232 VINN.n133 4.5005
R61770 VINN.n368 VINN.n133 4.5005
R61771 VINN.n231 VINN.n133 4.5005
R61772 VINN.n370 VINN.n133 4.5005
R61773 VINN.n230 VINN.n133 4.5005
R61774 VINN.n372 VINN.n133 4.5005
R61775 VINN.n229 VINN.n133 4.5005
R61776 VINN.n374 VINN.n133 4.5005
R61777 VINN.n228 VINN.n133 4.5005
R61778 VINN.n376 VINN.n133 4.5005
R61779 VINN.n227 VINN.n133 4.5005
R61780 VINN.n378 VINN.n133 4.5005
R61781 VINN.n226 VINN.n133 4.5005
R61782 VINN.n380 VINN.n133 4.5005
R61783 VINN.n225 VINN.n133 4.5005
R61784 VINN.n382 VINN.n133 4.5005
R61785 VINN.n224 VINN.n133 4.5005
R61786 VINN.n384 VINN.n133 4.5005
R61787 VINN.n223 VINN.n133 4.5005
R61788 VINN.n386 VINN.n133 4.5005
R61789 VINN.n222 VINN.n133 4.5005
R61790 VINN.n388 VINN.n133 4.5005
R61791 VINN.n221 VINN.n133 4.5005
R61792 VINN.n390 VINN.n133 4.5005
R61793 VINN.n220 VINN.n133 4.5005
R61794 VINN.n392 VINN.n133 4.5005
R61795 VINN.n219 VINN.n133 4.5005
R61796 VINN.n394 VINN.n133 4.5005
R61797 VINN.n218 VINN.n133 4.5005
R61798 VINN.n396 VINN.n133 4.5005
R61799 VINN.n217 VINN.n133 4.5005
R61800 VINN.n398 VINN.n133 4.5005
R61801 VINN.n216 VINN.n133 4.5005
R61802 VINN.n400 VINN.n133 4.5005
R61803 VINN.n215 VINN.n133 4.5005
R61804 VINN.n654 VINN.n133 4.5005
R61805 VINN.n656 VINN.n133 4.5005
R61806 VINN.n133 VINN.n0 4.5005
R61807 VINN.n278 VINN.n168 4.5005
R61808 VINN.n276 VINN.n168 4.5005
R61809 VINN.n280 VINN.n168 4.5005
R61810 VINN.n275 VINN.n168 4.5005
R61811 VINN.n282 VINN.n168 4.5005
R61812 VINN.n274 VINN.n168 4.5005
R61813 VINN.n284 VINN.n168 4.5005
R61814 VINN.n273 VINN.n168 4.5005
R61815 VINN.n286 VINN.n168 4.5005
R61816 VINN.n272 VINN.n168 4.5005
R61817 VINN.n288 VINN.n168 4.5005
R61818 VINN.n271 VINN.n168 4.5005
R61819 VINN.n290 VINN.n168 4.5005
R61820 VINN.n270 VINN.n168 4.5005
R61821 VINN.n292 VINN.n168 4.5005
R61822 VINN.n269 VINN.n168 4.5005
R61823 VINN.n294 VINN.n168 4.5005
R61824 VINN.n268 VINN.n168 4.5005
R61825 VINN.n296 VINN.n168 4.5005
R61826 VINN.n267 VINN.n168 4.5005
R61827 VINN.n298 VINN.n168 4.5005
R61828 VINN.n266 VINN.n168 4.5005
R61829 VINN.n300 VINN.n168 4.5005
R61830 VINN.n265 VINN.n168 4.5005
R61831 VINN.n302 VINN.n168 4.5005
R61832 VINN.n264 VINN.n168 4.5005
R61833 VINN.n304 VINN.n168 4.5005
R61834 VINN.n263 VINN.n168 4.5005
R61835 VINN.n306 VINN.n168 4.5005
R61836 VINN.n262 VINN.n168 4.5005
R61837 VINN.n308 VINN.n168 4.5005
R61838 VINN.n261 VINN.n168 4.5005
R61839 VINN.n310 VINN.n168 4.5005
R61840 VINN.n260 VINN.n168 4.5005
R61841 VINN.n312 VINN.n168 4.5005
R61842 VINN.n259 VINN.n168 4.5005
R61843 VINN.n314 VINN.n168 4.5005
R61844 VINN.n258 VINN.n168 4.5005
R61845 VINN.n316 VINN.n168 4.5005
R61846 VINN.n257 VINN.n168 4.5005
R61847 VINN.n318 VINN.n168 4.5005
R61848 VINN.n256 VINN.n168 4.5005
R61849 VINN.n320 VINN.n168 4.5005
R61850 VINN.n255 VINN.n168 4.5005
R61851 VINN.n322 VINN.n168 4.5005
R61852 VINN.n254 VINN.n168 4.5005
R61853 VINN.n324 VINN.n168 4.5005
R61854 VINN.n253 VINN.n168 4.5005
R61855 VINN.n326 VINN.n168 4.5005
R61856 VINN.n252 VINN.n168 4.5005
R61857 VINN.n328 VINN.n168 4.5005
R61858 VINN.n251 VINN.n168 4.5005
R61859 VINN.n330 VINN.n168 4.5005
R61860 VINN.n250 VINN.n168 4.5005
R61861 VINN.n332 VINN.n168 4.5005
R61862 VINN.n249 VINN.n168 4.5005
R61863 VINN.n334 VINN.n168 4.5005
R61864 VINN.n248 VINN.n168 4.5005
R61865 VINN.n336 VINN.n168 4.5005
R61866 VINN.n247 VINN.n168 4.5005
R61867 VINN.n338 VINN.n168 4.5005
R61868 VINN.n246 VINN.n168 4.5005
R61869 VINN.n340 VINN.n168 4.5005
R61870 VINN.n245 VINN.n168 4.5005
R61871 VINN.n342 VINN.n168 4.5005
R61872 VINN.n244 VINN.n168 4.5005
R61873 VINN.n344 VINN.n168 4.5005
R61874 VINN.n243 VINN.n168 4.5005
R61875 VINN.n346 VINN.n168 4.5005
R61876 VINN.n242 VINN.n168 4.5005
R61877 VINN.n348 VINN.n168 4.5005
R61878 VINN.n241 VINN.n168 4.5005
R61879 VINN.n350 VINN.n168 4.5005
R61880 VINN.n240 VINN.n168 4.5005
R61881 VINN.n352 VINN.n168 4.5005
R61882 VINN.n239 VINN.n168 4.5005
R61883 VINN.n354 VINN.n168 4.5005
R61884 VINN.n238 VINN.n168 4.5005
R61885 VINN.n356 VINN.n168 4.5005
R61886 VINN.n237 VINN.n168 4.5005
R61887 VINN.n358 VINN.n168 4.5005
R61888 VINN.n236 VINN.n168 4.5005
R61889 VINN.n360 VINN.n168 4.5005
R61890 VINN.n235 VINN.n168 4.5005
R61891 VINN.n362 VINN.n168 4.5005
R61892 VINN.n234 VINN.n168 4.5005
R61893 VINN.n364 VINN.n168 4.5005
R61894 VINN.n233 VINN.n168 4.5005
R61895 VINN.n366 VINN.n168 4.5005
R61896 VINN.n232 VINN.n168 4.5005
R61897 VINN.n368 VINN.n168 4.5005
R61898 VINN.n231 VINN.n168 4.5005
R61899 VINN.n370 VINN.n168 4.5005
R61900 VINN.n230 VINN.n168 4.5005
R61901 VINN.n372 VINN.n168 4.5005
R61902 VINN.n229 VINN.n168 4.5005
R61903 VINN.n374 VINN.n168 4.5005
R61904 VINN.n228 VINN.n168 4.5005
R61905 VINN.n376 VINN.n168 4.5005
R61906 VINN.n227 VINN.n168 4.5005
R61907 VINN.n378 VINN.n168 4.5005
R61908 VINN.n226 VINN.n168 4.5005
R61909 VINN.n380 VINN.n168 4.5005
R61910 VINN.n225 VINN.n168 4.5005
R61911 VINN.n382 VINN.n168 4.5005
R61912 VINN.n224 VINN.n168 4.5005
R61913 VINN.n384 VINN.n168 4.5005
R61914 VINN.n223 VINN.n168 4.5005
R61915 VINN.n386 VINN.n168 4.5005
R61916 VINN.n222 VINN.n168 4.5005
R61917 VINN.n388 VINN.n168 4.5005
R61918 VINN.n221 VINN.n168 4.5005
R61919 VINN.n390 VINN.n168 4.5005
R61920 VINN.n220 VINN.n168 4.5005
R61921 VINN.n392 VINN.n168 4.5005
R61922 VINN.n219 VINN.n168 4.5005
R61923 VINN.n394 VINN.n168 4.5005
R61924 VINN.n218 VINN.n168 4.5005
R61925 VINN.n396 VINN.n168 4.5005
R61926 VINN.n217 VINN.n168 4.5005
R61927 VINN.n398 VINN.n168 4.5005
R61928 VINN.n216 VINN.n168 4.5005
R61929 VINN.n400 VINN.n168 4.5005
R61930 VINN.n215 VINN.n168 4.5005
R61931 VINN.n654 VINN.n168 4.5005
R61932 VINN.n656 VINN.n168 4.5005
R61933 VINN.n168 VINN.n0 4.5005
R61934 VINN.n278 VINN.n132 4.5005
R61935 VINN.n276 VINN.n132 4.5005
R61936 VINN.n280 VINN.n132 4.5005
R61937 VINN.n275 VINN.n132 4.5005
R61938 VINN.n282 VINN.n132 4.5005
R61939 VINN.n274 VINN.n132 4.5005
R61940 VINN.n284 VINN.n132 4.5005
R61941 VINN.n273 VINN.n132 4.5005
R61942 VINN.n286 VINN.n132 4.5005
R61943 VINN.n272 VINN.n132 4.5005
R61944 VINN.n288 VINN.n132 4.5005
R61945 VINN.n271 VINN.n132 4.5005
R61946 VINN.n290 VINN.n132 4.5005
R61947 VINN.n270 VINN.n132 4.5005
R61948 VINN.n292 VINN.n132 4.5005
R61949 VINN.n269 VINN.n132 4.5005
R61950 VINN.n294 VINN.n132 4.5005
R61951 VINN.n268 VINN.n132 4.5005
R61952 VINN.n296 VINN.n132 4.5005
R61953 VINN.n267 VINN.n132 4.5005
R61954 VINN.n298 VINN.n132 4.5005
R61955 VINN.n266 VINN.n132 4.5005
R61956 VINN.n300 VINN.n132 4.5005
R61957 VINN.n265 VINN.n132 4.5005
R61958 VINN.n302 VINN.n132 4.5005
R61959 VINN.n264 VINN.n132 4.5005
R61960 VINN.n304 VINN.n132 4.5005
R61961 VINN.n263 VINN.n132 4.5005
R61962 VINN.n306 VINN.n132 4.5005
R61963 VINN.n262 VINN.n132 4.5005
R61964 VINN.n308 VINN.n132 4.5005
R61965 VINN.n261 VINN.n132 4.5005
R61966 VINN.n310 VINN.n132 4.5005
R61967 VINN.n260 VINN.n132 4.5005
R61968 VINN.n312 VINN.n132 4.5005
R61969 VINN.n259 VINN.n132 4.5005
R61970 VINN.n314 VINN.n132 4.5005
R61971 VINN.n258 VINN.n132 4.5005
R61972 VINN.n316 VINN.n132 4.5005
R61973 VINN.n257 VINN.n132 4.5005
R61974 VINN.n318 VINN.n132 4.5005
R61975 VINN.n256 VINN.n132 4.5005
R61976 VINN.n320 VINN.n132 4.5005
R61977 VINN.n255 VINN.n132 4.5005
R61978 VINN.n322 VINN.n132 4.5005
R61979 VINN.n254 VINN.n132 4.5005
R61980 VINN.n324 VINN.n132 4.5005
R61981 VINN.n253 VINN.n132 4.5005
R61982 VINN.n326 VINN.n132 4.5005
R61983 VINN.n252 VINN.n132 4.5005
R61984 VINN.n328 VINN.n132 4.5005
R61985 VINN.n251 VINN.n132 4.5005
R61986 VINN.n330 VINN.n132 4.5005
R61987 VINN.n250 VINN.n132 4.5005
R61988 VINN.n332 VINN.n132 4.5005
R61989 VINN.n249 VINN.n132 4.5005
R61990 VINN.n334 VINN.n132 4.5005
R61991 VINN.n248 VINN.n132 4.5005
R61992 VINN.n336 VINN.n132 4.5005
R61993 VINN.n247 VINN.n132 4.5005
R61994 VINN.n338 VINN.n132 4.5005
R61995 VINN.n246 VINN.n132 4.5005
R61996 VINN.n340 VINN.n132 4.5005
R61997 VINN.n245 VINN.n132 4.5005
R61998 VINN.n342 VINN.n132 4.5005
R61999 VINN.n244 VINN.n132 4.5005
R62000 VINN.n344 VINN.n132 4.5005
R62001 VINN.n243 VINN.n132 4.5005
R62002 VINN.n346 VINN.n132 4.5005
R62003 VINN.n242 VINN.n132 4.5005
R62004 VINN.n348 VINN.n132 4.5005
R62005 VINN.n241 VINN.n132 4.5005
R62006 VINN.n350 VINN.n132 4.5005
R62007 VINN.n240 VINN.n132 4.5005
R62008 VINN.n352 VINN.n132 4.5005
R62009 VINN.n239 VINN.n132 4.5005
R62010 VINN.n354 VINN.n132 4.5005
R62011 VINN.n238 VINN.n132 4.5005
R62012 VINN.n356 VINN.n132 4.5005
R62013 VINN.n237 VINN.n132 4.5005
R62014 VINN.n358 VINN.n132 4.5005
R62015 VINN.n236 VINN.n132 4.5005
R62016 VINN.n360 VINN.n132 4.5005
R62017 VINN.n235 VINN.n132 4.5005
R62018 VINN.n362 VINN.n132 4.5005
R62019 VINN.n234 VINN.n132 4.5005
R62020 VINN.n364 VINN.n132 4.5005
R62021 VINN.n233 VINN.n132 4.5005
R62022 VINN.n366 VINN.n132 4.5005
R62023 VINN.n232 VINN.n132 4.5005
R62024 VINN.n368 VINN.n132 4.5005
R62025 VINN.n231 VINN.n132 4.5005
R62026 VINN.n370 VINN.n132 4.5005
R62027 VINN.n230 VINN.n132 4.5005
R62028 VINN.n372 VINN.n132 4.5005
R62029 VINN.n229 VINN.n132 4.5005
R62030 VINN.n374 VINN.n132 4.5005
R62031 VINN.n228 VINN.n132 4.5005
R62032 VINN.n376 VINN.n132 4.5005
R62033 VINN.n227 VINN.n132 4.5005
R62034 VINN.n378 VINN.n132 4.5005
R62035 VINN.n226 VINN.n132 4.5005
R62036 VINN.n380 VINN.n132 4.5005
R62037 VINN.n225 VINN.n132 4.5005
R62038 VINN.n382 VINN.n132 4.5005
R62039 VINN.n224 VINN.n132 4.5005
R62040 VINN.n384 VINN.n132 4.5005
R62041 VINN.n223 VINN.n132 4.5005
R62042 VINN.n386 VINN.n132 4.5005
R62043 VINN.n222 VINN.n132 4.5005
R62044 VINN.n388 VINN.n132 4.5005
R62045 VINN.n221 VINN.n132 4.5005
R62046 VINN.n390 VINN.n132 4.5005
R62047 VINN.n220 VINN.n132 4.5005
R62048 VINN.n392 VINN.n132 4.5005
R62049 VINN.n219 VINN.n132 4.5005
R62050 VINN.n394 VINN.n132 4.5005
R62051 VINN.n218 VINN.n132 4.5005
R62052 VINN.n396 VINN.n132 4.5005
R62053 VINN.n217 VINN.n132 4.5005
R62054 VINN.n398 VINN.n132 4.5005
R62055 VINN.n216 VINN.n132 4.5005
R62056 VINN.n400 VINN.n132 4.5005
R62057 VINN.n215 VINN.n132 4.5005
R62058 VINN.n654 VINN.n132 4.5005
R62059 VINN.n656 VINN.n132 4.5005
R62060 VINN.n132 VINN.n0 4.5005
R62061 VINN.n278 VINN.n169 4.5005
R62062 VINN.n276 VINN.n169 4.5005
R62063 VINN.n280 VINN.n169 4.5005
R62064 VINN.n275 VINN.n169 4.5005
R62065 VINN.n282 VINN.n169 4.5005
R62066 VINN.n274 VINN.n169 4.5005
R62067 VINN.n284 VINN.n169 4.5005
R62068 VINN.n273 VINN.n169 4.5005
R62069 VINN.n286 VINN.n169 4.5005
R62070 VINN.n272 VINN.n169 4.5005
R62071 VINN.n288 VINN.n169 4.5005
R62072 VINN.n271 VINN.n169 4.5005
R62073 VINN.n290 VINN.n169 4.5005
R62074 VINN.n270 VINN.n169 4.5005
R62075 VINN.n292 VINN.n169 4.5005
R62076 VINN.n269 VINN.n169 4.5005
R62077 VINN.n294 VINN.n169 4.5005
R62078 VINN.n268 VINN.n169 4.5005
R62079 VINN.n296 VINN.n169 4.5005
R62080 VINN.n267 VINN.n169 4.5005
R62081 VINN.n298 VINN.n169 4.5005
R62082 VINN.n266 VINN.n169 4.5005
R62083 VINN.n300 VINN.n169 4.5005
R62084 VINN.n265 VINN.n169 4.5005
R62085 VINN.n302 VINN.n169 4.5005
R62086 VINN.n264 VINN.n169 4.5005
R62087 VINN.n304 VINN.n169 4.5005
R62088 VINN.n263 VINN.n169 4.5005
R62089 VINN.n306 VINN.n169 4.5005
R62090 VINN.n262 VINN.n169 4.5005
R62091 VINN.n308 VINN.n169 4.5005
R62092 VINN.n261 VINN.n169 4.5005
R62093 VINN.n310 VINN.n169 4.5005
R62094 VINN.n260 VINN.n169 4.5005
R62095 VINN.n312 VINN.n169 4.5005
R62096 VINN.n259 VINN.n169 4.5005
R62097 VINN.n314 VINN.n169 4.5005
R62098 VINN.n258 VINN.n169 4.5005
R62099 VINN.n316 VINN.n169 4.5005
R62100 VINN.n257 VINN.n169 4.5005
R62101 VINN.n318 VINN.n169 4.5005
R62102 VINN.n256 VINN.n169 4.5005
R62103 VINN.n320 VINN.n169 4.5005
R62104 VINN.n255 VINN.n169 4.5005
R62105 VINN.n322 VINN.n169 4.5005
R62106 VINN.n254 VINN.n169 4.5005
R62107 VINN.n324 VINN.n169 4.5005
R62108 VINN.n253 VINN.n169 4.5005
R62109 VINN.n326 VINN.n169 4.5005
R62110 VINN.n252 VINN.n169 4.5005
R62111 VINN.n328 VINN.n169 4.5005
R62112 VINN.n251 VINN.n169 4.5005
R62113 VINN.n330 VINN.n169 4.5005
R62114 VINN.n250 VINN.n169 4.5005
R62115 VINN.n332 VINN.n169 4.5005
R62116 VINN.n249 VINN.n169 4.5005
R62117 VINN.n334 VINN.n169 4.5005
R62118 VINN.n248 VINN.n169 4.5005
R62119 VINN.n336 VINN.n169 4.5005
R62120 VINN.n247 VINN.n169 4.5005
R62121 VINN.n338 VINN.n169 4.5005
R62122 VINN.n246 VINN.n169 4.5005
R62123 VINN.n340 VINN.n169 4.5005
R62124 VINN.n245 VINN.n169 4.5005
R62125 VINN.n342 VINN.n169 4.5005
R62126 VINN.n244 VINN.n169 4.5005
R62127 VINN.n344 VINN.n169 4.5005
R62128 VINN.n243 VINN.n169 4.5005
R62129 VINN.n346 VINN.n169 4.5005
R62130 VINN.n242 VINN.n169 4.5005
R62131 VINN.n348 VINN.n169 4.5005
R62132 VINN.n241 VINN.n169 4.5005
R62133 VINN.n350 VINN.n169 4.5005
R62134 VINN.n240 VINN.n169 4.5005
R62135 VINN.n352 VINN.n169 4.5005
R62136 VINN.n239 VINN.n169 4.5005
R62137 VINN.n354 VINN.n169 4.5005
R62138 VINN.n238 VINN.n169 4.5005
R62139 VINN.n356 VINN.n169 4.5005
R62140 VINN.n237 VINN.n169 4.5005
R62141 VINN.n358 VINN.n169 4.5005
R62142 VINN.n236 VINN.n169 4.5005
R62143 VINN.n360 VINN.n169 4.5005
R62144 VINN.n235 VINN.n169 4.5005
R62145 VINN.n362 VINN.n169 4.5005
R62146 VINN.n234 VINN.n169 4.5005
R62147 VINN.n364 VINN.n169 4.5005
R62148 VINN.n233 VINN.n169 4.5005
R62149 VINN.n366 VINN.n169 4.5005
R62150 VINN.n232 VINN.n169 4.5005
R62151 VINN.n368 VINN.n169 4.5005
R62152 VINN.n231 VINN.n169 4.5005
R62153 VINN.n370 VINN.n169 4.5005
R62154 VINN.n230 VINN.n169 4.5005
R62155 VINN.n372 VINN.n169 4.5005
R62156 VINN.n229 VINN.n169 4.5005
R62157 VINN.n374 VINN.n169 4.5005
R62158 VINN.n228 VINN.n169 4.5005
R62159 VINN.n376 VINN.n169 4.5005
R62160 VINN.n227 VINN.n169 4.5005
R62161 VINN.n378 VINN.n169 4.5005
R62162 VINN.n226 VINN.n169 4.5005
R62163 VINN.n380 VINN.n169 4.5005
R62164 VINN.n225 VINN.n169 4.5005
R62165 VINN.n382 VINN.n169 4.5005
R62166 VINN.n224 VINN.n169 4.5005
R62167 VINN.n384 VINN.n169 4.5005
R62168 VINN.n223 VINN.n169 4.5005
R62169 VINN.n386 VINN.n169 4.5005
R62170 VINN.n222 VINN.n169 4.5005
R62171 VINN.n388 VINN.n169 4.5005
R62172 VINN.n221 VINN.n169 4.5005
R62173 VINN.n390 VINN.n169 4.5005
R62174 VINN.n220 VINN.n169 4.5005
R62175 VINN.n392 VINN.n169 4.5005
R62176 VINN.n219 VINN.n169 4.5005
R62177 VINN.n394 VINN.n169 4.5005
R62178 VINN.n218 VINN.n169 4.5005
R62179 VINN.n396 VINN.n169 4.5005
R62180 VINN.n217 VINN.n169 4.5005
R62181 VINN.n398 VINN.n169 4.5005
R62182 VINN.n216 VINN.n169 4.5005
R62183 VINN.n400 VINN.n169 4.5005
R62184 VINN.n215 VINN.n169 4.5005
R62185 VINN.n654 VINN.n169 4.5005
R62186 VINN.n656 VINN.n169 4.5005
R62187 VINN.n169 VINN.n0 4.5005
R62188 VINN.n278 VINN.n131 4.5005
R62189 VINN.n276 VINN.n131 4.5005
R62190 VINN.n280 VINN.n131 4.5005
R62191 VINN.n275 VINN.n131 4.5005
R62192 VINN.n282 VINN.n131 4.5005
R62193 VINN.n274 VINN.n131 4.5005
R62194 VINN.n284 VINN.n131 4.5005
R62195 VINN.n273 VINN.n131 4.5005
R62196 VINN.n286 VINN.n131 4.5005
R62197 VINN.n272 VINN.n131 4.5005
R62198 VINN.n288 VINN.n131 4.5005
R62199 VINN.n271 VINN.n131 4.5005
R62200 VINN.n290 VINN.n131 4.5005
R62201 VINN.n270 VINN.n131 4.5005
R62202 VINN.n292 VINN.n131 4.5005
R62203 VINN.n269 VINN.n131 4.5005
R62204 VINN.n294 VINN.n131 4.5005
R62205 VINN.n268 VINN.n131 4.5005
R62206 VINN.n296 VINN.n131 4.5005
R62207 VINN.n267 VINN.n131 4.5005
R62208 VINN.n298 VINN.n131 4.5005
R62209 VINN.n266 VINN.n131 4.5005
R62210 VINN.n300 VINN.n131 4.5005
R62211 VINN.n265 VINN.n131 4.5005
R62212 VINN.n302 VINN.n131 4.5005
R62213 VINN.n264 VINN.n131 4.5005
R62214 VINN.n304 VINN.n131 4.5005
R62215 VINN.n263 VINN.n131 4.5005
R62216 VINN.n306 VINN.n131 4.5005
R62217 VINN.n262 VINN.n131 4.5005
R62218 VINN.n308 VINN.n131 4.5005
R62219 VINN.n261 VINN.n131 4.5005
R62220 VINN.n310 VINN.n131 4.5005
R62221 VINN.n260 VINN.n131 4.5005
R62222 VINN.n312 VINN.n131 4.5005
R62223 VINN.n259 VINN.n131 4.5005
R62224 VINN.n314 VINN.n131 4.5005
R62225 VINN.n258 VINN.n131 4.5005
R62226 VINN.n316 VINN.n131 4.5005
R62227 VINN.n257 VINN.n131 4.5005
R62228 VINN.n318 VINN.n131 4.5005
R62229 VINN.n256 VINN.n131 4.5005
R62230 VINN.n320 VINN.n131 4.5005
R62231 VINN.n255 VINN.n131 4.5005
R62232 VINN.n322 VINN.n131 4.5005
R62233 VINN.n254 VINN.n131 4.5005
R62234 VINN.n324 VINN.n131 4.5005
R62235 VINN.n253 VINN.n131 4.5005
R62236 VINN.n326 VINN.n131 4.5005
R62237 VINN.n252 VINN.n131 4.5005
R62238 VINN.n328 VINN.n131 4.5005
R62239 VINN.n251 VINN.n131 4.5005
R62240 VINN.n330 VINN.n131 4.5005
R62241 VINN.n250 VINN.n131 4.5005
R62242 VINN.n332 VINN.n131 4.5005
R62243 VINN.n249 VINN.n131 4.5005
R62244 VINN.n334 VINN.n131 4.5005
R62245 VINN.n248 VINN.n131 4.5005
R62246 VINN.n336 VINN.n131 4.5005
R62247 VINN.n247 VINN.n131 4.5005
R62248 VINN.n338 VINN.n131 4.5005
R62249 VINN.n246 VINN.n131 4.5005
R62250 VINN.n340 VINN.n131 4.5005
R62251 VINN.n245 VINN.n131 4.5005
R62252 VINN.n342 VINN.n131 4.5005
R62253 VINN.n244 VINN.n131 4.5005
R62254 VINN.n344 VINN.n131 4.5005
R62255 VINN.n243 VINN.n131 4.5005
R62256 VINN.n346 VINN.n131 4.5005
R62257 VINN.n242 VINN.n131 4.5005
R62258 VINN.n348 VINN.n131 4.5005
R62259 VINN.n241 VINN.n131 4.5005
R62260 VINN.n350 VINN.n131 4.5005
R62261 VINN.n240 VINN.n131 4.5005
R62262 VINN.n352 VINN.n131 4.5005
R62263 VINN.n239 VINN.n131 4.5005
R62264 VINN.n354 VINN.n131 4.5005
R62265 VINN.n238 VINN.n131 4.5005
R62266 VINN.n356 VINN.n131 4.5005
R62267 VINN.n237 VINN.n131 4.5005
R62268 VINN.n358 VINN.n131 4.5005
R62269 VINN.n236 VINN.n131 4.5005
R62270 VINN.n360 VINN.n131 4.5005
R62271 VINN.n235 VINN.n131 4.5005
R62272 VINN.n362 VINN.n131 4.5005
R62273 VINN.n234 VINN.n131 4.5005
R62274 VINN.n364 VINN.n131 4.5005
R62275 VINN.n233 VINN.n131 4.5005
R62276 VINN.n366 VINN.n131 4.5005
R62277 VINN.n232 VINN.n131 4.5005
R62278 VINN.n368 VINN.n131 4.5005
R62279 VINN.n231 VINN.n131 4.5005
R62280 VINN.n370 VINN.n131 4.5005
R62281 VINN.n230 VINN.n131 4.5005
R62282 VINN.n372 VINN.n131 4.5005
R62283 VINN.n229 VINN.n131 4.5005
R62284 VINN.n374 VINN.n131 4.5005
R62285 VINN.n228 VINN.n131 4.5005
R62286 VINN.n376 VINN.n131 4.5005
R62287 VINN.n227 VINN.n131 4.5005
R62288 VINN.n378 VINN.n131 4.5005
R62289 VINN.n226 VINN.n131 4.5005
R62290 VINN.n380 VINN.n131 4.5005
R62291 VINN.n225 VINN.n131 4.5005
R62292 VINN.n382 VINN.n131 4.5005
R62293 VINN.n224 VINN.n131 4.5005
R62294 VINN.n384 VINN.n131 4.5005
R62295 VINN.n223 VINN.n131 4.5005
R62296 VINN.n386 VINN.n131 4.5005
R62297 VINN.n222 VINN.n131 4.5005
R62298 VINN.n388 VINN.n131 4.5005
R62299 VINN.n221 VINN.n131 4.5005
R62300 VINN.n390 VINN.n131 4.5005
R62301 VINN.n220 VINN.n131 4.5005
R62302 VINN.n392 VINN.n131 4.5005
R62303 VINN.n219 VINN.n131 4.5005
R62304 VINN.n394 VINN.n131 4.5005
R62305 VINN.n218 VINN.n131 4.5005
R62306 VINN.n396 VINN.n131 4.5005
R62307 VINN.n217 VINN.n131 4.5005
R62308 VINN.n398 VINN.n131 4.5005
R62309 VINN.n216 VINN.n131 4.5005
R62310 VINN.n400 VINN.n131 4.5005
R62311 VINN.n215 VINN.n131 4.5005
R62312 VINN.n654 VINN.n131 4.5005
R62313 VINN.n656 VINN.n131 4.5005
R62314 VINN.n131 VINN.n0 4.5005
R62315 VINN.n278 VINN.n170 4.5005
R62316 VINN.n276 VINN.n170 4.5005
R62317 VINN.n280 VINN.n170 4.5005
R62318 VINN.n275 VINN.n170 4.5005
R62319 VINN.n282 VINN.n170 4.5005
R62320 VINN.n274 VINN.n170 4.5005
R62321 VINN.n284 VINN.n170 4.5005
R62322 VINN.n273 VINN.n170 4.5005
R62323 VINN.n286 VINN.n170 4.5005
R62324 VINN.n272 VINN.n170 4.5005
R62325 VINN.n288 VINN.n170 4.5005
R62326 VINN.n271 VINN.n170 4.5005
R62327 VINN.n290 VINN.n170 4.5005
R62328 VINN.n270 VINN.n170 4.5005
R62329 VINN.n292 VINN.n170 4.5005
R62330 VINN.n269 VINN.n170 4.5005
R62331 VINN.n294 VINN.n170 4.5005
R62332 VINN.n268 VINN.n170 4.5005
R62333 VINN.n296 VINN.n170 4.5005
R62334 VINN.n267 VINN.n170 4.5005
R62335 VINN.n298 VINN.n170 4.5005
R62336 VINN.n266 VINN.n170 4.5005
R62337 VINN.n300 VINN.n170 4.5005
R62338 VINN.n265 VINN.n170 4.5005
R62339 VINN.n302 VINN.n170 4.5005
R62340 VINN.n264 VINN.n170 4.5005
R62341 VINN.n304 VINN.n170 4.5005
R62342 VINN.n263 VINN.n170 4.5005
R62343 VINN.n306 VINN.n170 4.5005
R62344 VINN.n262 VINN.n170 4.5005
R62345 VINN.n308 VINN.n170 4.5005
R62346 VINN.n261 VINN.n170 4.5005
R62347 VINN.n310 VINN.n170 4.5005
R62348 VINN.n260 VINN.n170 4.5005
R62349 VINN.n312 VINN.n170 4.5005
R62350 VINN.n259 VINN.n170 4.5005
R62351 VINN.n314 VINN.n170 4.5005
R62352 VINN.n258 VINN.n170 4.5005
R62353 VINN.n316 VINN.n170 4.5005
R62354 VINN.n257 VINN.n170 4.5005
R62355 VINN.n318 VINN.n170 4.5005
R62356 VINN.n256 VINN.n170 4.5005
R62357 VINN.n320 VINN.n170 4.5005
R62358 VINN.n255 VINN.n170 4.5005
R62359 VINN.n322 VINN.n170 4.5005
R62360 VINN.n254 VINN.n170 4.5005
R62361 VINN.n324 VINN.n170 4.5005
R62362 VINN.n253 VINN.n170 4.5005
R62363 VINN.n326 VINN.n170 4.5005
R62364 VINN.n252 VINN.n170 4.5005
R62365 VINN.n328 VINN.n170 4.5005
R62366 VINN.n251 VINN.n170 4.5005
R62367 VINN.n330 VINN.n170 4.5005
R62368 VINN.n250 VINN.n170 4.5005
R62369 VINN.n332 VINN.n170 4.5005
R62370 VINN.n249 VINN.n170 4.5005
R62371 VINN.n334 VINN.n170 4.5005
R62372 VINN.n248 VINN.n170 4.5005
R62373 VINN.n336 VINN.n170 4.5005
R62374 VINN.n247 VINN.n170 4.5005
R62375 VINN.n338 VINN.n170 4.5005
R62376 VINN.n246 VINN.n170 4.5005
R62377 VINN.n340 VINN.n170 4.5005
R62378 VINN.n245 VINN.n170 4.5005
R62379 VINN.n342 VINN.n170 4.5005
R62380 VINN.n244 VINN.n170 4.5005
R62381 VINN.n344 VINN.n170 4.5005
R62382 VINN.n243 VINN.n170 4.5005
R62383 VINN.n346 VINN.n170 4.5005
R62384 VINN.n242 VINN.n170 4.5005
R62385 VINN.n348 VINN.n170 4.5005
R62386 VINN.n241 VINN.n170 4.5005
R62387 VINN.n350 VINN.n170 4.5005
R62388 VINN.n240 VINN.n170 4.5005
R62389 VINN.n352 VINN.n170 4.5005
R62390 VINN.n239 VINN.n170 4.5005
R62391 VINN.n354 VINN.n170 4.5005
R62392 VINN.n238 VINN.n170 4.5005
R62393 VINN.n356 VINN.n170 4.5005
R62394 VINN.n237 VINN.n170 4.5005
R62395 VINN.n358 VINN.n170 4.5005
R62396 VINN.n236 VINN.n170 4.5005
R62397 VINN.n360 VINN.n170 4.5005
R62398 VINN.n235 VINN.n170 4.5005
R62399 VINN.n362 VINN.n170 4.5005
R62400 VINN.n234 VINN.n170 4.5005
R62401 VINN.n364 VINN.n170 4.5005
R62402 VINN.n233 VINN.n170 4.5005
R62403 VINN.n366 VINN.n170 4.5005
R62404 VINN.n232 VINN.n170 4.5005
R62405 VINN.n368 VINN.n170 4.5005
R62406 VINN.n231 VINN.n170 4.5005
R62407 VINN.n370 VINN.n170 4.5005
R62408 VINN.n230 VINN.n170 4.5005
R62409 VINN.n372 VINN.n170 4.5005
R62410 VINN.n229 VINN.n170 4.5005
R62411 VINN.n374 VINN.n170 4.5005
R62412 VINN.n228 VINN.n170 4.5005
R62413 VINN.n376 VINN.n170 4.5005
R62414 VINN.n227 VINN.n170 4.5005
R62415 VINN.n378 VINN.n170 4.5005
R62416 VINN.n226 VINN.n170 4.5005
R62417 VINN.n380 VINN.n170 4.5005
R62418 VINN.n225 VINN.n170 4.5005
R62419 VINN.n382 VINN.n170 4.5005
R62420 VINN.n224 VINN.n170 4.5005
R62421 VINN.n384 VINN.n170 4.5005
R62422 VINN.n223 VINN.n170 4.5005
R62423 VINN.n386 VINN.n170 4.5005
R62424 VINN.n222 VINN.n170 4.5005
R62425 VINN.n388 VINN.n170 4.5005
R62426 VINN.n221 VINN.n170 4.5005
R62427 VINN.n390 VINN.n170 4.5005
R62428 VINN.n220 VINN.n170 4.5005
R62429 VINN.n392 VINN.n170 4.5005
R62430 VINN.n219 VINN.n170 4.5005
R62431 VINN.n394 VINN.n170 4.5005
R62432 VINN.n218 VINN.n170 4.5005
R62433 VINN.n396 VINN.n170 4.5005
R62434 VINN.n217 VINN.n170 4.5005
R62435 VINN.n398 VINN.n170 4.5005
R62436 VINN.n216 VINN.n170 4.5005
R62437 VINN.n400 VINN.n170 4.5005
R62438 VINN.n215 VINN.n170 4.5005
R62439 VINN.n654 VINN.n170 4.5005
R62440 VINN.n656 VINN.n170 4.5005
R62441 VINN.n170 VINN.n0 4.5005
R62442 VINN.n278 VINN.n130 4.5005
R62443 VINN.n276 VINN.n130 4.5005
R62444 VINN.n280 VINN.n130 4.5005
R62445 VINN.n275 VINN.n130 4.5005
R62446 VINN.n282 VINN.n130 4.5005
R62447 VINN.n274 VINN.n130 4.5005
R62448 VINN.n284 VINN.n130 4.5005
R62449 VINN.n273 VINN.n130 4.5005
R62450 VINN.n286 VINN.n130 4.5005
R62451 VINN.n272 VINN.n130 4.5005
R62452 VINN.n288 VINN.n130 4.5005
R62453 VINN.n271 VINN.n130 4.5005
R62454 VINN.n290 VINN.n130 4.5005
R62455 VINN.n270 VINN.n130 4.5005
R62456 VINN.n292 VINN.n130 4.5005
R62457 VINN.n269 VINN.n130 4.5005
R62458 VINN.n294 VINN.n130 4.5005
R62459 VINN.n268 VINN.n130 4.5005
R62460 VINN.n296 VINN.n130 4.5005
R62461 VINN.n267 VINN.n130 4.5005
R62462 VINN.n298 VINN.n130 4.5005
R62463 VINN.n266 VINN.n130 4.5005
R62464 VINN.n300 VINN.n130 4.5005
R62465 VINN.n265 VINN.n130 4.5005
R62466 VINN.n302 VINN.n130 4.5005
R62467 VINN.n264 VINN.n130 4.5005
R62468 VINN.n304 VINN.n130 4.5005
R62469 VINN.n263 VINN.n130 4.5005
R62470 VINN.n306 VINN.n130 4.5005
R62471 VINN.n262 VINN.n130 4.5005
R62472 VINN.n308 VINN.n130 4.5005
R62473 VINN.n261 VINN.n130 4.5005
R62474 VINN.n310 VINN.n130 4.5005
R62475 VINN.n260 VINN.n130 4.5005
R62476 VINN.n312 VINN.n130 4.5005
R62477 VINN.n259 VINN.n130 4.5005
R62478 VINN.n314 VINN.n130 4.5005
R62479 VINN.n258 VINN.n130 4.5005
R62480 VINN.n316 VINN.n130 4.5005
R62481 VINN.n257 VINN.n130 4.5005
R62482 VINN.n318 VINN.n130 4.5005
R62483 VINN.n256 VINN.n130 4.5005
R62484 VINN.n320 VINN.n130 4.5005
R62485 VINN.n255 VINN.n130 4.5005
R62486 VINN.n322 VINN.n130 4.5005
R62487 VINN.n254 VINN.n130 4.5005
R62488 VINN.n324 VINN.n130 4.5005
R62489 VINN.n253 VINN.n130 4.5005
R62490 VINN.n326 VINN.n130 4.5005
R62491 VINN.n252 VINN.n130 4.5005
R62492 VINN.n328 VINN.n130 4.5005
R62493 VINN.n251 VINN.n130 4.5005
R62494 VINN.n330 VINN.n130 4.5005
R62495 VINN.n250 VINN.n130 4.5005
R62496 VINN.n332 VINN.n130 4.5005
R62497 VINN.n249 VINN.n130 4.5005
R62498 VINN.n334 VINN.n130 4.5005
R62499 VINN.n248 VINN.n130 4.5005
R62500 VINN.n336 VINN.n130 4.5005
R62501 VINN.n247 VINN.n130 4.5005
R62502 VINN.n338 VINN.n130 4.5005
R62503 VINN.n246 VINN.n130 4.5005
R62504 VINN.n340 VINN.n130 4.5005
R62505 VINN.n245 VINN.n130 4.5005
R62506 VINN.n342 VINN.n130 4.5005
R62507 VINN.n244 VINN.n130 4.5005
R62508 VINN.n344 VINN.n130 4.5005
R62509 VINN.n243 VINN.n130 4.5005
R62510 VINN.n346 VINN.n130 4.5005
R62511 VINN.n242 VINN.n130 4.5005
R62512 VINN.n348 VINN.n130 4.5005
R62513 VINN.n241 VINN.n130 4.5005
R62514 VINN.n350 VINN.n130 4.5005
R62515 VINN.n240 VINN.n130 4.5005
R62516 VINN.n352 VINN.n130 4.5005
R62517 VINN.n239 VINN.n130 4.5005
R62518 VINN.n354 VINN.n130 4.5005
R62519 VINN.n238 VINN.n130 4.5005
R62520 VINN.n356 VINN.n130 4.5005
R62521 VINN.n237 VINN.n130 4.5005
R62522 VINN.n358 VINN.n130 4.5005
R62523 VINN.n236 VINN.n130 4.5005
R62524 VINN.n360 VINN.n130 4.5005
R62525 VINN.n235 VINN.n130 4.5005
R62526 VINN.n362 VINN.n130 4.5005
R62527 VINN.n234 VINN.n130 4.5005
R62528 VINN.n364 VINN.n130 4.5005
R62529 VINN.n233 VINN.n130 4.5005
R62530 VINN.n366 VINN.n130 4.5005
R62531 VINN.n232 VINN.n130 4.5005
R62532 VINN.n368 VINN.n130 4.5005
R62533 VINN.n231 VINN.n130 4.5005
R62534 VINN.n370 VINN.n130 4.5005
R62535 VINN.n230 VINN.n130 4.5005
R62536 VINN.n372 VINN.n130 4.5005
R62537 VINN.n229 VINN.n130 4.5005
R62538 VINN.n374 VINN.n130 4.5005
R62539 VINN.n228 VINN.n130 4.5005
R62540 VINN.n376 VINN.n130 4.5005
R62541 VINN.n227 VINN.n130 4.5005
R62542 VINN.n378 VINN.n130 4.5005
R62543 VINN.n226 VINN.n130 4.5005
R62544 VINN.n380 VINN.n130 4.5005
R62545 VINN.n225 VINN.n130 4.5005
R62546 VINN.n382 VINN.n130 4.5005
R62547 VINN.n224 VINN.n130 4.5005
R62548 VINN.n384 VINN.n130 4.5005
R62549 VINN.n223 VINN.n130 4.5005
R62550 VINN.n386 VINN.n130 4.5005
R62551 VINN.n222 VINN.n130 4.5005
R62552 VINN.n388 VINN.n130 4.5005
R62553 VINN.n221 VINN.n130 4.5005
R62554 VINN.n390 VINN.n130 4.5005
R62555 VINN.n220 VINN.n130 4.5005
R62556 VINN.n392 VINN.n130 4.5005
R62557 VINN.n219 VINN.n130 4.5005
R62558 VINN.n394 VINN.n130 4.5005
R62559 VINN.n218 VINN.n130 4.5005
R62560 VINN.n396 VINN.n130 4.5005
R62561 VINN.n217 VINN.n130 4.5005
R62562 VINN.n398 VINN.n130 4.5005
R62563 VINN.n216 VINN.n130 4.5005
R62564 VINN.n400 VINN.n130 4.5005
R62565 VINN.n215 VINN.n130 4.5005
R62566 VINN.n654 VINN.n130 4.5005
R62567 VINN.n656 VINN.n130 4.5005
R62568 VINN.n130 VINN.n0 4.5005
R62569 VINN.n278 VINN.n171 4.5005
R62570 VINN.n276 VINN.n171 4.5005
R62571 VINN.n280 VINN.n171 4.5005
R62572 VINN.n275 VINN.n171 4.5005
R62573 VINN.n282 VINN.n171 4.5005
R62574 VINN.n274 VINN.n171 4.5005
R62575 VINN.n284 VINN.n171 4.5005
R62576 VINN.n273 VINN.n171 4.5005
R62577 VINN.n286 VINN.n171 4.5005
R62578 VINN.n272 VINN.n171 4.5005
R62579 VINN.n288 VINN.n171 4.5005
R62580 VINN.n271 VINN.n171 4.5005
R62581 VINN.n290 VINN.n171 4.5005
R62582 VINN.n270 VINN.n171 4.5005
R62583 VINN.n292 VINN.n171 4.5005
R62584 VINN.n269 VINN.n171 4.5005
R62585 VINN.n294 VINN.n171 4.5005
R62586 VINN.n268 VINN.n171 4.5005
R62587 VINN.n296 VINN.n171 4.5005
R62588 VINN.n267 VINN.n171 4.5005
R62589 VINN.n298 VINN.n171 4.5005
R62590 VINN.n266 VINN.n171 4.5005
R62591 VINN.n300 VINN.n171 4.5005
R62592 VINN.n265 VINN.n171 4.5005
R62593 VINN.n302 VINN.n171 4.5005
R62594 VINN.n264 VINN.n171 4.5005
R62595 VINN.n304 VINN.n171 4.5005
R62596 VINN.n263 VINN.n171 4.5005
R62597 VINN.n306 VINN.n171 4.5005
R62598 VINN.n262 VINN.n171 4.5005
R62599 VINN.n308 VINN.n171 4.5005
R62600 VINN.n261 VINN.n171 4.5005
R62601 VINN.n310 VINN.n171 4.5005
R62602 VINN.n260 VINN.n171 4.5005
R62603 VINN.n312 VINN.n171 4.5005
R62604 VINN.n259 VINN.n171 4.5005
R62605 VINN.n314 VINN.n171 4.5005
R62606 VINN.n258 VINN.n171 4.5005
R62607 VINN.n316 VINN.n171 4.5005
R62608 VINN.n257 VINN.n171 4.5005
R62609 VINN.n318 VINN.n171 4.5005
R62610 VINN.n256 VINN.n171 4.5005
R62611 VINN.n320 VINN.n171 4.5005
R62612 VINN.n255 VINN.n171 4.5005
R62613 VINN.n322 VINN.n171 4.5005
R62614 VINN.n254 VINN.n171 4.5005
R62615 VINN.n324 VINN.n171 4.5005
R62616 VINN.n253 VINN.n171 4.5005
R62617 VINN.n326 VINN.n171 4.5005
R62618 VINN.n252 VINN.n171 4.5005
R62619 VINN.n328 VINN.n171 4.5005
R62620 VINN.n251 VINN.n171 4.5005
R62621 VINN.n330 VINN.n171 4.5005
R62622 VINN.n250 VINN.n171 4.5005
R62623 VINN.n332 VINN.n171 4.5005
R62624 VINN.n249 VINN.n171 4.5005
R62625 VINN.n334 VINN.n171 4.5005
R62626 VINN.n248 VINN.n171 4.5005
R62627 VINN.n336 VINN.n171 4.5005
R62628 VINN.n247 VINN.n171 4.5005
R62629 VINN.n338 VINN.n171 4.5005
R62630 VINN.n246 VINN.n171 4.5005
R62631 VINN.n340 VINN.n171 4.5005
R62632 VINN.n245 VINN.n171 4.5005
R62633 VINN.n342 VINN.n171 4.5005
R62634 VINN.n244 VINN.n171 4.5005
R62635 VINN.n344 VINN.n171 4.5005
R62636 VINN.n243 VINN.n171 4.5005
R62637 VINN.n346 VINN.n171 4.5005
R62638 VINN.n242 VINN.n171 4.5005
R62639 VINN.n348 VINN.n171 4.5005
R62640 VINN.n241 VINN.n171 4.5005
R62641 VINN.n350 VINN.n171 4.5005
R62642 VINN.n240 VINN.n171 4.5005
R62643 VINN.n352 VINN.n171 4.5005
R62644 VINN.n239 VINN.n171 4.5005
R62645 VINN.n354 VINN.n171 4.5005
R62646 VINN.n238 VINN.n171 4.5005
R62647 VINN.n356 VINN.n171 4.5005
R62648 VINN.n237 VINN.n171 4.5005
R62649 VINN.n358 VINN.n171 4.5005
R62650 VINN.n236 VINN.n171 4.5005
R62651 VINN.n360 VINN.n171 4.5005
R62652 VINN.n235 VINN.n171 4.5005
R62653 VINN.n362 VINN.n171 4.5005
R62654 VINN.n234 VINN.n171 4.5005
R62655 VINN.n364 VINN.n171 4.5005
R62656 VINN.n233 VINN.n171 4.5005
R62657 VINN.n366 VINN.n171 4.5005
R62658 VINN.n232 VINN.n171 4.5005
R62659 VINN.n368 VINN.n171 4.5005
R62660 VINN.n231 VINN.n171 4.5005
R62661 VINN.n370 VINN.n171 4.5005
R62662 VINN.n230 VINN.n171 4.5005
R62663 VINN.n372 VINN.n171 4.5005
R62664 VINN.n229 VINN.n171 4.5005
R62665 VINN.n374 VINN.n171 4.5005
R62666 VINN.n228 VINN.n171 4.5005
R62667 VINN.n376 VINN.n171 4.5005
R62668 VINN.n227 VINN.n171 4.5005
R62669 VINN.n378 VINN.n171 4.5005
R62670 VINN.n226 VINN.n171 4.5005
R62671 VINN.n380 VINN.n171 4.5005
R62672 VINN.n225 VINN.n171 4.5005
R62673 VINN.n382 VINN.n171 4.5005
R62674 VINN.n224 VINN.n171 4.5005
R62675 VINN.n384 VINN.n171 4.5005
R62676 VINN.n223 VINN.n171 4.5005
R62677 VINN.n386 VINN.n171 4.5005
R62678 VINN.n222 VINN.n171 4.5005
R62679 VINN.n388 VINN.n171 4.5005
R62680 VINN.n221 VINN.n171 4.5005
R62681 VINN.n390 VINN.n171 4.5005
R62682 VINN.n220 VINN.n171 4.5005
R62683 VINN.n392 VINN.n171 4.5005
R62684 VINN.n219 VINN.n171 4.5005
R62685 VINN.n394 VINN.n171 4.5005
R62686 VINN.n218 VINN.n171 4.5005
R62687 VINN.n396 VINN.n171 4.5005
R62688 VINN.n217 VINN.n171 4.5005
R62689 VINN.n398 VINN.n171 4.5005
R62690 VINN.n216 VINN.n171 4.5005
R62691 VINN.n400 VINN.n171 4.5005
R62692 VINN.n215 VINN.n171 4.5005
R62693 VINN.n654 VINN.n171 4.5005
R62694 VINN.n656 VINN.n171 4.5005
R62695 VINN.n171 VINN.n0 4.5005
R62696 VINN.n278 VINN.n129 4.5005
R62697 VINN.n276 VINN.n129 4.5005
R62698 VINN.n280 VINN.n129 4.5005
R62699 VINN.n275 VINN.n129 4.5005
R62700 VINN.n282 VINN.n129 4.5005
R62701 VINN.n274 VINN.n129 4.5005
R62702 VINN.n284 VINN.n129 4.5005
R62703 VINN.n273 VINN.n129 4.5005
R62704 VINN.n286 VINN.n129 4.5005
R62705 VINN.n272 VINN.n129 4.5005
R62706 VINN.n288 VINN.n129 4.5005
R62707 VINN.n271 VINN.n129 4.5005
R62708 VINN.n290 VINN.n129 4.5005
R62709 VINN.n270 VINN.n129 4.5005
R62710 VINN.n292 VINN.n129 4.5005
R62711 VINN.n269 VINN.n129 4.5005
R62712 VINN.n294 VINN.n129 4.5005
R62713 VINN.n268 VINN.n129 4.5005
R62714 VINN.n296 VINN.n129 4.5005
R62715 VINN.n267 VINN.n129 4.5005
R62716 VINN.n298 VINN.n129 4.5005
R62717 VINN.n266 VINN.n129 4.5005
R62718 VINN.n300 VINN.n129 4.5005
R62719 VINN.n265 VINN.n129 4.5005
R62720 VINN.n302 VINN.n129 4.5005
R62721 VINN.n264 VINN.n129 4.5005
R62722 VINN.n304 VINN.n129 4.5005
R62723 VINN.n263 VINN.n129 4.5005
R62724 VINN.n306 VINN.n129 4.5005
R62725 VINN.n262 VINN.n129 4.5005
R62726 VINN.n308 VINN.n129 4.5005
R62727 VINN.n261 VINN.n129 4.5005
R62728 VINN.n310 VINN.n129 4.5005
R62729 VINN.n260 VINN.n129 4.5005
R62730 VINN.n312 VINN.n129 4.5005
R62731 VINN.n259 VINN.n129 4.5005
R62732 VINN.n314 VINN.n129 4.5005
R62733 VINN.n258 VINN.n129 4.5005
R62734 VINN.n316 VINN.n129 4.5005
R62735 VINN.n257 VINN.n129 4.5005
R62736 VINN.n318 VINN.n129 4.5005
R62737 VINN.n256 VINN.n129 4.5005
R62738 VINN.n320 VINN.n129 4.5005
R62739 VINN.n255 VINN.n129 4.5005
R62740 VINN.n322 VINN.n129 4.5005
R62741 VINN.n254 VINN.n129 4.5005
R62742 VINN.n324 VINN.n129 4.5005
R62743 VINN.n253 VINN.n129 4.5005
R62744 VINN.n326 VINN.n129 4.5005
R62745 VINN.n252 VINN.n129 4.5005
R62746 VINN.n328 VINN.n129 4.5005
R62747 VINN.n251 VINN.n129 4.5005
R62748 VINN.n330 VINN.n129 4.5005
R62749 VINN.n250 VINN.n129 4.5005
R62750 VINN.n332 VINN.n129 4.5005
R62751 VINN.n249 VINN.n129 4.5005
R62752 VINN.n334 VINN.n129 4.5005
R62753 VINN.n248 VINN.n129 4.5005
R62754 VINN.n336 VINN.n129 4.5005
R62755 VINN.n247 VINN.n129 4.5005
R62756 VINN.n338 VINN.n129 4.5005
R62757 VINN.n246 VINN.n129 4.5005
R62758 VINN.n340 VINN.n129 4.5005
R62759 VINN.n245 VINN.n129 4.5005
R62760 VINN.n342 VINN.n129 4.5005
R62761 VINN.n244 VINN.n129 4.5005
R62762 VINN.n344 VINN.n129 4.5005
R62763 VINN.n243 VINN.n129 4.5005
R62764 VINN.n346 VINN.n129 4.5005
R62765 VINN.n242 VINN.n129 4.5005
R62766 VINN.n348 VINN.n129 4.5005
R62767 VINN.n241 VINN.n129 4.5005
R62768 VINN.n350 VINN.n129 4.5005
R62769 VINN.n240 VINN.n129 4.5005
R62770 VINN.n352 VINN.n129 4.5005
R62771 VINN.n239 VINN.n129 4.5005
R62772 VINN.n354 VINN.n129 4.5005
R62773 VINN.n238 VINN.n129 4.5005
R62774 VINN.n356 VINN.n129 4.5005
R62775 VINN.n237 VINN.n129 4.5005
R62776 VINN.n358 VINN.n129 4.5005
R62777 VINN.n236 VINN.n129 4.5005
R62778 VINN.n360 VINN.n129 4.5005
R62779 VINN.n235 VINN.n129 4.5005
R62780 VINN.n362 VINN.n129 4.5005
R62781 VINN.n234 VINN.n129 4.5005
R62782 VINN.n364 VINN.n129 4.5005
R62783 VINN.n233 VINN.n129 4.5005
R62784 VINN.n366 VINN.n129 4.5005
R62785 VINN.n232 VINN.n129 4.5005
R62786 VINN.n368 VINN.n129 4.5005
R62787 VINN.n231 VINN.n129 4.5005
R62788 VINN.n370 VINN.n129 4.5005
R62789 VINN.n230 VINN.n129 4.5005
R62790 VINN.n372 VINN.n129 4.5005
R62791 VINN.n229 VINN.n129 4.5005
R62792 VINN.n374 VINN.n129 4.5005
R62793 VINN.n228 VINN.n129 4.5005
R62794 VINN.n376 VINN.n129 4.5005
R62795 VINN.n227 VINN.n129 4.5005
R62796 VINN.n378 VINN.n129 4.5005
R62797 VINN.n226 VINN.n129 4.5005
R62798 VINN.n380 VINN.n129 4.5005
R62799 VINN.n225 VINN.n129 4.5005
R62800 VINN.n382 VINN.n129 4.5005
R62801 VINN.n224 VINN.n129 4.5005
R62802 VINN.n384 VINN.n129 4.5005
R62803 VINN.n223 VINN.n129 4.5005
R62804 VINN.n386 VINN.n129 4.5005
R62805 VINN.n222 VINN.n129 4.5005
R62806 VINN.n388 VINN.n129 4.5005
R62807 VINN.n221 VINN.n129 4.5005
R62808 VINN.n390 VINN.n129 4.5005
R62809 VINN.n220 VINN.n129 4.5005
R62810 VINN.n392 VINN.n129 4.5005
R62811 VINN.n219 VINN.n129 4.5005
R62812 VINN.n394 VINN.n129 4.5005
R62813 VINN.n218 VINN.n129 4.5005
R62814 VINN.n396 VINN.n129 4.5005
R62815 VINN.n217 VINN.n129 4.5005
R62816 VINN.n398 VINN.n129 4.5005
R62817 VINN.n216 VINN.n129 4.5005
R62818 VINN.n400 VINN.n129 4.5005
R62819 VINN.n215 VINN.n129 4.5005
R62820 VINN.n654 VINN.n129 4.5005
R62821 VINN.n656 VINN.n129 4.5005
R62822 VINN.n129 VINN.n0 4.5005
R62823 VINN.n278 VINN.n172 4.5005
R62824 VINN.n276 VINN.n172 4.5005
R62825 VINN.n280 VINN.n172 4.5005
R62826 VINN.n275 VINN.n172 4.5005
R62827 VINN.n282 VINN.n172 4.5005
R62828 VINN.n274 VINN.n172 4.5005
R62829 VINN.n284 VINN.n172 4.5005
R62830 VINN.n273 VINN.n172 4.5005
R62831 VINN.n286 VINN.n172 4.5005
R62832 VINN.n272 VINN.n172 4.5005
R62833 VINN.n288 VINN.n172 4.5005
R62834 VINN.n271 VINN.n172 4.5005
R62835 VINN.n290 VINN.n172 4.5005
R62836 VINN.n270 VINN.n172 4.5005
R62837 VINN.n292 VINN.n172 4.5005
R62838 VINN.n269 VINN.n172 4.5005
R62839 VINN.n294 VINN.n172 4.5005
R62840 VINN.n268 VINN.n172 4.5005
R62841 VINN.n296 VINN.n172 4.5005
R62842 VINN.n267 VINN.n172 4.5005
R62843 VINN.n298 VINN.n172 4.5005
R62844 VINN.n266 VINN.n172 4.5005
R62845 VINN.n300 VINN.n172 4.5005
R62846 VINN.n265 VINN.n172 4.5005
R62847 VINN.n302 VINN.n172 4.5005
R62848 VINN.n264 VINN.n172 4.5005
R62849 VINN.n304 VINN.n172 4.5005
R62850 VINN.n263 VINN.n172 4.5005
R62851 VINN.n306 VINN.n172 4.5005
R62852 VINN.n262 VINN.n172 4.5005
R62853 VINN.n308 VINN.n172 4.5005
R62854 VINN.n261 VINN.n172 4.5005
R62855 VINN.n310 VINN.n172 4.5005
R62856 VINN.n260 VINN.n172 4.5005
R62857 VINN.n312 VINN.n172 4.5005
R62858 VINN.n259 VINN.n172 4.5005
R62859 VINN.n314 VINN.n172 4.5005
R62860 VINN.n258 VINN.n172 4.5005
R62861 VINN.n316 VINN.n172 4.5005
R62862 VINN.n257 VINN.n172 4.5005
R62863 VINN.n318 VINN.n172 4.5005
R62864 VINN.n256 VINN.n172 4.5005
R62865 VINN.n320 VINN.n172 4.5005
R62866 VINN.n255 VINN.n172 4.5005
R62867 VINN.n322 VINN.n172 4.5005
R62868 VINN.n254 VINN.n172 4.5005
R62869 VINN.n324 VINN.n172 4.5005
R62870 VINN.n253 VINN.n172 4.5005
R62871 VINN.n326 VINN.n172 4.5005
R62872 VINN.n252 VINN.n172 4.5005
R62873 VINN.n328 VINN.n172 4.5005
R62874 VINN.n251 VINN.n172 4.5005
R62875 VINN.n330 VINN.n172 4.5005
R62876 VINN.n250 VINN.n172 4.5005
R62877 VINN.n332 VINN.n172 4.5005
R62878 VINN.n249 VINN.n172 4.5005
R62879 VINN.n334 VINN.n172 4.5005
R62880 VINN.n248 VINN.n172 4.5005
R62881 VINN.n336 VINN.n172 4.5005
R62882 VINN.n247 VINN.n172 4.5005
R62883 VINN.n338 VINN.n172 4.5005
R62884 VINN.n246 VINN.n172 4.5005
R62885 VINN.n340 VINN.n172 4.5005
R62886 VINN.n245 VINN.n172 4.5005
R62887 VINN.n342 VINN.n172 4.5005
R62888 VINN.n244 VINN.n172 4.5005
R62889 VINN.n344 VINN.n172 4.5005
R62890 VINN.n243 VINN.n172 4.5005
R62891 VINN.n346 VINN.n172 4.5005
R62892 VINN.n242 VINN.n172 4.5005
R62893 VINN.n348 VINN.n172 4.5005
R62894 VINN.n241 VINN.n172 4.5005
R62895 VINN.n350 VINN.n172 4.5005
R62896 VINN.n240 VINN.n172 4.5005
R62897 VINN.n352 VINN.n172 4.5005
R62898 VINN.n239 VINN.n172 4.5005
R62899 VINN.n354 VINN.n172 4.5005
R62900 VINN.n238 VINN.n172 4.5005
R62901 VINN.n356 VINN.n172 4.5005
R62902 VINN.n237 VINN.n172 4.5005
R62903 VINN.n358 VINN.n172 4.5005
R62904 VINN.n236 VINN.n172 4.5005
R62905 VINN.n360 VINN.n172 4.5005
R62906 VINN.n235 VINN.n172 4.5005
R62907 VINN.n362 VINN.n172 4.5005
R62908 VINN.n234 VINN.n172 4.5005
R62909 VINN.n364 VINN.n172 4.5005
R62910 VINN.n233 VINN.n172 4.5005
R62911 VINN.n366 VINN.n172 4.5005
R62912 VINN.n232 VINN.n172 4.5005
R62913 VINN.n368 VINN.n172 4.5005
R62914 VINN.n231 VINN.n172 4.5005
R62915 VINN.n370 VINN.n172 4.5005
R62916 VINN.n230 VINN.n172 4.5005
R62917 VINN.n372 VINN.n172 4.5005
R62918 VINN.n229 VINN.n172 4.5005
R62919 VINN.n374 VINN.n172 4.5005
R62920 VINN.n228 VINN.n172 4.5005
R62921 VINN.n376 VINN.n172 4.5005
R62922 VINN.n227 VINN.n172 4.5005
R62923 VINN.n378 VINN.n172 4.5005
R62924 VINN.n226 VINN.n172 4.5005
R62925 VINN.n380 VINN.n172 4.5005
R62926 VINN.n225 VINN.n172 4.5005
R62927 VINN.n382 VINN.n172 4.5005
R62928 VINN.n224 VINN.n172 4.5005
R62929 VINN.n384 VINN.n172 4.5005
R62930 VINN.n223 VINN.n172 4.5005
R62931 VINN.n386 VINN.n172 4.5005
R62932 VINN.n222 VINN.n172 4.5005
R62933 VINN.n388 VINN.n172 4.5005
R62934 VINN.n221 VINN.n172 4.5005
R62935 VINN.n390 VINN.n172 4.5005
R62936 VINN.n220 VINN.n172 4.5005
R62937 VINN.n392 VINN.n172 4.5005
R62938 VINN.n219 VINN.n172 4.5005
R62939 VINN.n394 VINN.n172 4.5005
R62940 VINN.n218 VINN.n172 4.5005
R62941 VINN.n396 VINN.n172 4.5005
R62942 VINN.n217 VINN.n172 4.5005
R62943 VINN.n398 VINN.n172 4.5005
R62944 VINN.n216 VINN.n172 4.5005
R62945 VINN.n400 VINN.n172 4.5005
R62946 VINN.n215 VINN.n172 4.5005
R62947 VINN.n654 VINN.n172 4.5005
R62948 VINN.n656 VINN.n172 4.5005
R62949 VINN.n172 VINN.n0 4.5005
R62950 VINN.n278 VINN.n128 4.5005
R62951 VINN.n276 VINN.n128 4.5005
R62952 VINN.n280 VINN.n128 4.5005
R62953 VINN.n275 VINN.n128 4.5005
R62954 VINN.n282 VINN.n128 4.5005
R62955 VINN.n274 VINN.n128 4.5005
R62956 VINN.n284 VINN.n128 4.5005
R62957 VINN.n273 VINN.n128 4.5005
R62958 VINN.n286 VINN.n128 4.5005
R62959 VINN.n272 VINN.n128 4.5005
R62960 VINN.n288 VINN.n128 4.5005
R62961 VINN.n271 VINN.n128 4.5005
R62962 VINN.n290 VINN.n128 4.5005
R62963 VINN.n270 VINN.n128 4.5005
R62964 VINN.n292 VINN.n128 4.5005
R62965 VINN.n269 VINN.n128 4.5005
R62966 VINN.n294 VINN.n128 4.5005
R62967 VINN.n268 VINN.n128 4.5005
R62968 VINN.n296 VINN.n128 4.5005
R62969 VINN.n267 VINN.n128 4.5005
R62970 VINN.n298 VINN.n128 4.5005
R62971 VINN.n266 VINN.n128 4.5005
R62972 VINN.n300 VINN.n128 4.5005
R62973 VINN.n265 VINN.n128 4.5005
R62974 VINN.n302 VINN.n128 4.5005
R62975 VINN.n264 VINN.n128 4.5005
R62976 VINN.n304 VINN.n128 4.5005
R62977 VINN.n263 VINN.n128 4.5005
R62978 VINN.n306 VINN.n128 4.5005
R62979 VINN.n262 VINN.n128 4.5005
R62980 VINN.n308 VINN.n128 4.5005
R62981 VINN.n261 VINN.n128 4.5005
R62982 VINN.n310 VINN.n128 4.5005
R62983 VINN.n260 VINN.n128 4.5005
R62984 VINN.n312 VINN.n128 4.5005
R62985 VINN.n259 VINN.n128 4.5005
R62986 VINN.n314 VINN.n128 4.5005
R62987 VINN.n258 VINN.n128 4.5005
R62988 VINN.n316 VINN.n128 4.5005
R62989 VINN.n257 VINN.n128 4.5005
R62990 VINN.n318 VINN.n128 4.5005
R62991 VINN.n256 VINN.n128 4.5005
R62992 VINN.n320 VINN.n128 4.5005
R62993 VINN.n255 VINN.n128 4.5005
R62994 VINN.n322 VINN.n128 4.5005
R62995 VINN.n254 VINN.n128 4.5005
R62996 VINN.n324 VINN.n128 4.5005
R62997 VINN.n253 VINN.n128 4.5005
R62998 VINN.n326 VINN.n128 4.5005
R62999 VINN.n252 VINN.n128 4.5005
R63000 VINN.n328 VINN.n128 4.5005
R63001 VINN.n251 VINN.n128 4.5005
R63002 VINN.n330 VINN.n128 4.5005
R63003 VINN.n250 VINN.n128 4.5005
R63004 VINN.n332 VINN.n128 4.5005
R63005 VINN.n249 VINN.n128 4.5005
R63006 VINN.n334 VINN.n128 4.5005
R63007 VINN.n248 VINN.n128 4.5005
R63008 VINN.n336 VINN.n128 4.5005
R63009 VINN.n247 VINN.n128 4.5005
R63010 VINN.n338 VINN.n128 4.5005
R63011 VINN.n246 VINN.n128 4.5005
R63012 VINN.n340 VINN.n128 4.5005
R63013 VINN.n245 VINN.n128 4.5005
R63014 VINN.n342 VINN.n128 4.5005
R63015 VINN.n244 VINN.n128 4.5005
R63016 VINN.n344 VINN.n128 4.5005
R63017 VINN.n243 VINN.n128 4.5005
R63018 VINN.n346 VINN.n128 4.5005
R63019 VINN.n242 VINN.n128 4.5005
R63020 VINN.n348 VINN.n128 4.5005
R63021 VINN.n241 VINN.n128 4.5005
R63022 VINN.n350 VINN.n128 4.5005
R63023 VINN.n240 VINN.n128 4.5005
R63024 VINN.n352 VINN.n128 4.5005
R63025 VINN.n239 VINN.n128 4.5005
R63026 VINN.n354 VINN.n128 4.5005
R63027 VINN.n238 VINN.n128 4.5005
R63028 VINN.n356 VINN.n128 4.5005
R63029 VINN.n237 VINN.n128 4.5005
R63030 VINN.n358 VINN.n128 4.5005
R63031 VINN.n236 VINN.n128 4.5005
R63032 VINN.n360 VINN.n128 4.5005
R63033 VINN.n235 VINN.n128 4.5005
R63034 VINN.n362 VINN.n128 4.5005
R63035 VINN.n234 VINN.n128 4.5005
R63036 VINN.n364 VINN.n128 4.5005
R63037 VINN.n233 VINN.n128 4.5005
R63038 VINN.n366 VINN.n128 4.5005
R63039 VINN.n232 VINN.n128 4.5005
R63040 VINN.n368 VINN.n128 4.5005
R63041 VINN.n231 VINN.n128 4.5005
R63042 VINN.n370 VINN.n128 4.5005
R63043 VINN.n230 VINN.n128 4.5005
R63044 VINN.n372 VINN.n128 4.5005
R63045 VINN.n229 VINN.n128 4.5005
R63046 VINN.n374 VINN.n128 4.5005
R63047 VINN.n228 VINN.n128 4.5005
R63048 VINN.n376 VINN.n128 4.5005
R63049 VINN.n227 VINN.n128 4.5005
R63050 VINN.n378 VINN.n128 4.5005
R63051 VINN.n226 VINN.n128 4.5005
R63052 VINN.n380 VINN.n128 4.5005
R63053 VINN.n225 VINN.n128 4.5005
R63054 VINN.n382 VINN.n128 4.5005
R63055 VINN.n224 VINN.n128 4.5005
R63056 VINN.n384 VINN.n128 4.5005
R63057 VINN.n223 VINN.n128 4.5005
R63058 VINN.n386 VINN.n128 4.5005
R63059 VINN.n222 VINN.n128 4.5005
R63060 VINN.n388 VINN.n128 4.5005
R63061 VINN.n221 VINN.n128 4.5005
R63062 VINN.n390 VINN.n128 4.5005
R63063 VINN.n220 VINN.n128 4.5005
R63064 VINN.n392 VINN.n128 4.5005
R63065 VINN.n219 VINN.n128 4.5005
R63066 VINN.n394 VINN.n128 4.5005
R63067 VINN.n218 VINN.n128 4.5005
R63068 VINN.n396 VINN.n128 4.5005
R63069 VINN.n217 VINN.n128 4.5005
R63070 VINN.n398 VINN.n128 4.5005
R63071 VINN.n216 VINN.n128 4.5005
R63072 VINN.n400 VINN.n128 4.5005
R63073 VINN.n215 VINN.n128 4.5005
R63074 VINN.n654 VINN.n128 4.5005
R63075 VINN.n656 VINN.n128 4.5005
R63076 VINN.n128 VINN.n0 4.5005
R63077 VINN.n278 VINN.n173 4.5005
R63078 VINN.n276 VINN.n173 4.5005
R63079 VINN.n280 VINN.n173 4.5005
R63080 VINN.n275 VINN.n173 4.5005
R63081 VINN.n282 VINN.n173 4.5005
R63082 VINN.n274 VINN.n173 4.5005
R63083 VINN.n284 VINN.n173 4.5005
R63084 VINN.n273 VINN.n173 4.5005
R63085 VINN.n286 VINN.n173 4.5005
R63086 VINN.n272 VINN.n173 4.5005
R63087 VINN.n288 VINN.n173 4.5005
R63088 VINN.n271 VINN.n173 4.5005
R63089 VINN.n290 VINN.n173 4.5005
R63090 VINN.n270 VINN.n173 4.5005
R63091 VINN.n292 VINN.n173 4.5005
R63092 VINN.n269 VINN.n173 4.5005
R63093 VINN.n294 VINN.n173 4.5005
R63094 VINN.n268 VINN.n173 4.5005
R63095 VINN.n296 VINN.n173 4.5005
R63096 VINN.n267 VINN.n173 4.5005
R63097 VINN.n298 VINN.n173 4.5005
R63098 VINN.n266 VINN.n173 4.5005
R63099 VINN.n300 VINN.n173 4.5005
R63100 VINN.n265 VINN.n173 4.5005
R63101 VINN.n302 VINN.n173 4.5005
R63102 VINN.n264 VINN.n173 4.5005
R63103 VINN.n304 VINN.n173 4.5005
R63104 VINN.n263 VINN.n173 4.5005
R63105 VINN.n306 VINN.n173 4.5005
R63106 VINN.n262 VINN.n173 4.5005
R63107 VINN.n308 VINN.n173 4.5005
R63108 VINN.n261 VINN.n173 4.5005
R63109 VINN.n310 VINN.n173 4.5005
R63110 VINN.n260 VINN.n173 4.5005
R63111 VINN.n312 VINN.n173 4.5005
R63112 VINN.n259 VINN.n173 4.5005
R63113 VINN.n314 VINN.n173 4.5005
R63114 VINN.n258 VINN.n173 4.5005
R63115 VINN.n316 VINN.n173 4.5005
R63116 VINN.n257 VINN.n173 4.5005
R63117 VINN.n318 VINN.n173 4.5005
R63118 VINN.n256 VINN.n173 4.5005
R63119 VINN.n320 VINN.n173 4.5005
R63120 VINN.n255 VINN.n173 4.5005
R63121 VINN.n322 VINN.n173 4.5005
R63122 VINN.n254 VINN.n173 4.5005
R63123 VINN.n324 VINN.n173 4.5005
R63124 VINN.n253 VINN.n173 4.5005
R63125 VINN.n326 VINN.n173 4.5005
R63126 VINN.n252 VINN.n173 4.5005
R63127 VINN.n328 VINN.n173 4.5005
R63128 VINN.n251 VINN.n173 4.5005
R63129 VINN.n330 VINN.n173 4.5005
R63130 VINN.n250 VINN.n173 4.5005
R63131 VINN.n332 VINN.n173 4.5005
R63132 VINN.n249 VINN.n173 4.5005
R63133 VINN.n334 VINN.n173 4.5005
R63134 VINN.n248 VINN.n173 4.5005
R63135 VINN.n336 VINN.n173 4.5005
R63136 VINN.n247 VINN.n173 4.5005
R63137 VINN.n338 VINN.n173 4.5005
R63138 VINN.n246 VINN.n173 4.5005
R63139 VINN.n340 VINN.n173 4.5005
R63140 VINN.n245 VINN.n173 4.5005
R63141 VINN.n342 VINN.n173 4.5005
R63142 VINN.n244 VINN.n173 4.5005
R63143 VINN.n344 VINN.n173 4.5005
R63144 VINN.n243 VINN.n173 4.5005
R63145 VINN.n346 VINN.n173 4.5005
R63146 VINN.n242 VINN.n173 4.5005
R63147 VINN.n348 VINN.n173 4.5005
R63148 VINN.n241 VINN.n173 4.5005
R63149 VINN.n350 VINN.n173 4.5005
R63150 VINN.n240 VINN.n173 4.5005
R63151 VINN.n352 VINN.n173 4.5005
R63152 VINN.n239 VINN.n173 4.5005
R63153 VINN.n354 VINN.n173 4.5005
R63154 VINN.n238 VINN.n173 4.5005
R63155 VINN.n356 VINN.n173 4.5005
R63156 VINN.n237 VINN.n173 4.5005
R63157 VINN.n358 VINN.n173 4.5005
R63158 VINN.n236 VINN.n173 4.5005
R63159 VINN.n360 VINN.n173 4.5005
R63160 VINN.n235 VINN.n173 4.5005
R63161 VINN.n362 VINN.n173 4.5005
R63162 VINN.n234 VINN.n173 4.5005
R63163 VINN.n364 VINN.n173 4.5005
R63164 VINN.n233 VINN.n173 4.5005
R63165 VINN.n366 VINN.n173 4.5005
R63166 VINN.n232 VINN.n173 4.5005
R63167 VINN.n368 VINN.n173 4.5005
R63168 VINN.n231 VINN.n173 4.5005
R63169 VINN.n370 VINN.n173 4.5005
R63170 VINN.n230 VINN.n173 4.5005
R63171 VINN.n372 VINN.n173 4.5005
R63172 VINN.n229 VINN.n173 4.5005
R63173 VINN.n374 VINN.n173 4.5005
R63174 VINN.n228 VINN.n173 4.5005
R63175 VINN.n376 VINN.n173 4.5005
R63176 VINN.n227 VINN.n173 4.5005
R63177 VINN.n378 VINN.n173 4.5005
R63178 VINN.n226 VINN.n173 4.5005
R63179 VINN.n380 VINN.n173 4.5005
R63180 VINN.n225 VINN.n173 4.5005
R63181 VINN.n382 VINN.n173 4.5005
R63182 VINN.n224 VINN.n173 4.5005
R63183 VINN.n384 VINN.n173 4.5005
R63184 VINN.n223 VINN.n173 4.5005
R63185 VINN.n386 VINN.n173 4.5005
R63186 VINN.n222 VINN.n173 4.5005
R63187 VINN.n388 VINN.n173 4.5005
R63188 VINN.n221 VINN.n173 4.5005
R63189 VINN.n390 VINN.n173 4.5005
R63190 VINN.n220 VINN.n173 4.5005
R63191 VINN.n392 VINN.n173 4.5005
R63192 VINN.n219 VINN.n173 4.5005
R63193 VINN.n394 VINN.n173 4.5005
R63194 VINN.n218 VINN.n173 4.5005
R63195 VINN.n396 VINN.n173 4.5005
R63196 VINN.n217 VINN.n173 4.5005
R63197 VINN.n398 VINN.n173 4.5005
R63198 VINN.n216 VINN.n173 4.5005
R63199 VINN.n400 VINN.n173 4.5005
R63200 VINN.n215 VINN.n173 4.5005
R63201 VINN.n654 VINN.n173 4.5005
R63202 VINN.n656 VINN.n173 4.5005
R63203 VINN.n173 VINN.n0 4.5005
R63204 VINN.n278 VINN.n127 4.5005
R63205 VINN.n276 VINN.n127 4.5005
R63206 VINN.n280 VINN.n127 4.5005
R63207 VINN.n275 VINN.n127 4.5005
R63208 VINN.n282 VINN.n127 4.5005
R63209 VINN.n274 VINN.n127 4.5005
R63210 VINN.n284 VINN.n127 4.5005
R63211 VINN.n273 VINN.n127 4.5005
R63212 VINN.n286 VINN.n127 4.5005
R63213 VINN.n272 VINN.n127 4.5005
R63214 VINN.n288 VINN.n127 4.5005
R63215 VINN.n271 VINN.n127 4.5005
R63216 VINN.n290 VINN.n127 4.5005
R63217 VINN.n270 VINN.n127 4.5005
R63218 VINN.n292 VINN.n127 4.5005
R63219 VINN.n269 VINN.n127 4.5005
R63220 VINN.n294 VINN.n127 4.5005
R63221 VINN.n268 VINN.n127 4.5005
R63222 VINN.n296 VINN.n127 4.5005
R63223 VINN.n267 VINN.n127 4.5005
R63224 VINN.n298 VINN.n127 4.5005
R63225 VINN.n266 VINN.n127 4.5005
R63226 VINN.n300 VINN.n127 4.5005
R63227 VINN.n265 VINN.n127 4.5005
R63228 VINN.n302 VINN.n127 4.5005
R63229 VINN.n264 VINN.n127 4.5005
R63230 VINN.n304 VINN.n127 4.5005
R63231 VINN.n263 VINN.n127 4.5005
R63232 VINN.n306 VINN.n127 4.5005
R63233 VINN.n262 VINN.n127 4.5005
R63234 VINN.n308 VINN.n127 4.5005
R63235 VINN.n261 VINN.n127 4.5005
R63236 VINN.n310 VINN.n127 4.5005
R63237 VINN.n260 VINN.n127 4.5005
R63238 VINN.n312 VINN.n127 4.5005
R63239 VINN.n259 VINN.n127 4.5005
R63240 VINN.n314 VINN.n127 4.5005
R63241 VINN.n258 VINN.n127 4.5005
R63242 VINN.n316 VINN.n127 4.5005
R63243 VINN.n257 VINN.n127 4.5005
R63244 VINN.n318 VINN.n127 4.5005
R63245 VINN.n256 VINN.n127 4.5005
R63246 VINN.n320 VINN.n127 4.5005
R63247 VINN.n255 VINN.n127 4.5005
R63248 VINN.n322 VINN.n127 4.5005
R63249 VINN.n254 VINN.n127 4.5005
R63250 VINN.n324 VINN.n127 4.5005
R63251 VINN.n253 VINN.n127 4.5005
R63252 VINN.n326 VINN.n127 4.5005
R63253 VINN.n252 VINN.n127 4.5005
R63254 VINN.n328 VINN.n127 4.5005
R63255 VINN.n251 VINN.n127 4.5005
R63256 VINN.n330 VINN.n127 4.5005
R63257 VINN.n250 VINN.n127 4.5005
R63258 VINN.n332 VINN.n127 4.5005
R63259 VINN.n249 VINN.n127 4.5005
R63260 VINN.n334 VINN.n127 4.5005
R63261 VINN.n248 VINN.n127 4.5005
R63262 VINN.n336 VINN.n127 4.5005
R63263 VINN.n247 VINN.n127 4.5005
R63264 VINN.n338 VINN.n127 4.5005
R63265 VINN.n246 VINN.n127 4.5005
R63266 VINN.n340 VINN.n127 4.5005
R63267 VINN.n245 VINN.n127 4.5005
R63268 VINN.n342 VINN.n127 4.5005
R63269 VINN.n244 VINN.n127 4.5005
R63270 VINN.n344 VINN.n127 4.5005
R63271 VINN.n243 VINN.n127 4.5005
R63272 VINN.n346 VINN.n127 4.5005
R63273 VINN.n242 VINN.n127 4.5005
R63274 VINN.n348 VINN.n127 4.5005
R63275 VINN.n241 VINN.n127 4.5005
R63276 VINN.n350 VINN.n127 4.5005
R63277 VINN.n240 VINN.n127 4.5005
R63278 VINN.n352 VINN.n127 4.5005
R63279 VINN.n239 VINN.n127 4.5005
R63280 VINN.n354 VINN.n127 4.5005
R63281 VINN.n238 VINN.n127 4.5005
R63282 VINN.n356 VINN.n127 4.5005
R63283 VINN.n237 VINN.n127 4.5005
R63284 VINN.n358 VINN.n127 4.5005
R63285 VINN.n236 VINN.n127 4.5005
R63286 VINN.n360 VINN.n127 4.5005
R63287 VINN.n235 VINN.n127 4.5005
R63288 VINN.n362 VINN.n127 4.5005
R63289 VINN.n234 VINN.n127 4.5005
R63290 VINN.n364 VINN.n127 4.5005
R63291 VINN.n233 VINN.n127 4.5005
R63292 VINN.n366 VINN.n127 4.5005
R63293 VINN.n232 VINN.n127 4.5005
R63294 VINN.n368 VINN.n127 4.5005
R63295 VINN.n231 VINN.n127 4.5005
R63296 VINN.n370 VINN.n127 4.5005
R63297 VINN.n230 VINN.n127 4.5005
R63298 VINN.n372 VINN.n127 4.5005
R63299 VINN.n229 VINN.n127 4.5005
R63300 VINN.n374 VINN.n127 4.5005
R63301 VINN.n228 VINN.n127 4.5005
R63302 VINN.n376 VINN.n127 4.5005
R63303 VINN.n227 VINN.n127 4.5005
R63304 VINN.n378 VINN.n127 4.5005
R63305 VINN.n226 VINN.n127 4.5005
R63306 VINN.n380 VINN.n127 4.5005
R63307 VINN.n225 VINN.n127 4.5005
R63308 VINN.n382 VINN.n127 4.5005
R63309 VINN.n224 VINN.n127 4.5005
R63310 VINN.n384 VINN.n127 4.5005
R63311 VINN.n223 VINN.n127 4.5005
R63312 VINN.n386 VINN.n127 4.5005
R63313 VINN.n222 VINN.n127 4.5005
R63314 VINN.n388 VINN.n127 4.5005
R63315 VINN.n221 VINN.n127 4.5005
R63316 VINN.n390 VINN.n127 4.5005
R63317 VINN.n220 VINN.n127 4.5005
R63318 VINN.n392 VINN.n127 4.5005
R63319 VINN.n219 VINN.n127 4.5005
R63320 VINN.n394 VINN.n127 4.5005
R63321 VINN.n218 VINN.n127 4.5005
R63322 VINN.n396 VINN.n127 4.5005
R63323 VINN.n217 VINN.n127 4.5005
R63324 VINN.n398 VINN.n127 4.5005
R63325 VINN.n216 VINN.n127 4.5005
R63326 VINN.n400 VINN.n127 4.5005
R63327 VINN.n215 VINN.n127 4.5005
R63328 VINN.n654 VINN.n127 4.5005
R63329 VINN.n656 VINN.n127 4.5005
R63330 VINN.n127 VINN.n0 4.5005
R63331 VINN.n278 VINN.n174 4.5005
R63332 VINN.n276 VINN.n174 4.5005
R63333 VINN.n280 VINN.n174 4.5005
R63334 VINN.n275 VINN.n174 4.5005
R63335 VINN.n282 VINN.n174 4.5005
R63336 VINN.n274 VINN.n174 4.5005
R63337 VINN.n284 VINN.n174 4.5005
R63338 VINN.n273 VINN.n174 4.5005
R63339 VINN.n286 VINN.n174 4.5005
R63340 VINN.n272 VINN.n174 4.5005
R63341 VINN.n288 VINN.n174 4.5005
R63342 VINN.n271 VINN.n174 4.5005
R63343 VINN.n290 VINN.n174 4.5005
R63344 VINN.n270 VINN.n174 4.5005
R63345 VINN.n292 VINN.n174 4.5005
R63346 VINN.n269 VINN.n174 4.5005
R63347 VINN.n294 VINN.n174 4.5005
R63348 VINN.n268 VINN.n174 4.5005
R63349 VINN.n296 VINN.n174 4.5005
R63350 VINN.n267 VINN.n174 4.5005
R63351 VINN.n298 VINN.n174 4.5005
R63352 VINN.n266 VINN.n174 4.5005
R63353 VINN.n300 VINN.n174 4.5005
R63354 VINN.n265 VINN.n174 4.5005
R63355 VINN.n302 VINN.n174 4.5005
R63356 VINN.n264 VINN.n174 4.5005
R63357 VINN.n304 VINN.n174 4.5005
R63358 VINN.n263 VINN.n174 4.5005
R63359 VINN.n306 VINN.n174 4.5005
R63360 VINN.n262 VINN.n174 4.5005
R63361 VINN.n308 VINN.n174 4.5005
R63362 VINN.n261 VINN.n174 4.5005
R63363 VINN.n310 VINN.n174 4.5005
R63364 VINN.n260 VINN.n174 4.5005
R63365 VINN.n312 VINN.n174 4.5005
R63366 VINN.n259 VINN.n174 4.5005
R63367 VINN.n314 VINN.n174 4.5005
R63368 VINN.n258 VINN.n174 4.5005
R63369 VINN.n316 VINN.n174 4.5005
R63370 VINN.n257 VINN.n174 4.5005
R63371 VINN.n318 VINN.n174 4.5005
R63372 VINN.n256 VINN.n174 4.5005
R63373 VINN.n320 VINN.n174 4.5005
R63374 VINN.n255 VINN.n174 4.5005
R63375 VINN.n322 VINN.n174 4.5005
R63376 VINN.n254 VINN.n174 4.5005
R63377 VINN.n324 VINN.n174 4.5005
R63378 VINN.n253 VINN.n174 4.5005
R63379 VINN.n326 VINN.n174 4.5005
R63380 VINN.n252 VINN.n174 4.5005
R63381 VINN.n328 VINN.n174 4.5005
R63382 VINN.n251 VINN.n174 4.5005
R63383 VINN.n330 VINN.n174 4.5005
R63384 VINN.n250 VINN.n174 4.5005
R63385 VINN.n332 VINN.n174 4.5005
R63386 VINN.n249 VINN.n174 4.5005
R63387 VINN.n334 VINN.n174 4.5005
R63388 VINN.n248 VINN.n174 4.5005
R63389 VINN.n336 VINN.n174 4.5005
R63390 VINN.n247 VINN.n174 4.5005
R63391 VINN.n338 VINN.n174 4.5005
R63392 VINN.n246 VINN.n174 4.5005
R63393 VINN.n340 VINN.n174 4.5005
R63394 VINN.n245 VINN.n174 4.5005
R63395 VINN.n342 VINN.n174 4.5005
R63396 VINN.n244 VINN.n174 4.5005
R63397 VINN.n344 VINN.n174 4.5005
R63398 VINN.n243 VINN.n174 4.5005
R63399 VINN.n346 VINN.n174 4.5005
R63400 VINN.n242 VINN.n174 4.5005
R63401 VINN.n348 VINN.n174 4.5005
R63402 VINN.n241 VINN.n174 4.5005
R63403 VINN.n350 VINN.n174 4.5005
R63404 VINN.n240 VINN.n174 4.5005
R63405 VINN.n352 VINN.n174 4.5005
R63406 VINN.n239 VINN.n174 4.5005
R63407 VINN.n354 VINN.n174 4.5005
R63408 VINN.n238 VINN.n174 4.5005
R63409 VINN.n356 VINN.n174 4.5005
R63410 VINN.n237 VINN.n174 4.5005
R63411 VINN.n358 VINN.n174 4.5005
R63412 VINN.n236 VINN.n174 4.5005
R63413 VINN.n360 VINN.n174 4.5005
R63414 VINN.n235 VINN.n174 4.5005
R63415 VINN.n362 VINN.n174 4.5005
R63416 VINN.n234 VINN.n174 4.5005
R63417 VINN.n364 VINN.n174 4.5005
R63418 VINN.n233 VINN.n174 4.5005
R63419 VINN.n366 VINN.n174 4.5005
R63420 VINN.n232 VINN.n174 4.5005
R63421 VINN.n368 VINN.n174 4.5005
R63422 VINN.n231 VINN.n174 4.5005
R63423 VINN.n370 VINN.n174 4.5005
R63424 VINN.n230 VINN.n174 4.5005
R63425 VINN.n372 VINN.n174 4.5005
R63426 VINN.n229 VINN.n174 4.5005
R63427 VINN.n374 VINN.n174 4.5005
R63428 VINN.n228 VINN.n174 4.5005
R63429 VINN.n376 VINN.n174 4.5005
R63430 VINN.n227 VINN.n174 4.5005
R63431 VINN.n378 VINN.n174 4.5005
R63432 VINN.n226 VINN.n174 4.5005
R63433 VINN.n380 VINN.n174 4.5005
R63434 VINN.n225 VINN.n174 4.5005
R63435 VINN.n382 VINN.n174 4.5005
R63436 VINN.n224 VINN.n174 4.5005
R63437 VINN.n384 VINN.n174 4.5005
R63438 VINN.n223 VINN.n174 4.5005
R63439 VINN.n386 VINN.n174 4.5005
R63440 VINN.n222 VINN.n174 4.5005
R63441 VINN.n388 VINN.n174 4.5005
R63442 VINN.n221 VINN.n174 4.5005
R63443 VINN.n390 VINN.n174 4.5005
R63444 VINN.n220 VINN.n174 4.5005
R63445 VINN.n392 VINN.n174 4.5005
R63446 VINN.n219 VINN.n174 4.5005
R63447 VINN.n394 VINN.n174 4.5005
R63448 VINN.n218 VINN.n174 4.5005
R63449 VINN.n396 VINN.n174 4.5005
R63450 VINN.n217 VINN.n174 4.5005
R63451 VINN.n398 VINN.n174 4.5005
R63452 VINN.n216 VINN.n174 4.5005
R63453 VINN.n400 VINN.n174 4.5005
R63454 VINN.n215 VINN.n174 4.5005
R63455 VINN.n654 VINN.n174 4.5005
R63456 VINN.n656 VINN.n174 4.5005
R63457 VINN.n174 VINN.n0 4.5005
R63458 VINN.n278 VINN.n126 4.5005
R63459 VINN.n276 VINN.n126 4.5005
R63460 VINN.n280 VINN.n126 4.5005
R63461 VINN.n275 VINN.n126 4.5005
R63462 VINN.n282 VINN.n126 4.5005
R63463 VINN.n274 VINN.n126 4.5005
R63464 VINN.n284 VINN.n126 4.5005
R63465 VINN.n273 VINN.n126 4.5005
R63466 VINN.n286 VINN.n126 4.5005
R63467 VINN.n272 VINN.n126 4.5005
R63468 VINN.n288 VINN.n126 4.5005
R63469 VINN.n271 VINN.n126 4.5005
R63470 VINN.n290 VINN.n126 4.5005
R63471 VINN.n270 VINN.n126 4.5005
R63472 VINN.n292 VINN.n126 4.5005
R63473 VINN.n269 VINN.n126 4.5005
R63474 VINN.n294 VINN.n126 4.5005
R63475 VINN.n268 VINN.n126 4.5005
R63476 VINN.n296 VINN.n126 4.5005
R63477 VINN.n267 VINN.n126 4.5005
R63478 VINN.n298 VINN.n126 4.5005
R63479 VINN.n266 VINN.n126 4.5005
R63480 VINN.n300 VINN.n126 4.5005
R63481 VINN.n265 VINN.n126 4.5005
R63482 VINN.n302 VINN.n126 4.5005
R63483 VINN.n264 VINN.n126 4.5005
R63484 VINN.n304 VINN.n126 4.5005
R63485 VINN.n263 VINN.n126 4.5005
R63486 VINN.n306 VINN.n126 4.5005
R63487 VINN.n262 VINN.n126 4.5005
R63488 VINN.n308 VINN.n126 4.5005
R63489 VINN.n261 VINN.n126 4.5005
R63490 VINN.n310 VINN.n126 4.5005
R63491 VINN.n260 VINN.n126 4.5005
R63492 VINN.n312 VINN.n126 4.5005
R63493 VINN.n259 VINN.n126 4.5005
R63494 VINN.n314 VINN.n126 4.5005
R63495 VINN.n258 VINN.n126 4.5005
R63496 VINN.n316 VINN.n126 4.5005
R63497 VINN.n257 VINN.n126 4.5005
R63498 VINN.n318 VINN.n126 4.5005
R63499 VINN.n256 VINN.n126 4.5005
R63500 VINN.n320 VINN.n126 4.5005
R63501 VINN.n255 VINN.n126 4.5005
R63502 VINN.n322 VINN.n126 4.5005
R63503 VINN.n254 VINN.n126 4.5005
R63504 VINN.n324 VINN.n126 4.5005
R63505 VINN.n253 VINN.n126 4.5005
R63506 VINN.n326 VINN.n126 4.5005
R63507 VINN.n252 VINN.n126 4.5005
R63508 VINN.n328 VINN.n126 4.5005
R63509 VINN.n251 VINN.n126 4.5005
R63510 VINN.n330 VINN.n126 4.5005
R63511 VINN.n250 VINN.n126 4.5005
R63512 VINN.n332 VINN.n126 4.5005
R63513 VINN.n249 VINN.n126 4.5005
R63514 VINN.n334 VINN.n126 4.5005
R63515 VINN.n248 VINN.n126 4.5005
R63516 VINN.n336 VINN.n126 4.5005
R63517 VINN.n247 VINN.n126 4.5005
R63518 VINN.n338 VINN.n126 4.5005
R63519 VINN.n246 VINN.n126 4.5005
R63520 VINN.n340 VINN.n126 4.5005
R63521 VINN.n245 VINN.n126 4.5005
R63522 VINN.n342 VINN.n126 4.5005
R63523 VINN.n244 VINN.n126 4.5005
R63524 VINN.n344 VINN.n126 4.5005
R63525 VINN.n243 VINN.n126 4.5005
R63526 VINN.n346 VINN.n126 4.5005
R63527 VINN.n242 VINN.n126 4.5005
R63528 VINN.n348 VINN.n126 4.5005
R63529 VINN.n241 VINN.n126 4.5005
R63530 VINN.n350 VINN.n126 4.5005
R63531 VINN.n240 VINN.n126 4.5005
R63532 VINN.n352 VINN.n126 4.5005
R63533 VINN.n239 VINN.n126 4.5005
R63534 VINN.n354 VINN.n126 4.5005
R63535 VINN.n238 VINN.n126 4.5005
R63536 VINN.n356 VINN.n126 4.5005
R63537 VINN.n237 VINN.n126 4.5005
R63538 VINN.n358 VINN.n126 4.5005
R63539 VINN.n236 VINN.n126 4.5005
R63540 VINN.n360 VINN.n126 4.5005
R63541 VINN.n235 VINN.n126 4.5005
R63542 VINN.n362 VINN.n126 4.5005
R63543 VINN.n234 VINN.n126 4.5005
R63544 VINN.n364 VINN.n126 4.5005
R63545 VINN.n233 VINN.n126 4.5005
R63546 VINN.n366 VINN.n126 4.5005
R63547 VINN.n232 VINN.n126 4.5005
R63548 VINN.n368 VINN.n126 4.5005
R63549 VINN.n231 VINN.n126 4.5005
R63550 VINN.n370 VINN.n126 4.5005
R63551 VINN.n230 VINN.n126 4.5005
R63552 VINN.n372 VINN.n126 4.5005
R63553 VINN.n229 VINN.n126 4.5005
R63554 VINN.n374 VINN.n126 4.5005
R63555 VINN.n228 VINN.n126 4.5005
R63556 VINN.n376 VINN.n126 4.5005
R63557 VINN.n227 VINN.n126 4.5005
R63558 VINN.n378 VINN.n126 4.5005
R63559 VINN.n226 VINN.n126 4.5005
R63560 VINN.n380 VINN.n126 4.5005
R63561 VINN.n225 VINN.n126 4.5005
R63562 VINN.n382 VINN.n126 4.5005
R63563 VINN.n224 VINN.n126 4.5005
R63564 VINN.n384 VINN.n126 4.5005
R63565 VINN.n223 VINN.n126 4.5005
R63566 VINN.n386 VINN.n126 4.5005
R63567 VINN.n222 VINN.n126 4.5005
R63568 VINN.n388 VINN.n126 4.5005
R63569 VINN.n221 VINN.n126 4.5005
R63570 VINN.n390 VINN.n126 4.5005
R63571 VINN.n220 VINN.n126 4.5005
R63572 VINN.n392 VINN.n126 4.5005
R63573 VINN.n219 VINN.n126 4.5005
R63574 VINN.n394 VINN.n126 4.5005
R63575 VINN.n218 VINN.n126 4.5005
R63576 VINN.n396 VINN.n126 4.5005
R63577 VINN.n217 VINN.n126 4.5005
R63578 VINN.n398 VINN.n126 4.5005
R63579 VINN.n216 VINN.n126 4.5005
R63580 VINN.n400 VINN.n126 4.5005
R63581 VINN.n215 VINN.n126 4.5005
R63582 VINN.n654 VINN.n126 4.5005
R63583 VINN.n656 VINN.n126 4.5005
R63584 VINN.n126 VINN.n0 4.5005
R63585 VINN.n278 VINN.n175 4.5005
R63586 VINN.n276 VINN.n175 4.5005
R63587 VINN.n280 VINN.n175 4.5005
R63588 VINN.n275 VINN.n175 4.5005
R63589 VINN.n282 VINN.n175 4.5005
R63590 VINN.n274 VINN.n175 4.5005
R63591 VINN.n284 VINN.n175 4.5005
R63592 VINN.n273 VINN.n175 4.5005
R63593 VINN.n286 VINN.n175 4.5005
R63594 VINN.n272 VINN.n175 4.5005
R63595 VINN.n288 VINN.n175 4.5005
R63596 VINN.n271 VINN.n175 4.5005
R63597 VINN.n290 VINN.n175 4.5005
R63598 VINN.n270 VINN.n175 4.5005
R63599 VINN.n292 VINN.n175 4.5005
R63600 VINN.n269 VINN.n175 4.5005
R63601 VINN.n294 VINN.n175 4.5005
R63602 VINN.n268 VINN.n175 4.5005
R63603 VINN.n296 VINN.n175 4.5005
R63604 VINN.n267 VINN.n175 4.5005
R63605 VINN.n298 VINN.n175 4.5005
R63606 VINN.n266 VINN.n175 4.5005
R63607 VINN.n300 VINN.n175 4.5005
R63608 VINN.n265 VINN.n175 4.5005
R63609 VINN.n302 VINN.n175 4.5005
R63610 VINN.n264 VINN.n175 4.5005
R63611 VINN.n304 VINN.n175 4.5005
R63612 VINN.n263 VINN.n175 4.5005
R63613 VINN.n306 VINN.n175 4.5005
R63614 VINN.n262 VINN.n175 4.5005
R63615 VINN.n308 VINN.n175 4.5005
R63616 VINN.n261 VINN.n175 4.5005
R63617 VINN.n310 VINN.n175 4.5005
R63618 VINN.n260 VINN.n175 4.5005
R63619 VINN.n312 VINN.n175 4.5005
R63620 VINN.n259 VINN.n175 4.5005
R63621 VINN.n314 VINN.n175 4.5005
R63622 VINN.n258 VINN.n175 4.5005
R63623 VINN.n316 VINN.n175 4.5005
R63624 VINN.n257 VINN.n175 4.5005
R63625 VINN.n318 VINN.n175 4.5005
R63626 VINN.n256 VINN.n175 4.5005
R63627 VINN.n320 VINN.n175 4.5005
R63628 VINN.n255 VINN.n175 4.5005
R63629 VINN.n322 VINN.n175 4.5005
R63630 VINN.n254 VINN.n175 4.5005
R63631 VINN.n324 VINN.n175 4.5005
R63632 VINN.n253 VINN.n175 4.5005
R63633 VINN.n326 VINN.n175 4.5005
R63634 VINN.n252 VINN.n175 4.5005
R63635 VINN.n328 VINN.n175 4.5005
R63636 VINN.n251 VINN.n175 4.5005
R63637 VINN.n330 VINN.n175 4.5005
R63638 VINN.n250 VINN.n175 4.5005
R63639 VINN.n332 VINN.n175 4.5005
R63640 VINN.n249 VINN.n175 4.5005
R63641 VINN.n334 VINN.n175 4.5005
R63642 VINN.n248 VINN.n175 4.5005
R63643 VINN.n336 VINN.n175 4.5005
R63644 VINN.n247 VINN.n175 4.5005
R63645 VINN.n338 VINN.n175 4.5005
R63646 VINN.n246 VINN.n175 4.5005
R63647 VINN.n340 VINN.n175 4.5005
R63648 VINN.n245 VINN.n175 4.5005
R63649 VINN.n342 VINN.n175 4.5005
R63650 VINN.n244 VINN.n175 4.5005
R63651 VINN.n344 VINN.n175 4.5005
R63652 VINN.n243 VINN.n175 4.5005
R63653 VINN.n346 VINN.n175 4.5005
R63654 VINN.n242 VINN.n175 4.5005
R63655 VINN.n348 VINN.n175 4.5005
R63656 VINN.n241 VINN.n175 4.5005
R63657 VINN.n350 VINN.n175 4.5005
R63658 VINN.n240 VINN.n175 4.5005
R63659 VINN.n352 VINN.n175 4.5005
R63660 VINN.n239 VINN.n175 4.5005
R63661 VINN.n354 VINN.n175 4.5005
R63662 VINN.n238 VINN.n175 4.5005
R63663 VINN.n356 VINN.n175 4.5005
R63664 VINN.n237 VINN.n175 4.5005
R63665 VINN.n358 VINN.n175 4.5005
R63666 VINN.n236 VINN.n175 4.5005
R63667 VINN.n360 VINN.n175 4.5005
R63668 VINN.n235 VINN.n175 4.5005
R63669 VINN.n362 VINN.n175 4.5005
R63670 VINN.n234 VINN.n175 4.5005
R63671 VINN.n364 VINN.n175 4.5005
R63672 VINN.n233 VINN.n175 4.5005
R63673 VINN.n366 VINN.n175 4.5005
R63674 VINN.n232 VINN.n175 4.5005
R63675 VINN.n368 VINN.n175 4.5005
R63676 VINN.n231 VINN.n175 4.5005
R63677 VINN.n370 VINN.n175 4.5005
R63678 VINN.n230 VINN.n175 4.5005
R63679 VINN.n372 VINN.n175 4.5005
R63680 VINN.n229 VINN.n175 4.5005
R63681 VINN.n374 VINN.n175 4.5005
R63682 VINN.n228 VINN.n175 4.5005
R63683 VINN.n376 VINN.n175 4.5005
R63684 VINN.n227 VINN.n175 4.5005
R63685 VINN.n378 VINN.n175 4.5005
R63686 VINN.n226 VINN.n175 4.5005
R63687 VINN.n380 VINN.n175 4.5005
R63688 VINN.n225 VINN.n175 4.5005
R63689 VINN.n382 VINN.n175 4.5005
R63690 VINN.n224 VINN.n175 4.5005
R63691 VINN.n384 VINN.n175 4.5005
R63692 VINN.n223 VINN.n175 4.5005
R63693 VINN.n386 VINN.n175 4.5005
R63694 VINN.n222 VINN.n175 4.5005
R63695 VINN.n388 VINN.n175 4.5005
R63696 VINN.n221 VINN.n175 4.5005
R63697 VINN.n390 VINN.n175 4.5005
R63698 VINN.n220 VINN.n175 4.5005
R63699 VINN.n392 VINN.n175 4.5005
R63700 VINN.n219 VINN.n175 4.5005
R63701 VINN.n394 VINN.n175 4.5005
R63702 VINN.n218 VINN.n175 4.5005
R63703 VINN.n396 VINN.n175 4.5005
R63704 VINN.n217 VINN.n175 4.5005
R63705 VINN.n398 VINN.n175 4.5005
R63706 VINN.n216 VINN.n175 4.5005
R63707 VINN.n400 VINN.n175 4.5005
R63708 VINN.n215 VINN.n175 4.5005
R63709 VINN.n654 VINN.n175 4.5005
R63710 VINN.n656 VINN.n175 4.5005
R63711 VINN.n175 VINN.n0 4.5005
R63712 VINN.n278 VINN.n125 4.5005
R63713 VINN.n276 VINN.n125 4.5005
R63714 VINN.n280 VINN.n125 4.5005
R63715 VINN.n275 VINN.n125 4.5005
R63716 VINN.n282 VINN.n125 4.5005
R63717 VINN.n274 VINN.n125 4.5005
R63718 VINN.n284 VINN.n125 4.5005
R63719 VINN.n273 VINN.n125 4.5005
R63720 VINN.n286 VINN.n125 4.5005
R63721 VINN.n272 VINN.n125 4.5005
R63722 VINN.n288 VINN.n125 4.5005
R63723 VINN.n271 VINN.n125 4.5005
R63724 VINN.n290 VINN.n125 4.5005
R63725 VINN.n270 VINN.n125 4.5005
R63726 VINN.n292 VINN.n125 4.5005
R63727 VINN.n269 VINN.n125 4.5005
R63728 VINN.n294 VINN.n125 4.5005
R63729 VINN.n268 VINN.n125 4.5005
R63730 VINN.n296 VINN.n125 4.5005
R63731 VINN.n267 VINN.n125 4.5005
R63732 VINN.n298 VINN.n125 4.5005
R63733 VINN.n266 VINN.n125 4.5005
R63734 VINN.n300 VINN.n125 4.5005
R63735 VINN.n265 VINN.n125 4.5005
R63736 VINN.n302 VINN.n125 4.5005
R63737 VINN.n264 VINN.n125 4.5005
R63738 VINN.n304 VINN.n125 4.5005
R63739 VINN.n263 VINN.n125 4.5005
R63740 VINN.n306 VINN.n125 4.5005
R63741 VINN.n262 VINN.n125 4.5005
R63742 VINN.n308 VINN.n125 4.5005
R63743 VINN.n261 VINN.n125 4.5005
R63744 VINN.n310 VINN.n125 4.5005
R63745 VINN.n260 VINN.n125 4.5005
R63746 VINN.n312 VINN.n125 4.5005
R63747 VINN.n259 VINN.n125 4.5005
R63748 VINN.n314 VINN.n125 4.5005
R63749 VINN.n258 VINN.n125 4.5005
R63750 VINN.n316 VINN.n125 4.5005
R63751 VINN.n257 VINN.n125 4.5005
R63752 VINN.n318 VINN.n125 4.5005
R63753 VINN.n256 VINN.n125 4.5005
R63754 VINN.n320 VINN.n125 4.5005
R63755 VINN.n255 VINN.n125 4.5005
R63756 VINN.n322 VINN.n125 4.5005
R63757 VINN.n254 VINN.n125 4.5005
R63758 VINN.n324 VINN.n125 4.5005
R63759 VINN.n253 VINN.n125 4.5005
R63760 VINN.n326 VINN.n125 4.5005
R63761 VINN.n252 VINN.n125 4.5005
R63762 VINN.n328 VINN.n125 4.5005
R63763 VINN.n251 VINN.n125 4.5005
R63764 VINN.n330 VINN.n125 4.5005
R63765 VINN.n250 VINN.n125 4.5005
R63766 VINN.n332 VINN.n125 4.5005
R63767 VINN.n249 VINN.n125 4.5005
R63768 VINN.n334 VINN.n125 4.5005
R63769 VINN.n248 VINN.n125 4.5005
R63770 VINN.n336 VINN.n125 4.5005
R63771 VINN.n247 VINN.n125 4.5005
R63772 VINN.n338 VINN.n125 4.5005
R63773 VINN.n246 VINN.n125 4.5005
R63774 VINN.n340 VINN.n125 4.5005
R63775 VINN.n245 VINN.n125 4.5005
R63776 VINN.n342 VINN.n125 4.5005
R63777 VINN.n244 VINN.n125 4.5005
R63778 VINN.n344 VINN.n125 4.5005
R63779 VINN.n243 VINN.n125 4.5005
R63780 VINN.n346 VINN.n125 4.5005
R63781 VINN.n242 VINN.n125 4.5005
R63782 VINN.n348 VINN.n125 4.5005
R63783 VINN.n241 VINN.n125 4.5005
R63784 VINN.n350 VINN.n125 4.5005
R63785 VINN.n240 VINN.n125 4.5005
R63786 VINN.n352 VINN.n125 4.5005
R63787 VINN.n239 VINN.n125 4.5005
R63788 VINN.n354 VINN.n125 4.5005
R63789 VINN.n238 VINN.n125 4.5005
R63790 VINN.n356 VINN.n125 4.5005
R63791 VINN.n237 VINN.n125 4.5005
R63792 VINN.n358 VINN.n125 4.5005
R63793 VINN.n236 VINN.n125 4.5005
R63794 VINN.n360 VINN.n125 4.5005
R63795 VINN.n235 VINN.n125 4.5005
R63796 VINN.n362 VINN.n125 4.5005
R63797 VINN.n234 VINN.n125 4.5005
R63798 VINN.n364 VINN.n125 4.5005
R63799 VINN.n233 VINN.n125 4.5005
R63800 VINN.n366 VINN.n125 4.5005
R63801 VINN.n232 VINN.n125 4.5005
R63802 VINN.n368 VINN.n125 4.5005
R63803 VINN.n231 VINN.n125 4.5005
R63804 VINN.n370 VINN.n125 4.5005
R63805 VINN.n230 VINN.n125 4.5005
R63806 VINN.n372 VINN.n125 4.5005
R63807 VINN.n229 VINN.n125 4.5005
R63808 VINN.n374 VINN.n125 4.5005
R63809 VINN.n228 VINN.n125 4.5005
R63810 VINN.n376 VINN.n125 4.5005
R63811 VINN.n227 VINN.n125 4.5005
R63812 VINN.n378 VINN.n125 4.5005
R63813 VINN.n226 VINN.n125 4.5005
R63814 VINN.n380 VINN.n125 4.5005
R63815 VINN.n225 VINN.n125 4.5005
R63816 VINN.n382 VINN.n125 4.5005
R63817 VINN.n224 VINN.n125 4.5005
R63818 VINN.n384 VINN.n125 4.5005
R63819 VINN.n223 VINN.n125 4.5005
R63820 VINN.n386 VINN.n125 4.5005
R63821 VINN.n222 VINN.n125 4.5005
R63822 VINN.n388 VINN.n125 4.5005
R63823 VINN.n221 VINN.n125 4.5005
R63824 VINN.n390 VINN.n125 4.5005
R63825 VINN.n220 VINN.n125 4.5005
R63826 VINN.n392 VINN.n125 4.5005
R63827 VINN.n219 VINN.n125 4.5005
R63828 VINN.n394 VINN.n125 4.5005
R63829 VINN.n218 VINN.n125 4.5005
R63830 VINN.n396 VINN.n125 4.5005
R63831 VINN.n217 VINN.n125 4.5005
R63832 VINN.n398 VINN.n125 4.5005
R63833 VINN.n216 VINN.n125 4.5005
R63834 VINN.n400 VINN.n125 4.5005
R63835 VINN.n215 VINN.n125 4.5005
R63836 VINN.n654 VINN.n125 4.5005
R63837 VINN.n656 VINN.n125 4.5005
R63838 VINN.n125 VINN.n0 4.5005
R63839 VINN.n278 VINN.n176 4.5005
R63840 VINN.n276 VINN.n176 4.5005
R63841 VINN.n280 VINN.n176 4.5005
R63842 VINN.n275 VINN.n176 4.5005
R63843 VINN.n282 VINN.n176 4.5005
R63844 VINN.n274 VINN.n176 4.5005
R63845 VINN.n284 VINN.n176 4.5005
R63846 VINN.n273 VINN.n176 4.5005
R63847 VINN.n286 VINN.n176 4.5005
R63848 VINN.n272 VINN.n176 4.5005
R63849 VINN.n288 VINN.n176 4.5005
R63850 VINN.n271 VINN.n176 4.5005
R63851 VINN.n290 VINN.n176 4.5005
R63852 VINN.n270 VINN.n176 4.5005
R63853 VINN.n292 VINN.n176 4.5005
R63854 VINN.n269 VINN.n176 4.5005
R63855 VINN.n294 VINN.n176 4.5005
R63856 VINN.n268 VINN.n176 4.5005
R63857 VINN.n296 VINN.n176 4.5005
R63858 VINN.n267 VINN.n176 4.5005
R63859 VINN.n298 VINN.n176 4.5005
R63860 VINN.n266 VINN.n176 4.5005
R63861 VINN.n300 VINN.n176 4.5005
R63862 VINN.n265 VINN.n176 4.5005
R63863 VINN.n302 VINN.n176 4.5005
R63864 VINN.n264 VINN.n176 4.5005
R63865 VINN.n304 VINN.n176 4.5005
R63866 VINN.n263 VINN.n176 4.5005
R63867 VINN.n306 VINN.n176 4.5005
R63868 VINN.n262 VINN.n176 4.5005
R63869 VINN.n308 VINN.n176 4.5005
R63870 VINN.n261 VINN.n176 4.5005
R63871 VINN.n310 VINN.n176 4.5005
R63872 VINN.n260 VINN.n176 4.5005
R63873 VINN.n312 VINN.n176 4.5005
R63874 VINN.n259 VINN.n176 4.5005
R63875 VINN.n314 VINN.n176 4.5005
R63876 VINN.n258 VINN.n176 4.5005
R63877 VINN.n316 VINN.n176 4.5005
R63878 VINN.n257 VINN.n176 4.5005
R63879 VINN.n318 VINN.n176 4.5005
R63880 VINN.n256 VINN.n176 4.5005
R63881 VINN.n320 VINN.n176 4.5005
R63882 VINN.n255 VINN.n176 4.5005
R63883 VINN.n322 VINN.n176 4.5005
R63884 VINN.n254 VINN.n176 4.5005
R63885 VINN.n324 VINN.n176 4.5005
R63886 VINN.n253 VINN.n176 4.5005
R63887 VINN.n326 VINN.n176 4.5005
R63888 VINN.n252 VINN.n176 4.5005
R63889 VINN.n328 VINN.n176 4.5005
R63890 VINN.n251 VINN.n176 4.5005
R63891 VINN.n330 VINN.n176 4.5005
R63892 VINN.n250 VINN.n176 4.5005
R63893 VINN.n332 VINN.n176 4.5005
R63894 VINN.n249 VINN.n176 4.5005
R63895 VINN.n334 VINN.n176 4.5005
R63896 VINN.n248 VINN.n176 4.5005
R63897 VINN.n336 VINN.n176 4.5005
R63898 VINN.n247 VINN.n176 4.5005
R63899 VINN.n338 VINN.n176 4.5005
R63900 VINN.n246 VINN.n176 4.5005
R63901 VINN.n340 VINN.n176 4.5005
R63902 VINN.n245 VINN.n176 4.5005
R63903 VINN.n342 VINN.n176 4.5005
R63904 VINN.n244 VINN.n176 4.5005
R63905 VINN.n344 VINN.n176 4.5005
R63906 VINN.n243 VINN.n176 4.5005
R63907 VINN.n346 VINN.n176 4.5005
R63908 VINN.n242 VINN.n176 4.5005
R63909 VINN.n348 VINN.n176 4.5005
R63910 VINN.n241 VINN.n176 4.5005
R63911 VINN.n350 VINN.n176 4.5005
R63912 VINN.n240 VINN.n176 4.5005
R63913 VINN.n352 VINN.n176 4.5005
R63914 VINN.n239 VINN.n176 4.5005
R63915 VINN.n354 VINN.n176 4.5005
R63916 VINN.n238 VINN.n176 4.5005
R63917 VINN.n356 VINN.n176 4.5005
R63918 VINN.n237 VINN.n176 4.5005
R63919 VINN.n358 VINN.n176 4.5005
R63920 VINN.n236 VINN.n176 4.5005
R63921 VINN.n360 VINN.n176 4.5005
R63922 VINN.n235 VINN.n176 4.5005
R63923 VINN.n362 VINN.n176 4.5005
R63924 VINN.n234 VINN.n176 4.5005
R63925 VINN.n364 VINN.n176 4.5005
R63926 VINN.n233 VINN.n176 4.5005
R63927 VINN.n366 VINN.n176 4.5005
R63928 VINN.n232 VINN.n176 4.5005
R63929 VINN.n368 VINN.n176 4.5005
R63930 VINN.n231 VINN.n176 4.5005
R63931 VINN.n370 VINN.n176 4.5005
R63932 VINN.n230 VINN.n176 4.5005
R63933 VINN.n372 VINN.n176 4.5005
R63934 VINN.n229 VINN.n176 4.5005
R63935 VINN.n374 VINN.n176 4.5005
R63936 VINN.n228 VINN.n176 4.5005
R63937 VINN.n376 VINN.n176 4.5005
R63938 VINN.n227 VINN.n176 4.5005
R63939 VINN.n378 VINN.n176 4.5005
R63940 VINN.n226 VINN.n176 4.5005
R63941 VINN.n380 VINN.n176 4.5005
R63942 VINN.n225 VINN.n176 4.5005
R63943 VINN.n382 VINN.n176 4.5005
R63944 VINN.n224 VINN.n176 4.5005
R63945 VINN.n384 VINN.n176 4.5005
R63946 VINN.n223 VINN.n176 4.5005
R63947 VINN.n386 VINN.n176 4.5005
R63948 VINN.n222 VINN.n176 4.5005
R63949 VINN.n388 VINN.n176 4.5005
R63950 VINN.n221 VINN.n176 4.5005
R63951 VINN.n390 VINN.n176 4.5005
R63952 VINN.n220 VINN.n176 4.5005
R63953 VINN.n392 VINN.n176 4.5005
R63954 VINN.n219 VINN.n176 4.5005
R63955 VINN.n394 VINN.n176 4.5005
R63956 VINN.n218 VINN.n176 4.5005
R63957 VINN.n396 VINN.n176 4.5005
R63958 VINN.n217 VINN.n176 4.5005
R63959 VINN.n398 VINN.n176 4.5005
R63960 VINN.n216 VINN.n176 4.5005
R63961 VINN.n400 VINN.n176 4.5005
R63962 VINN.n215 VINN.n176 4.5005
R63963 VINN.n654 VINN.n176 4.5005
R63964 VINN.n656 VINN.n176 4.5005
R63965 VINN.n176 VINN.n0 4.5005
R63966 VINN.n278 VINN.n124 4.5005
R63967 VINN.n276 VINN.n124 4.5005
R63968 VINN.n280 VINN.n124 4.5005
R63969 VINN.n275 VINN.n124 4.5005
R63970 VINN.n282 VINN.n124 4.5005
R63971 VINN.n274 VINN.n124 4.5005
R63972 VINN.n284 VINN.n124 4.5005
R63973 VINN.n273 VINN.n124 4.5005
R63974 VINN.n286 VINN.n124 4.5005
R63975 VINN.n272 VINN.n124 4.5005
R63976 VINN.n288 VINN.n124 4.5005
R63977 VINN.n271 VINN.n124 4.5005
R63978 VINN.n290 VINN.n124 4.5005
R63979 VINN.n270 VINN.n124 4.5005
R63980 VINN.n292 VINN.n124 4.5005
R63981 VINN.n269 VINN.n124 4.5005
R63982 VINN.n294 VINN.n124 4.5005
R63983 VINN.n268 VINN.n124 4.5005
R63984 VINN.n296 VINN.n124 4.5005
R63985 VINN.n267 VINN.n124 4.5005
R63986 VINN.n298 VINN.n124 4.5005
R63987 VINN.n266 VINN.n124 4.5005
R63988 VINN.n300 VINN.n124 4.5005
R63989 VINN.n265 VINN.n124 4.5005
R63990 VINN.n302 VINN.n124 4.5005
R63991 VINN.n264 VINN.n124 4.5005
R63992 VINN.n304 VINN.n124 4.5005
R63993 VINN.n263 VINN.n124 4.5005
R63994 VINN.n306 VINN.n124 4.5005
R63995 VINN.n262 VINN.n124 4.5005
R63996 VINN.n308 VINN.n124 4.5005
R63997 VINN.n261 VINN.n124 4.5005
R63998 VINN.n310 VINN.n124 4.5005
R63999 VINN.n260 VINN.n124 4.5005
R64000 VINN.n312 VINN.n124 4.5005
R64001 VINN.n259 VINN.n124 4.5005
R64002 VINN.n314 VINN.n124 4.5005
R64003 VINN.n258 VINN.n124 4.5005
R64004 VINN.n316 VINN.n124 4.5005
R64005 VINN.n257 VINN.n124 4.5005
R64006 VINN.n318 VINN.n124 4.5005
R64007 VINN.n256 VINN.n124 4.5005
R64008 VINN.n320 VINN.n124 4.5005
R64009 VINN.n255 VINN.n124 4.5005
R64010 VINN.n322 VINN.n124 4.5005
R64011 VINN.n254 VINN.n124 4.5005
R64012 VINN.n324 VINN.n124 4.5005
R64013 VINN.n253 VINN.n124 4.5005
R64014 VINN.n326 VINN.n124 4.5005
R64015 VINN.n252 VINN.n124 4.5005
R64016 VINN.n328 VINN.n124 4.5005
R64017 VINN.n251 VINN.n124 4.5005
R64018 VINN.n330 VINN.n124 4.5005
R64019 VINN.n250 VINN.n124 4.5005
R64020 VINN.n332 VINN.n124 4.5005
R64021 VINN.n249 VINN.n124 4.5005
R64022 VINN.n334 VINN.n124 4.5005
R64023 VINN.n248 VINN.n124 4.5005
R64024 VINN.n336 VINN.n124 4.5005
R64025 VINN.n247 VINN.n124 4.5005
R64026 VINN.n338 VINN.n124 4.5005
R64027 VINN.n246 VINN.n124 4.5005
R64028 VINN.n340 VINN.n124 4.5005
R64029 VINN.n245 VINN.n124 4.5005
R64030 VINN.n342 VINN.n124 4.5005
R64031 VINN.n244 VINN.n124 4.5005
R64032 VINN.n344 VINN.n124 4.5005
R64033 VINN.n243 VINN.n124 4.5005
R64034 VINN.n346 VINN.n124 4.5005
R64035 VINN.n242 VINN.n124 4.5005
R64036 VINN.n348 VINN.n124 4.5005
R64037 VINN.n241 VINN.n124 4.5005
R64038 VINN.n350 VINN.n124 4.5005
R64039 VINN.n240 VINN.n124 4.5005
R64040 VINN.n352 VINN.n124 4.5005
R64041 VINN.n239 VINN.n124 4.5005
R64042 VINN.n354 VINN.n124 4.5005
R64043 VINN.n238 VINN.n124 4.5005
R64044 VINN.n356 VINN.n124 4.5005
R64045 VINN.n237 VINN.n124 4.5005
R64046 VINN.n358 VINN.n124 4.5005
R64047 VINN.n236 VINN.n124 4.5005
R64048 VINN.n360 VINN.n124 4.5005
R64049 VINN.n235 VINN.n124 4.5005
R64050 VINN.n362 VINN.n124 4.5005
R64051 VINN.n234 VINN.n124 4.5005
R64052 VINN.n364 VINN.n124 4.5005
R64053 VINN.n233 VINN.n124 4.5005
R64054 VINN.n366 VINN.n124 4.5005
R64055 VINN.n232 VINN.n124 4.5005
R64056 VINN.n368 VINN.n124 4.5005
R64057 VINN.n231 VINN.n124 4.5005
R64058 VINN.n370 VINN.n124 4.5005
R64059 VINN.n230 VINN.n124 4.5005
R64060 VINN.n372 VINN.n124 4.5005
R64061 VINN.n229 VINN.n124 4.5005
R64062 VINN.n374 VINN.n124 4.5005
R64063 VINN.n228 VINN.n124 4.5005
R64064 VINN.n376 VINN.n124 4.5005
R64065 VINN.n227 VINN.n124 4.5005
R64066 VINN.n378 VINN.n124 4.5005
R64067 VINN.n226 VINN.n124 4.5005
R64068 VINN.n380 VINN.n124 4.5005
R64069 VINN.n225 VINN.n124 4.5005
R64070 VINN.n382 VINN.n124 4.5005
R64071 VINN.n224 VINN.n124 4.5005
R64072 VINN.n384 VINN.n124 4.5005
R64073 VINN.n223 VINN.n124 4.5005
R64074 VINN.n386 VINN.n124 4.5005
R64075 VINN.n222 VINN.n124 4.5005
R64076 VINN.n388 VINN.n124 4.5005
R64077 VINN.n221 VINN.n124 4.5005
R64078 VINN.n390 VINN.n124 4.5005
R64079 VINN.n220 VINN.n124 4.5005
R64080 VINN.n392 VINN.n124 4.5005
R64081 VINN.n219 VINN.n124 4.5005
R64082 VINN.n394 VINN.n124 4.5005
R64083 VINN.n218 VINN.n124 4.5005
R64084 VINN.n396 VINN.n124 4.5005
R64085 VINN.n217 VINN.n124 4.5005
R64086 VINN.n398 VINN.n124 4.5005
R64087 VINN.n216 VINN.n124 4.5005
R64088 VINN.n400 VINN.n124 4.5005
R64089 VINN.n215 VINN.n124 4.5005
R64090 VINN.n654 VINN.n124 4.5005
R64091 VINN.n656 VINN.n124 4.5005
R64092 VINN.n124 VINN.n0 4.5005
R64093 VINN.n278 VINN.n177 4.5005
R64094 VINN.n276 VINN.n177 4.5005
R64095 VINN.n280 VINN.n177 4.5005
R64096 VINN.n275 VINN.n177 4.5005
R64097 VINN.n282 VINN.n177 4.5005
R64098 VINN.n274 VINN.n177 4.5005
R64099 VINN.n284 VINN.n177 4.5005
R64100 VINN.n273 VINN.n177 4.5005
R64101 VINN.n286 VINN.n177 4.5005
R64102 VINN.n272 VINN.n177 4.5005
R64103 VINN.n288 VINN.n177 4.5005
R64104 VINN.n271 VINN.n177 4.5005
R64105 VINN.n290 VINN.n177 4.5005
R64106 VINN.n270 VINN.n177 4.5005
R64107 VINN.n292 VINN.n177 4.5005
R64108 VINN.n269 VINN.n177 4.5005
R64109 VINN.n294 VINN.n177 4.5005
R64110 VINN.n268 VINN.n177 4.5005
R64111 VINN.n296 VINN.n177 4.5005
R64112 VINN.n267 VINN.n177 4.5005
R64113 VINN.n298 VINN.n177 4.5005
R64114 VINN.n266 VINN.n177 4.5005
R64115 VINN.n300 VINN.n177 4.5005
R64116 VINN.n265 VINN.n177 4.5005
R64117 VINN.n302 VINN.n177 4.5005
R64118 VINN.n264 VINN.n177 4.5005
R64119 VINN.n304 VINN.n177 4.5005
R64120 VINN.n263 VINN.n177 4.5005
R64121 VINN.n306 VINN.n177 4.5005
R64122 VINN.n262 VINN.n177 4.5005
R64123 VINN.n308 VINN.n177 4.5005
R64124 VINN.n261 VINN.n177 4.5005
R64125 VINN.n310 VINN.n177 4.5005
R64126 VINN.n260 VINN.n177 4.5005
R64127 VINN.n312 VINN.n177 4.5005
R64128 VINN.n259 VINN.n177 4.5005
R64129 VINN.n314 VINN.n177 4.5005
R64130 VINN.n258 VINN.n177 4.5005
R64131 VINN.n316 VINN.n177 4.5005
R64132 VINN.n257 VINN.n177 4.5005
R64133 VINN.n318 VINN.n177 4.5005
R64134 VINN.n256 VINN.n177 4.5005
R64135 VINN.n320 VINN.n177 4.5005
R64136 VINN.n255 VINN.n177 4.5005
R64137 VINN.n322 VINN.n177 4.5005
R64138 VINN.n254 VINN.n177 4.5005
R64139 VINN.n324 VINN.n177 4.5005
R64140 VINN.n253 VINN.n177 4.5005
R64141 VINN.n326 VINN.n177 4.5005
R64142 VINN.n252 VINN.n177 4.5005
R64143 VINN.n328 VINN.n177 4.5005
R64144 VINN.n251 VINN.n177 4.5005
R64145 VINN.n330 VINN.n177 4.5005
R64146 VINN.n250 VINN.n177 4.5005
R64147 VINN.n332 VINN.n177 4.5005
R64148 VINN.n249 VINN.n177 4.5005
R64149 VINN.n334 VINN.n177 4.5005
R64150 VINN.n248 VINN.n177 4.5005
R64151 VINN.n336 VINN.n177 4.5005
R64152 VINN.n247 VINN.n177 4.5005
R64153 VINN.n338 VINN.n177 4.5005
R64154 VINN.n246 VINN.n177 4.5005
R64155 VINN.n340 VINN.n177 4.5005
R64156 VINN.n245 VINN.n177 4.5005
R64157 VINN.n342 VINN.n177 4.5005
R64158 VINN.n244 VINN.n177 4.5005
R64159 VINN.n344 VINN.n177 4.5005
R64160 VINN.n243 VINN.n177 4.5005
R64161 VINN.n346 VINN.n177 4.5005
R64162 VINN.n242 VINN.n177 4.5005
R64163 VINN.n348 VINN.n177 4.5005
R64164 VINN.n241 VINN.n177 4.5005
R64165 VINN.n350 VINN.n177 4.5005
R64166 VINN.n240 VINN.n177 4.5005
R64167 VINN.n352 VINN.n177 4.5005
R64168 VINN.n239 VINN.n177 4.5005
R64169 VINN.n354 VINN.n177 4.5005
R64170 VINN.n238 VINN.n177 4.5005
R64171 VINN.n356 VINN.n177 4.5005
R64172 VINN.n237 VINN.n177 4.5005
R64173 VINN.n358 VINN.n177 4.5005
R64174 VINN.n236 VINN.n177 4.5005
R64175 VINN.n360 VINN.n177 4.5005
R64176 VINN.n235 VINN.n177 4.5005
R64177 VINN.n362 VINN.n177 4.5005
R64178 VINN.n234 VINN.n177 4.5005
R64179 VINN.n364 VINN.n177 4.5005
R64180 VINN.n233 VINN.n177 4.5005
R64181 VINN.n366 VINN.n177 4.5005
R64182 VINN.n232 VINN.n177 4.5005
R64183 VINN.n368 VINN.n177 4.5005
R64184 VINN.n231 VINN.n177 4.5005
R64185 VINN.n370 VINN.n177 4.5005
R64186 VINN.n230 VINN.n177 4.5005
R64187 VINN.n372 VINN.n177 4.5005
R64188 VINN.n229 VINN.n177 4.5005
R64189 VINN.n374 VINN.n177 4.5005
R64190 VINN.n228 VINN.n177 4.5005
R64191 VINN.n376 VINN.n177 4.5005
R64192 VINN.n227 VINN.n177 4.5005
R64193 VINN.n378 VINN.n177 4.5005
R64194 VINN.n226 VINN.n177 4.5005
R64195 VINN.n380 VINN.n177 4.5005
R64196 VINN.n225 VINN.n177 4.5005
R64197 VINN.n382 VINN.n177 4.5005
R64198 VINN.n224 VINN.n177 4.5005
R64199 VINN.n384 VINN.n177 4.5005
R64200 VINN.n223 VINN.n177 4.5005
R64201 VINN.n386 VINN.n177 4.5005
R64202 VINN.n222 VINN.n177 4.5005
R64203 VINN.n388 VINN.n177 4.5005
R64204 VINN.n221 VINN.n177 4.5005
R64205 VINN.n390 VINN.n177 4.5005
R64206 VINN.n220 VINN.n177 4.5005
R64207 VINN.n392 VINN.n177 4.5005
R64208 VINN.n219 VINN.n177 4.5005
R64209 VINN.n394 VINN.n177 4.5005
R64210 VINN.n218 VINN.n177 4.5005
R64211 VINN.n396 VINN.n177 4.5005
R64212 VINN.n217 VINN.n177 4.5005
R64213 VINN.n398 VINN.n177 4.5005
R64214 VINN.n216 VINN.n177 4.5005
R64215 VINN.n400 VINN.n177 4.5005
R64216 VINN.n215 VINN.n177 4.5005
R64217 VINN.n654 VINN.n177 4.5005
R64218 VINN.n656 VINN.n177 4.5005
R64219 VINN.n177 VINN.n0 4.5005
R64220 VINN.n278 VINN.n123 4.5005
R64221 VINN.n276 VINN.n123 4.5005
R64222 VINN.n280 VINN.n123 4.5005
R64223 VINN.n275 VINN.n123 4.5005
R64224 VINN.n282 VINN.n123 4.5005
R64225 VINN.n274 VINN.n123 4.5005
R64226 VINN.n284 VINN.n123 4.5005
R64227 VINN.n273 VINN.n123 4.5005
R64228 VINN.n286 VINN.n123 4.5005
R64229 VINN.n272 VINN.n123 4.5005
R64230 VINN.n288 VINN.n123 4.5005
R64231 VINN.n271 VINN.n123 4.5005
R64232 VINN.n290 VINN.n123 4.5005
R64233 VINN.n270 VINN.n123 4.5005
R64234 VINN.n292 VINN.n123 4.5005
R64235 VINN.n269 VINN.n123 4.5005
R64236 VINN.n294 VINN.n123 4.5005
R64237 VINN.n268 VINN.n123 4.5005
R64238 VINN.n296 VINN.n123 4.5005
R64239 VINN.n267 VINN.n123 4.5005
R64240 VINN.n298 VINN.n123 4.5005
R64241 VINN.n266 VINN.n123 4.5005
R64242 VINN.n300 VINN.n123 4.5005
R64243 VINN.n265 VINN.n123 4.5005
R64244 VINN.n302 VINN.n123 4.5005
R64245 VINN.n264 VINN.n123 4.5005
R64246 VINN.n304 VINN.n123 4.5005
R64247 VINN.n263 VINN.n123 4.5005
R64248 VINN.n306 VINN.n123 4.5005
R64249 VINN.n262 VINN.n123 4.5005
R64250 VINN.n308 VINN.n123 4.5005
R64251 VINN.n261 VINN.n123 4.5005
R64252 VINN.n310 VINN.n123 4.5005
R64253 VINN.n260 VINN.n123 4.5005
R64254 VINN.n312 VINN.n123 4.5005
R64255 VINN.n259 VINN.n123 4.5005
R64256 VINN.n314 VINN.n123 4.5005
R64257 VINN.n258 VINN.n123 4.5005
R64258 VINN.n316 VINN.n123 4.5005
R64259 VINN.n257 VINN.n123 4.5005
R64260 VINN.n318 VINN.n123 4.5005
R64261 VINN.n256 VINN.n123 4.5005
R64262 VINN.n320 VINN.n123 4.5005
R64263 VINN.n255 VINN.n123 4.5005
R64264 VINN.n322 VINN.n123 4.5005
R64265 VINN.n254 VINN.n123 4.5005
R64266 VINN.n324 VINN.n123 4.5005
R64267 VINN.n253 VINN.n123 4.5005
R64268 VINN.n326 VINN.n123 4.5005
R64269 VINN.n252 VINN.n123 4.5005
R64270 VINN.n328 VINN.n123 4.5005
R64271 VINN.n251 VINN.n123 4.5005
R64272 VINN.n330 VINN.n123 4.5005
R64273 VINN.n250 VINN.n123 4.5005
R64274 VINN.n332 VINN.n123 4.5005
R64275 VINN.n249 VINN.n123 4.5005
R64276 VINN.n334 VINN.n123 4.5005
R64277 VINN.n248 VINN.n123 4.5005
R64278 VINN.n336 VINN.n123 4.5005
R64279 VINN.n247 VINN.n123 4.5005
R64280 VINN.n338 VINN.n123 4.5005
R64281 VINN.n246 VINN.n123 4.5005
R64282 VINN.n340 VINN.n123 4.5005
R64283 VINN.n245 VINN.n123 4.5005
R64284 VINN.n342 VINN.n123 4.5005
R64285 VINN.n244 VINN.n123 4.5005
R64286 VINN.n344 VINN.n123 4.5005
R64287 VINN.n243 VINN.n123 4.5005
R64288 VINN.n346 VINN.n123 4.5005
R64289 VINN.n242 VINN.n123 4.5005
R64290 VINN.n348 VINN.n123 4.5005
R64291 VINN.n241 VINN.n123 4.5005
R64292 VINN.n350 VINN.n123 4.5005
R64293 VINN.n240 VINN.n123 4.5005
R64294 VINN.n352 VINN.n123 4.5005
R64295 VINN.n239 VINN.n123 4.5005
R64296 VINN.n354 VINN.n123 4.5005
R64297 VINN.n238 VINN.n123 4.5005
R64298 VINN.n356 VINN.n123 4.5005
R64299 VINN.n237 VINN.n123 4.5005
R64300 VINN.n358 VINN.n123 4.5005
R64301 VINN.n236 VINN.n123 4.5005
R64302 VINN.n360 VINN.n123 4.5005
R64303 VINN.n235 VINN.n123 4.5005
R64304 VINN.n362 VINN.n123 4.5005
R64305 VINN.n234 VINN.n123 4.5005
R64306 VINN.n364 VINN.n123 4.5005
R64307 VINN.n233 VINN.n123 4.5005
R64308 VINN.n366 VINN.n123 4.5005
R64309 VINN.n232 VINN.n123 4.5005
R64310 VINN.n368 VINN.n123 4.5005
R64311 VINN.n231 VINN.n123 4.5005
R64312 VINN.n370 VINN.n123 4.5005
R64313 VINN.n230 VINN.n123 4.5005
R64314 VINN.n372 VINN.n123 4.5005
R64315 VINN.n229 VINN.n123 4.5005
R64316 VINN.n374 VINN.n123 4.5005
R64317 VINN.n228 VINN.n123 4.5005
R64318 VINN.n376 VINN.n123 4.5005
R64319 VINN.n227 VINN.n123 4.5005
R64320 VINN.n378 VINN.n123 4.5005
R64321 VINN.n226 VINN.n123 4.5005
R64322 VINN.n380 VINN.n123 4.5005
R64323 VINN.n225 VINN.n123 4.5005
R64324 VINN.n382 VINN.n123 4.5005
R64325 VINN.n224 VINN.n123 4.5005
R64326 VINN.n384 VINN.n123 4.5005
R64327 VINN.n223 VINN.n123 4.5005
R64328 VINN.n386 VINN.n123 4.5005
R64329 VINN.n222 VINN.n123 4.5005
R64330 VINN.n388 VINN.n123 4.5005
R64331 VINN.n221 VINN.n123 4.5005
R64332 VINN.n390 VINN.n123 4.5005
R64333 VINN.n220 VINN.n123 4.5005
R64334 VINN.n392 VINN.n123 4.5005
R64335 VINN.n219 VINN.n123 4.5005
R64336 VINN.n394 VINN.n123 4.5005
R64337 VINN.n218 VINN.n123 4.5005
R64338 VINN.n396 VINN.n123 4.5005
R64339 VINN.n217 VINN.n123 4.5005
R64340 VINN.n398 VINN.n123 4.5005
R64341 VINN.n216 VINN.n123 4.5005
R64342 VINN.n400 VINN.n123 4.5005
R64343 VINN.n215 VINN.n123 4.5005
R64344 VINN.n654 VINN.n123 4.5005
R64345 VINN.n656 VINN.n123 4.5005
R64346 VINN.n123 VINN.n0 4.5005
R64347 VINN.n278 VINN.n178 4.5005
R64348 VINN.n276 VINN.n178 4.5005
R64349 VINN.n280 VINN.n178 4.5005
R64350 VINN.n275 VINN.n178 4.5005
R64351 VINN.n282 VINN.n178 4.5005
R64352 VINN.n274 VINN.n178 4.5005
R64353 VINN.n284 VINN.n178 4.5005
R64354 VINN.n273 VINN.n178 4.5005
R64355 VINN.n286 VINN.n178 4.5005
R64356 VINN.n272 VINN.n178 4.5005
R64357 VINN.n288 VINN.n178 4.5005
R64358 VINN.n271 VINN.n178 4.5005
R64359 VINN.n290 VINN.n178 4.5005
R64360 VINN.n270 VINN.n178 4.5005
R64361 VINN.n292 VINN.n178 4.5005
R64362 VINN.n269 VINN.n178 4.5005
R64363 VINN.n294 VINN.n178 4.5005
R64364 VINN.n268 VINN.n178 4.5005
R64365 VINN.n296 VINN.n178 4.5005
R64366 VINN.n267 VINN.n178 4.5005
R64367 VINN.n298 VINN.n178 4.5005
R64368 VINN.n266 VINN.n178 4.5005
R64369 VINN.n300 VINN.n178 4.5005
R64370 VINN.n265 VINN.n178 4.5005
R64371 VINN.n302 VINN.n178 4.5005
R64372 VINN.n264 VINN.n178 4.5005
R64373 VINN.n304 VINN.n178 4.5005
R64374 VINN.n263 VINN.n178 4.5005
R64375 VINN.n306 VINN.n178 4.5005
R64376 VINN.n262 VINN.n178 4.5005
R64377 VINN.n308 VINN.n178 4.5005
R64378 VINN.n261 VINN.n178 4.5005
R64379 VINN.n310 VINN.n178 4.5005
R64380 VINN.n260 VINN.n178 4.5005
R64381 VINN.n312 VINN.n178 4.5005
R64382 VINN.n259 VINN.n178 4.5005
R64383 VINN.n314 VINN.n178 4.5005
R64384 VINN.n258 VINN.n178 4.5005
R64385 VINN.n316 VINN.n178 4.5005
R64386 VINN.n257 VINN.n178 4.5005
R64387 VINN.n318 VINN.n178 4.5005
R64388 VINN.n256 VINN.n178 4.5005
R64389 VINN.n320 VINN.n178 4.5005
R64390 VINN.n255 VINN.n178 4.5005
R64391 VINN.n322 VINN.n178 4.5005
R64392 VINN.n254 VINN.n178 4.5005
R64393 VINN.n324 VINN.n178 4.5005
R64394 VINN.n253 VINN.n178 4.5005
R64395 VINN.n326 VINN.n178 4.5005
R64396 VINN.n252 VINN.n178 4.5005
R64397 VINN.n328 VINN.n178 4.5005
R64398 VINN.n251 VINN.n178 4.5005
R64399 VINN.n330 VINN.n178 4.5005
R64400 VINN.n250 VINN.n178 4.5005
R64401 VINN.n332 VINN.n178 4.5005
R64402 VINN.n249 VINN.n178 4.5005
R64403 VINN.n334 VINN.n178 4.5005
R64404 VINN.n248 VINN.n178 4.5005
R64405 VINN.n336 VINN.n178 4.5005
R64406 VINN.n247 VINN.n178 4.5005
R64407 VINN.n338 VINN.n178 4.5005
R64408 VINN.n246 VINN.n178 4.5005
R64409 VINN.n340 VINN.n178 4.5005
R64410 VINN.n245 VINN.n178 4.5005
R64411 VINN.n342 VINN.n178 4.5005
R64412 VINN.n244 VINN.n178 4.5005
R64413 VINN.n344 VINN.n178 4.5005
R64414 VINN.n243 VINN.n178 4.5005
R64415 VINN.n346 VINN.n178 4.5005
R64416 VINN.n242 VINN.n178 4.5005
R64417 VINN.n348 VINN.n178 4.5005
R64418 VINN.n241 VINN.n178 4.5005
R64419 VINN.n350 VINN.n178 4.5005
R64420 VINN.n240 VINN.n178 4.5005
R64421 VINN.n352 VINN.n178 4.5005
R64422 VINN.n239 VINN.n178 4.5005
R64423 VINN.n354 VINN.n178 4.5005
R64424 VINN.n238 VINN.n178 4.5005
R64425 VINN.n356 VINN.n178 4.5005
R64426 VINN.n237 VINN.n178 4.5005
R64427 VINN.n358 VINN.n178 4.5005
R64428 VINN.n236 VINN.n178 4.5005
R64429 VINN.n360 VINN.n178 4.5005
R64430 VINN.n235 VINN.n178 4.5005
R64431 VINN.n362 VINN.n178 4.5005
R64432 VINN.n234 VINN.n178 4.5005
R64433 VINN.n364 VINN.n178 4.5005
R64434 VINN.n233 VINN.n178 4.5005
R64435 VINN.n366 VINN.n178 4.5005
R64436 VINN.n232 VINN.n178 4.5005
R64437 VINN.n368 VINN.n178 4.5005
R64438 VINN.n231 VINN.n178 4.5005
R64439 VINN.n370 VINN.n178 4.5005
R64440 VINN.n230 VINN.n178 4.5005
R64441 VINN.n372 VINN.n178 4.5005
R64442 VINN.n229 VINN.n178 4.5005
R64443 VINN.n374 VINN.n178 4.5005
R64444 VINN.n228 VINN.n178 4.5005
R64445 VINN.n376 VINN.n178 4.5005
R64446 VINN.n227 VINN.n178 4.5005
R64447 VINN.n378 VINN.n178 4.5005
R64448 VINN.n226 VINN.n178 4.5005
R64449 VINN.n380 VINN.n178 4.5005
R64450 VINN.n225 VINN.n178 4.5005
R64451 VINN.n382 VINN.n178 4.5005
R64452 VINN.n224 VINN.n178 4.5005
R64453 VINN.n384 VINN.n178 4.5005
R64454 VINN.n223 VINN.n178 4.5005
R64455 VINN.n386 VINN.n178 4.5005
R64456 VINN.n222 VINN.n178 4.5005
R64457 VINN.n388 VINN.n178 4.5005
R64458 VINN.n221 VINN.n178 4.5005
R64459 VINN.n390 VINN.n178 4.5005
R64460 VINN.n220 VINN.n178 4.5005
R64461 VINN.n392 VINN.n178 4.5005
R64462 VINN.n219 VINN.n178 4.5005
R64463 VINN.n394 VINN.n178 4.5005
R64464 VINN.n218 VINN.n178 4.5005
R64465 VINN.n396 VINN.n178 4.5005
R64466 VINN.n217 VINN.n178 4.5005
R64467 VINN.n398 VINN.n178 4.5005
R64468 VINN.n216 VINN.n178 4.5005
R64469 VINN.n400 VINN.n178 4.5005
R64470 VINN.n215 VINN.n178 4.5005
R64471 VINN.n654 VINN.n178 4.5005
R64472 VINN.n656 VINN.n178 4.5005
R64473 VINN.n178 VINN.n0 4.5005
R64474 VINN.n278 VINN.n122 4.5005
R64475 VINN.n276 VINN.n122 4.5005
R64476 VINN.n280 VINN.n122 4.5005
R64477 VINN.n275 VINN.n122 4.5005
R64478 VINN.n282 VINN.n122 4.5005
R64479 VINN.n274 VINN.n122 4.5005
R64480 VINN.n284 VINN.n122 4.5005
R64481 VINN.n273 VINN.n122 4.5005
R64482 VINN.n286 VINN.n122 4.5005
R64483 VINN.n272 VINN.n122 4.5005
R64484 VINN.n288 VINN.n122 4.5005
R64485 VINN.n271 VINN.n122 4.5005
R64486 VINN.n290 VINN.n122 4.5005
R64487 VINN.n270 VINN.n122 4.5005
R64488 VINN.n292 VINN.n122 4.5005
R64489 VINN.n269 VINN.n122 4.5005
R64490 VINN.n294 VINN.n122 4.5005
R64491 VINN.n268 VINN.n122 4.5005
R64492 VINN.n296 VINN.n122 4.5005
R64493 VINN.n267 VINN.n122 4.5005
R64494 VINN.n298 VINN.n122 4.5005
R64495 VINN.n266 VINN.n122 4.5005
R64496 VINN.n300 VINN.n122 4.5005
R64497 VINN.n265 VINN.n122 4.5005
R64498 VINN.n302 VINN.n122 4.5005
R64499 VINN.n264 VINN.n122 4.5005
R64500 VINN.n304 VINN.n122 4.5005
R64501 VINN.n263 VINN.n122 4.5005
R64502 VINN.n306 VINN.n122 4.5005
R64503 VINN.n262 VINN.n122 4.5005
R64504 VINN.n308 VINN.n122 4.5005
R64505 VINN.n261 VINN.n122 4.5005
R64506 VINN.n310 VINN.n122 4.5005
R64507 VINN.n260 VINN.n122 4.5005
R64508 VINN.n312 VINN.n122 4.5005
R64509 VINN.n259 VINN.n122 4.5005
R64510 VINN.n314 VINN.n122 4.5005
R64511 VINN.n258 VINN.n122 4.5005
R64512 VINN.n316 VINN.n122 4.5005
R64513 VINN.n257 VINN.n122 4.5005
R64514 VINN.n318 VINN.n122 4.5005
R64515 VINN.n256 VINN.n122 4.5005
R64516 VINN.n320 VINN.n122 4.5005
R64517 VINN.n255 VINN.n122 4.5005
R64518 VINN.n322 VINN.n122 4.5005
R64519 VINN.n254 VINN.n122 4.5005
R64520 VINN.n324 VINN.n122 4.5005
R64521 VINN.n253 VINN.n122 4.5005
R64522 VINN.n326 VINN.n122 4.5005
R64523 VINN.n252 VINN.n122 4.5005
R64524 VINN.n328 VINN.n122 4.5005
R64525 VINN.n251 VINN.n122 4.5005
R64526 VINN.n330 VINN.n122 4.5005
R64527 VINN.n250 VINN.n122 4.5005
R64528 VINN.n332 VINN.n122 4.5005
R64529 VINN.n249 VINN.n122 4.5005
R64530 VINN.n334 VINN.n122 4.5005
R64531 VINN.n248 VINN.n122 4.5005
R64532 VINN.n336 VINN.n122 4.5005
R64533 VINN.n247 VINN.n122 4.5005
R64534 VINN.n338 VINN.n122 4.5005
R64535 VINN.n246 VINN.n122 4.5005
R64536 VINN.n340 VINN.n122 4.5005
R64537 VINN.n245 VINN.n122 4.5005
R64538 VINN.n342 VINN.n122 4.5005
R64539 VINN.n244 VINN.n122 4.5005
R64540 VINN.n344 VINN.n122 4.5005
R64541 VINN.n243 VINN.n122 4.5005
R64542 VINN.n346 VINN.n122 4.5005
R64543 VINN.n242 VINN.n122 4.5005
R64544 VINN.n348 VINN.n122 4.5005
R64545 VINN.n241 VINN.n122 4.5005
R64546 VINN.n350 VINN.n122 4.5005
R64547 VINN.n240 VINN.n122 4.5005
R64548 VINN.n352 VINN.n122 4.5005
R64549 VINN.n239 VINN.n122 4.5005
R64550 VINN.n354 VINN.n122 4.5005
R64551 VINN.n238 VINN.n122 4.5005
R64552 VINN.n356 VINN.n122 4.5005
R64553 VINN.n237 VINN.n122 4.5005
R64554 VINN.n358 VINN.n122 4.5005
R64555 VINN.n236 VINN.n122 4.5005
R64556 VINN.n360 VINN.n122 4.5005
R64557 VINN.n235 VINN.n122 4.5005
R64558 VINN.n362 VINN.n122 4.5005
R64559 VINN.n234 VINN.n122 4.5005
R64560 VINN.n364 VINN.n122 4.5005
R64561 VINN.n233 VINN.n122 4.5005
R64562 VINN.n366 VINN.n122 4.5005
R64563 VINN.n232 VINN.n122 4.5005
R64564 VINN.n368 VINN.n122 4.5005
R64565 VINN.n231 VINN.n122 4.5005
R64566 VINN.n370 VINN.n122 4.5005
R64567 VINN.n230 VINN.n122 4.5005
R64568 VINN.n372 VINN.n122 4.5005
R64569 VINN.n229 VINN.n122 4.5005
R64570 VINN.n374 VINN.n122 4.5005
R64571 VINN.n228 VINN.n122 4.5005
R64572 VINN.n376 VINN.n122 4.5005
R64573 VINN.n227 VINN.n122 4.5005
R64574 VINN.n378 VINN.n122 4.5005
R64575 VINN.n226 VINN.n122 4.5005
R64576 VINN.n380 VINN.n122 4.5005
R64577 VINN.n225 VINN.n122 4.5005
R64578 VINN.n382 VINN.n122 4.5005
R64579 VINN.n224 VINN.n122 4.5005
R64580 VINN.n384 VINN.n122 4.5005
R64581 VINN.n223 VINN.n122 4.5005
R64582 VINN.n386 VINN.n122 4.5005
R64583 VINN.n222 VINN.n122 4.5005
R64584 VINN.n388 VINN.n122 4.5005
R64585 VINN.n221 VINN.n122 4.5005
R64586 VINN.n390 VINN.n122 4.5005
R64587 VINN.n220 VINN.n122 4.5005
R64588 VINN.n392 VINN.n122 4.5005
R64589 VINN.n219 VINN.n122 4.5005
R64590 VINN.n394 VINN.n122 4.5005
R64591 VINN.n218 VINN.n122 4.5005
R64592 VINN.n396 VINN.n122 4.5005
R64593 VINN.n217 VINN.n122 4.5005
R64594 VINN.n398 VINN.n122 4.5005
R64595 VINN.n216 VINN.n122 4.5005
R64596 VINN.n400 VINN.n122 4.5005
R64597 VINN.n215 VINN.n122 4.5005
R64598 VINN.n654 VINN.n122 4.5005
R64599 VINN.n656 VINN.n122 4.5005
R64600 VINN.n122 VINN.n0 4.5005
R64601 VINN.n278 VINN.n179 4.5005
R64602 VINN.n276 VINN.n179 4.5005
R64603 VINN.n280 VINN.n179 4.5005
R64604 VINN.n275 VINN.n179 4.5005
R64605 VINN.n282 VINN.n179 4.5005
R64606 VINN.n274 VINN.n179 4.5005
R64607 VINN.n284 VINN.n179 4.5005
R64608 VINN.n273 VINN.n179 4.5005
R64609 VINN.n286 VINN.n179 4.5005
R64610 VINN.n272 VINN.n179 4.5005
R64611 VINN.n288 VINN.n179 4.5005
R64612 VINN.n271 VINN.n179 4.5005
R64613 VINN.n290 VINN.n179 4.5005
R64614 VINN.n270 VINN.n179 4.5005
R64615 VINN.n292 VINN.n179 4.5005
R64616 VINN.n269 VINN.n179 4.5005
R64617 VINN.n294 VINN.n179 4.5005
R64618 VINN.n268 VINN.n179 4.5005
R64619 VINN.n296 VINN.n179 4.5005
R64620 VINN.n267 VINN.n179 4.5005
R64621 VINN.n298 VINN.n179 4.5005
R64622 VINN.n266 VINN.n179 4.5005
R64623 VINN.n300 VINN.n179 4.5005
R64624 VINN.n265 VINN.n179 4.5005
R64625 VINN.n302 VINN.n179 4.5005
R64626 VINN.n264 VINN.n179 4.5005
R64627 VINN.n304 VINN.n179 4.5005
R64628 VINN.n263 VINN.n179 4.5005
R64629 VINN.n306 VINN.n179 4.5005
R64630 VINN.n262 VINN.n179 4.5005
R64631 VINN.n308 VINN.n179 4.5005
R64632 VINN.n261 VINN.n179 4.5005
R64633 VINN.n310 VINN.n179 4.5005
R64634 VINN.n260 VINN.n179 4.5005
R64635 VINN.n312 VINN.n179 4.5005
R64636 VINN.n259 VINN.n179 4.5005
R64637 VINN.n314 VINN.n179 4.5005
R64638 VINN.n258 VINN.n179 4.5005
R64639 VINN.n316 VINN.n179 4.5005
R64640 VINN.n257 VINN.n179 4.5005
R64641 VINN.n318 VINN.n179 4.5005
R64642 VINN.n256 VINN.n179 4.5005
R64643 VINN.n320 VINN.n179 4.5005
R64644 VINN.n255 VINN.n179 4.5005
R64645 VINN.n322 VINN.n179 4.5005
R64646 VINN.n254 VINN.n179 4.5005
R64647 VINN.n324 VINN.n179 4.5005
R64648 VINN.n253 VINN.n179 4.5005
R64649 VINN.n326 VINN.n179 4.5005
R64650 VINN.n252 VINN.n179 4.5005
R64651 VINN.n328 VINN.n179 4.5005
R64652 VINN.n251 VINN.n179 4.5005
R64653 VINN.n330 VINN.n179 4.5005
R64654 VINN.n250 VINN.n179 4.5005
R64655 VINN.n332 VINN.n179 4.5005
R64656 VINN.n249 VINN.n179 4.5005
R64657 VINN.n334 VINN.n179 4.5005
R64658 VINN.n248 VINN.n179 4.5005
R64659 VINN.n336 VINN.n179 4.5005
R64660 VINN.n247 VINN.n179 4.5005
R64661 VINN.n338 VINN.n179 4.5005
R64662 VINN.n246 VINN.n179 4.5005
R64663 VINN.n340 VINN.n179 4.5005
R64664 VINN.n245 VINN.n179 4.5005
R64665 VINN.n342 VINN.n179 4.5005
R64666 VINN.n244 VINN.n179 4.5005
R64667 VINN.n344 VINN.n179 4.5005
R64668 VINN.n243 VINN.n179 4.5005
R64669 VINN.n346 VINN.n179 4.5005
R64670 VINN.n242 VINN.n179 4.5005
R64671 VINN.n348 VINN.n179 4.5005
R64672 VINN.n241 VINN.n179 4.5005
R64673 VINN.n350 VINN.n179 4.5005
R64674 VINN.n240 VINN.n179 4.5005
R64675 VINN.n352 VINN.n179 4.5005
R64676 VINN.n239 VINN.n179 4.5005
R64677 VINN.n354 VINN.n179 4.5005
R64678 VINN.n238 VINN.n179 4.5005
R64679 VINN.n356 VINN.n179 4.5005
R64680 VINN.n237 VINN.n179 4.5005
R64681 VINN.n358 VINN.n179 4.5005
R64682 VINN.n236 VINN.n179 4.5005
R64683 VINN.n360 VINN.n179 4.5005
R64684 VINN.n235 VINN.n179 4.5005
R64685 VINN.n362 VINN.n179 4.5005
R64686 VINN.n234 VINN.n179 4.5005
R64687 VINN.n364 VINN.n179 4.5005
R64688 VINN.n233 VINN.n179 4.5005
R64689 VINN.n366 VINN.n179 4.5005
R64690 VINN.n232 VINN.n179 4.5005
R64691 VINN.n368 VINN.n179 4.5005
R64692 VINN.n231 VINN.n179 4.5005
R64693 VINN.n370 VINN.n179 4.5005
R64694 VINN.n230 VINN.n179 4.5005
R64695 VINN.n372 VINN.n179 4.5005
R64696 VINN.n229 VINN.n179 4.5005
R64697 VINN.n374 VINN.n179 4.5005
R64698 VINN.n228 VINN.n179 4.5005
R64699 VINN.n376 VINN.n179 4.5005
R64700 VINN.n227 VINN.n179 4.5005
R64701 VINN.n378 VINN.n179 4.5005
R64702 VINN.n226 VINN.n179 4.5005
R64703 VINN.n380 VINN.n179 4.5005
R64704 VINN.n225 VINN.n179 4.5005
R64705 VINN.n382 VINN.n179 4.5005
R64706 VINN.n224 VINN.n179 4.5005
R64707 VINN.n384 VINN.n179 4.5005
R64708 VINN.n223 VINN.n179 4.5005
R64709 VINN.n386 VINN.n179 4.5005
R64710 VINN.n222 VINN.n179 4.5005
R64711 VINN.n388 VINN.n179 4.5005
R64712 VINN.n221 VINN.n179 4.5005
R64713 VINN.n390 VINN.n179 4.5005
R64714 VINN.n220 VINN.n179 4.5005
R64715 VINN.n392 VINN.n179 4.5005
R64716 VINN.n219 VINN.n179 4.5005
R64717 VINN.n394 VINN.n179 4.5005
R64718 VINN.n218 VINN.n179 4.5005
R64719 VINN.n396 VINN.n179 4.5005
R64720 VINN.n217 VINN.n179 4.5005
R64721 VINN.n398 VINN.n179 4.5005
R64722 VINN.n216 VINN.n179 4.5005
R64723 VINN.n400 VINN.n179 4.5005
R64724 VINN.n215 VINN.n179 4.5005
R64725 VINN.n654 VINN.n179 4.5005
R64726 VINN.n656 VINN.n179 4.5005
R64727 VINN.n179 VINN.n0 4.5005
R64728 VINN.n278 VINN.n121 4.5005
R64729 VINN.n276 VINN.n121 4.5005
R64730 VINN.n280 VINN.n121 4.5005
R64731 VINN.n275 VINN.n121 4.5005
R64732 VINN.n282 VINN.n121 4.5005
R64733 VINN.n274 VINN.n121 4.5005
R64734 VINN.n284 VINN.n121 4.5005
R64735 VINN.n273 VINN.n121 4.5005
R64736 VINN.n286 VINN.n121 4.5005
R64737 VINN.n272 VINN.n121 4.5005
R64738 VINN.n288 VINN.n121 4.5005
R64739 VINN.n271 VINN.n121 4.5005
R64740 VINN.n290 VINN.n121 4.5005
R64741 VINN.n270 VINN.n121 4.5005
R64742 VINN.n292 VINN.n121 4.5005
R64743 VINN.n269 VINN.n121 4.5005
R64744 VINN.n294 VINN.n121 4.5005
R64745 VINN.n268 VINN.n121 4.5005
R64746 VINN.n296 VINN.n121 4.5005
R64747 VINN.n267 VINN.n121 4.5005
R64748 VINN.n298 VINN.n121 4.5005
R64749 VINN.n266 VINN.n121 4.5005
R64750 VINN.n300 VINN.n121 4.5005
R64751 VINN.n265 VINN.n121 4.5005
R64752 VINN.n302 VINN.n121 4.5005
R64753 VINN.n264 VINN.n121 4.5005
R64754 VINN.n304 VINN.n121 4.5005
R64755 VINN.n263 VINN.n121 4.5005
R64756 VINN.n306 VINN.n121 4.5005
R64757 VINN.n262 VINN.n121 4.5005
R64758 VINN.n308 VINN.n121 4.5005
R64759 VINN.n261 VINN.n121 4.5005
R64760 VINN.n310 VINN.n121 4.5005
R64761 VINN.n260 VINN.n121 4.5005
R64762 VINN.n312 VINN.n121 4.5005
R64763 VINN.n259 VINN.n121 4.5005
R64764 VINN.n314 VINN.n121 4.5005
R64765 VINN.n258 VINN.n121 4.5005
R64766 VINN.n316 VINN.n121 4.5005
R64767 VINN.n257 VINN.n121 4.5005
R64768 VINN.n318 VINN.n121 4.5005
R64769 VINN.n256 VINN.n121 4.5005
R64770 VINN.n320 VINN.n121 4.5005
R64771 VINN.n255 VINN.n121 4.5005
R64772 VINN.n322 VINN.n121 4.5005
R64773 VINN.n254 VINN.n121 4.5005
R64774 VINN.n324 VINN.n121 4.5005
R64775 VINN.n253 VINN.n121 4.5005
R64776 VINN.n326 VINN.n121 4.5005
R64777 VINN.n252 VINN.n121 4.5005
R64778 VINN.n328 VINN.n121 4.5005
R64779 VINN.n251 VINN.n121 4.5005
R64780 VINN.n330 VINN.n121 4.5005
R64781 VINN.n250 VINN.n121 4.5005
R64782 VINN.n332 VINN.n121 4.5005
R64783 VINN.n249 VINN.n121 4.5005
R64784 VINN.n334 VINN.n121 4.5005
R64785 VINN.n248 VINN.n121 4.5005
R64786 VINN.n336 VINN.n121 4.5005
R64787 VINN.n247 VINN.n121 4.5005
R64788 VINN.n338 VINN.n121 4.5005
R64789 VINN.n246 VINN.n121 4.5005
R64790 VINN.n340 VINN.n121 4.5005
R64791 VINN.n245 VINN.n121 4.5005
R64792 VINN.n342 VINN.n121 4.5005
R64793 VINN.n244 VINN.n121 4.5005
R64794 VINN.n344 VINN.n121 4.5005
R64795 VINN.n243 VINN.n121 4.5005
R64796 VINN.n346 VINN.n121 4.5005
R64797 VINN.n242 VINN.n121 4.5005
R64798 VINN.n348 VINN.n121 4.5005
R64799 VINN.n241 VINN.n121 4.5005
R64800 VINN.n350 VINN.n121 4.5005
R64801 VINN.n240 VINN.n121 4.5005
R64802 VINN.n352 VINN.n121 4.5005
R64803 VINN.n239 VINN.n121 4.5005
R64804 VINN.n354 VINN.n121 4.5005
R64805 VINN.n238 VINN.n121 4.5005
R64806 VINN.n356 VINN.n121 4.5005
R64807 VINN.n237 VINN.n121 4.5005
R64808 VINN.n358 VINN.n121 4.5005
R64809 VINN.n236 VINN.n121 4.5005
R64810 VINN.n360 VINN.n121 4.5005
R64811 VINN.n235 VINN.n121 4.5005
R64812 VINN.n362 VINN.n121 4.5005
R64813 VINN.n234 VINN.n121 4.5005
R64814 VINN.n364 VINN.n121 4.5005
R64815 VINN.n233 VINN.n121 4.5005
R64816 VINN.n366 VINN.n121 4.5005
R64817 VINN.n232 VINN.n121 4.5005
R64818 VINN.n368 VINN.n121 4.5005
R64819 VINN.n231 VINN.n121 4.5005
R64820 VINN.n370 VINN.n121 4.5005
R64821 VINN.n230 VINN.n121 4.5005
R64822 VINN.n372 VINN.n121 4.5005
R64823 VINN.n229 VINN.n121 4.5005
R64824 VINN.n374 VINN.n121 4.5005
R64825 VINN.n228 VINN.n121 4.5005
R64826 VINN.n376 VINN.n121 4.5005
R64827 VINN.n227 VINN.n121 4.5005
R64828 VINN.n378 VINN.n121 4.5005
R64829 VINN.n226 VINN.n121 4.5005
R64830 VINN.n380 VINN.n121 4.5005
R64831 VINN.n225 VINN.n121 4.5005
R64832 VINN.n382 VINN.n121 4.5005
R64833 VINN.n224 VINN.n121 4.5005
R64834 VINN.n384 VINN.n121 4.5005
R64835 VINN.n223 VINN.n121 4.5005
R64836 VINN.n386 VINN.n121 4.5005
R64837 VINN.n222 VINN.n121 4.5005
R64838 VINN.n388 VINN.n121 4.5005
R64839 VINN.n221 VINN.n121 4.5005
R64840 VINN.n390 VINN.n121 4.5005
R64841 VINN.n220 VINN.n121 4.5005
R64842 VINN.n392 VINN.n121 4.5005
R64843 VINN.n219 VINN.n121 4.5005
R64844 VINN.n394 VINN.n121 4.5005
R64845 VINN.n218 VINN.n121 4.5005
R64846 VINN.n396 VINN.n121 4.5005
R64847 VINN.n217 VINN.n121 4.5005
R64848 VINN.n398 VINN.n121 4.5005
R64849 VINN.n216 VINN.n121 4.5005
R64850 VINN.n400 VINN.n121 4.5005
R64851 VINN.n215 VINN.n121 4.5005
R64852 VINN.n654 VINN.n121 4.5005
R64853 VINN.n656 VINN.n121 4.5005
R64854 VINN.n121 VINN.n0 4.5005
R64855 VINN.n278 VINN.n180 4.5005
R64856 VINN.n276 VINN.n180 4.5005
R64857 VINN.n280 VINN.n180 4.5005
R64858 VINN.n275 VINN.n180 4.5005
R64859 VINN.n282 VINN.n180 4.5005
R64860 VINN.n274 VINN.n180 4.5005
R64861 VINN.n284 VINN.n180 4.5005
R64862 VINN.n273 VINN.n180 4.5005
R64863 VINN.n286 VINN.n180 4.5005
R64864 VINN.n272 VINN.n180 4.5005
R64865 VINN.n288 VINN.n180 4.5005
R64866 VINN.n271 VINN.n180 4.5005
R64867 VINN.n290 VINN.n180 4.5005
R64868 VINN.n270 VINN.n180 4.5005
R64869 VINN.n292 VINN.n180 4.5005
R64870 VINN.n269 VINN.n180 4.5005
R64871 VINN.n294 VINN.n180 4.5005
R64872 VINN.n268 VINN.n180 4.5005
R64873 VINN.n296 VINN.n180 4.5005
R64874 VINN.n267 VINN.n180 4.5005
R64875 VINN.n298 VINN.n180 4.5005
R64876 VINN.n266 VINN.n180 4.5005
R64877 VINN.n300 VINN.n180 4.5005
R64878 VINN.n265 VINN.n180 4.5005
R64879 VINN.n302 VINN.n180 4.5005
R64880 VINN.n264 VINN.n180 4.5005
R64881 VINN.n304 VINN.n180 4.5005
R64882 VINN.n263 VINN.n180 4.5005
R64883 VINN.n306 VINN.n180 4.5005
R64884 VINN.n262 VINN.n180 4.5005
R64885 VINN.n308 VINN.n180 4.5005
R64886 VINN.n261 VINN.n180 4.5005
R64887 VINN.n310 VINN.n180 4.5005
R64888 VINN.n260 VINN.n180 4.5005
R64889 VINN.n312 VINN.n180 4.5005
R64890 VINN.n259 VINN.n180 4.5005
R64891 VINN.n314 VINN.n180 4.5005
R64892 VINN.n258 VINN.n180 4.5005
R64893 VINN.n316 VINN.n180 4.5005
R64894 VINN.n257 VINN.n180 4.5005
R64895 VINN.n318 VINN.n180 4.5005
R64896 VINN.n256 VINN.n180 4.5005
R64897 VINN.n320 VINN.n180 4.5005
R64898 VINN.n255 VINN.n180 4.5005
R64899 VINN.n322 VINN.n180 4.5005
R64900 VINN.n254 VINN.n180 4.5005
R64901 VINN.n324 VINN.n180 4.5005
R64902 VINN.n253 VINN.n180 4.5005
R64903 VINN.n326 VINN.n180 4.5005
R64904 VINN.n252 VINN.n180 4.5005
R64905 VINN.n328 VINN.n180 4.5005
R64906 VINN.n251 VINN.n180 4.5005
R64907 VINN.n330 VINN.n180 4.5005
R64908 VINN.n250 VINN.n180 4.5005
R64909 VINN.n332 VINN.n180 4.5005
R64910 VINN.n249 VINN.n180 4.5005
R64911 VINN.n334 VINN.n180 4.5005
R64912 VINN.n248 VINN.n180 4.5005
R64913 VINN.n336 VINN.n180 4.5005
R64914 VINN.n247 VINN.n180 4.5005
R64915 VINN.n338 VINN.n180 4.5005
R64916 VINN.n246 VINN.n180 4.5005
R64917 VINN.n340 VINN.n180 4.5005
R64918 VINN.n245 VINN.n180 4.5005
R64919 VINN.n342 VINN.n180 4.5005
R64920 VINN.n244 VINN.n180 4.5005
R64921 VINN.n344 VINN.n180 4.5005
R64922 VINN.n243 VINN.n180 4.5005
R64923 VINN.n346 VINN.n180 4.5005
R64924 VINN.n242 VINN.n180 4.5005
R64925 VINN.n348 VINN.n180 4.5005
R64926 VINN.n241 VINN.n180 4.5005
R64927 VINN.n350 VINN.n180 4.5005
R64928 VINN.n240 VINN.n180 4.5005
R64929 VINN.n352 VINN.n180 4.5005
R64930 VINN.n239 VINN.n180 4.5005
R64931 VINN.n354 VINN.n180 4.5005
R64932 VINN.n238 VINN.n180 4.5005
R64933 VINN.n356 VINN.n180 4.5005
R64934 VINN.n237 VINN.n180 4.5005
R64935 VINN.n358 VINN.n180 4.5005
R64936 VINN.n236 VINN.n180 4.5005
R64937 VINN.n360 VINN.n180 4.5005
R64938 VINN.n235 VINN.n180 4.5005
R64939 VINN.n362 VINN.n180 4.5005
R64940 VINN.n234 VINN.n180 4.5005
R64941 VINN.n364 VINN.n180 4.5005
R64942 VINN.n233 VINN.n180 4.5005
R64943 VINN.n366 VINN.n180 4.5005
R64944 VINN.n232 VINN.n180 4.5005
R64945 VINN.n368 VINN.n180 4.5005
R64946 VINN.n231 VINN.n180 4.5005
R64947 VINN.n370 VINN.n180 4.5005
R64948 VINN.n230 VINN.n180 4.5005
R64949 VINN.n372 VINN.n180 4.5005
R64950 VINN.n229 VINN.n180 4.5005
R64951 VINN.n374 VINN.n180 4.5005
R64952 VINN.n228 VINN.n180 4.5005
R64953 VINN.n376 VINN.n180 4.5005
R64954 VINN.n227 VINN.n180 4.5005
R64955 VINN.n378 VINN.n180 4.5005
R64956 VINN.n226 VINN.n180 4.5005
R64957 VINN.n380 VINN.n180 4.5005
R64958 VINN.n225 VINN.n180 4.5005
R64959 VINN.n382 VINN.n180 4.5005
R64960 VINN.n224 VINN.n180 4.5005
R64961 VINN.n384 VINN.n180 4.5005
R64962 VINN.n223 VINN.n180 4.5005
R64963 VINN.n386 VINN.n180 4.5005
R64964 VINN.n222 VINN.n180 4.5005
R64965 VINN.n388 VINN.n180 4.5005
R64966 VINN.n221 VINN.n180 4.5005
R64967 VINN.n390 VINN.n180 4.5005
R64968 VINN.n220 VINN.n180 4.5005
R64969 VINN.n392 VINN.n180 4.5005
R64970 VINN.n219 VINN.n180 4.5005
R64971 VINN.n394 VINN.n180 4.5005
R64972 VINN.n218 VINN.n180 4.5005
R64973 VINN.n396 VINN.n180 4.5005
R64974 VINN.n217 VINN.n180 4.5005
R64975 VINN.n398 VINN.n180 4.5005
R64976 VINN.n216 VINN.n180 4.5005
R64977 VINN.n400 VINN.n180 4.5005
R64978 VINN.n215 VINN.n180 4.5005
R64979 VINN.n654 VINN.n180 4.5005
R64980 VINN.n656 VINN.n180 4.5005
R64981 VINN.n180 VINN.n0 4.5005
R64982 VINN.n278 VINN.n120 4.5005
R64983 VINN.n276 VINN.n120 4.5005
R64984 VINN.n280 VINN.n120 4.5005
R64985 VINN.n275 VINN.n120 4.5005
R64986 VINN.n282 VINN.n120 4.5005
R64987 VINN.n274 VINN.n120 4.5005
R64988 VINN.n284 VINN.n120 4.5005
R64989 VINN.n273 VINN.n120 4.5005
R64990 VINN.n286 VINN.n120 4.5005
R64991 VINN.n272 VINN.n120 4.5005
R64992 VINN.n288 VINN.n120 4.5005
R64993 VINN.n271 VINN.n120 4.5005
R64994 VINN.n290 VINN.n120 4.5005
R64995 VINN.n270 VINN.n120 4.5005
R64996 VINN.n292 VINN.n120 4.5005
R64997 VINN.n269 VINN.n120 4.5005
R64998 VINN.n294 VINN.n120 4.5005
R64999 VINN.n268 VINN.n120 4.5005
R65000 VINN.n296 VINN.n120 4.5005
R65001 VINN.n267 VINN.n120 4.5005
R65002 VINN.n298 VINN.n120 4.5005
R65003 VINN.n266 VINN.n120 4.5005
R65004 VINN.n300 VINN.n120 4.5005
R65005 VINN.n265 VINN.n120 4.5005
R65006 VINN.n302 VINN.n120 4.5005
R65007 VINN.n264 VINN.n120 4.5005
R65008 VINN.n304 VINN.n120 4.5005
R65009 VINN.n263 VINN.n120 4.5005
R65010 VINN.n306 VINN.n120 4.5005
R65011 VINN.n262 VINN.n120 4.5005
R65012 VINN.n308 VINN.n120 4.5005
R65013 VINN.n261 VINN.n120 4.5005
R65014 VINN.n310 VINN.n120 4.5005
R65015 VINN.n260 VINN.n120 4.5005
R65016 VINN.n312 VINN.n120 4.5005
R65017 VINN.n259 VINN.n120 4.5005
R65018 VINN.n314 VINN.n120 4.5005
R65019 VINN.n258 VINN.n120 4.5005
R65020 VINN.n316 VINN.n120 4.5005
R65021 VINN.n257 VINN.n120 4.5005
R65022 VINN.n318 VINN.n120 4.5005
R65023 VINN.n256 VINN.n120 4.5005
R65024 VINN.n320 VINN.n120 4.5005
R65025 VINN.n255 VINN.n120 4.5005
R65026 VINN.n322 VINN.n120 4.5005
R65027 VINN.n254 VINN.n120 4.5005
R65028 VINN.n324 VINN.n120 4.5005
R65029 VINN.n253 VINN.n120 4.5005
R65030 VINN.n326 VINN.n120 4.5005
R65031 VINN.n252 VINN.n120 4.5005
R65032 VINN.n328 VINN.n120 4.5005
R65033 VINN.n251 VINN.n120 4.5005
R65034 VINN.n330 VINN.n120 4.5005
R65035 VINN.n250 VINN.n120 4.5005
R65036 VINN.n332 VINN.n120 4.5005
R65037 VINN.n249 VINN.n120 4.5005
R65038 VINN.n334 VINN.n120 4.5005
R65039 VINN.n248 VINN.n120 4.5005
R65040 VINN.n336 VINN.n120 4.5005
R65041 VINN.n247 VINN.n120 4.5005
R65042 VINN.n338 VINN.n120 4.5005
R65043 VINN.n246 VINN.n120 4.5005
R65044 VINN.n340 VINN.n120 4.5005
R65045 VINN.n245 VINN.n120 4.5005
R65046 VINN.n342 VINN.n120 4.5005
R65047 VINN.n244 VINN.n120 4.5005
R65048 VINN.n344 VINN.n120 4.5005
R65049 VINN.n243 VINN.n120 4.5005
R65050 VINN.n346 VINN.n120 4.5005
R65051 VINN.n242 VINN.n120 4.5005
R65052 VINN.n348 VINN.n120 4.5005
R65053 VINN.n241 VINN.n120 4.5005
R65054 VINN.n350 VINN.n120 4.5005
R65055 VINN.n240 VINN.n120 4.5005
R65056 VINN.n352 VINN.n120 4.5005
R65057 VINN.n239 VINN.n120 4.5005
R65058 VINN.n354 VINN.n120 4.5005
R65059 VINN.n238 VINN.n120 4.5005
R65060 VINN.n356 VINN.n120 4.5005
R65061 VINN.n237 VINN.n120 4.5005
R65062 VINN.n358 VINN.n120 4.5005
R65063 VINN.n236 VINN.n120 4.5005
R65064 VINN.n360 VINN.n120 4.5005
R65065 VINN.n235 VINN.n120 4.5005
R65066 VINN.n362 VINN.n120 4.5005
R65067 VINN.n234 VINN.n120 4.5005
R65068 VINN.n364 VINN.n120 4.5005
R65069 VINN.n233 VINN.n120 4.5005
R65070 VINN.n366 VINN.n120 4.5005
R65071 VINN.n232 VINN.n120 4.5005
R65072 VINN.n368 VINN.n120 4.5005
R65073 VINN.n231 VINN.n120 4.5005
R65074 VINN.n370 VINN.n120 4.5005
R65075 VINN.n230 VINN.n120 4.5005
R65076 VINN.n372 VINN.n120 4.5005
R65077 VINN.n229 VINN.n120 4.5005
R65078 VINN.n374 VINN.n120 4.5005
R65079 VINN.n228 VINN.n120 4.5005
R65080 VINN.n376 VINN.n120 4.5005
R65081 VINN.n227 VINN.n120 4.5005
R65082 VINN.n378 VINN.n120 4.5005
R65083 VINN.n226 VINN.n120 4.5005
R65084 VINN.n380 VINN.n120 4.5005
R65085 VINN.n225 VINN.n120 4.5005
R65086 VINN.n382 VINN.n120 4.5005
R65087 VINN.n224 VINN.n120 4.5005
R65088 VINN.n384 VINN.n120 4.5005
R65089 VINN.n223 VINN.n120 4.5005
R65090 VINN.n386 VINN.n120 4.5005
R65091 VINN.n222 VINN.n120 4.5005
R65092 VINN.n388 VINN.n120 4.5005
R65093 VINN.n221 VINN.n120 4.5005
R65094 VINN.n390 VINN.n120 4.5005
R65095 VINN.n220 VINN.n120 4.5005
R65096 VINN.n392 VINN.n120 4.5005
R65097 VINN.n219 VINN.n120 4.5005
R65098 VINN.n394 VINN.n120 4.5005
R65099 VINN.n218 VINN.n120 4.5005
R65100 VINN.n396 VINN.n120 4.5005
R65101 VINN.n217 VINN.n120 4.5005
R65102 VINN.n398 VINN.n120 4.5005
R65103 VINN.n216 VINN.n120 4.5005
R65104 VINN.n400 VINN.n120 4.5005
R65105 VINN.n215 VINN.n120 4.5005
R65106 VINN.n654 VINN.n120 4.5005
R65107 VINN.n656 VINN.n120 4.5005
R65108 VINN.n120 VINN.n0 4.5005
R65109 VINN.n278 VINN.n181 4.5005
R65110 VINN.n276 VINN.n181 4.5005
R65111 VINN.n280 VINN.n181 4.5005
R65112 VINN.n275 VINN.n181 4.5005
R65113 VINN.n282 VINN.n181 4.5005
R65114 VINN.n274 VINN.n181 4.5005
R65115 VINN.n284 VINN.n181 4.5005
R65116 VINN.n273 VINN.n181 4.5005
R65117 VINN.n286 VINN.n181 4.5005
R65118 VINN.n272 VINN.n181 4.5005
R65119 VINN.n288 VINN.n181 4.5005
R65120 VINN.n271 VINN.n181 4.5005
R65121 VINN.n290 VINN.n181 4.5005
R65122 VINN.n270 VINN.n181 4.5005
R65123 VINN.n292 VINN.n181 4.5005
R65124 VINN.n269 VINN.n181 4.5005
R65125 VINN.n294 VINN.n181 4.5005
R65126 VINN.n268 VINN.n181 4.5005
R65127 VINN.n296 VINN.n181 4.5005
R65128 VINN.n267 VINN.n181 4.5005
R65129 VINN.n298 VINN.n181 4.5005
R65130 VINN.n266 VINN.n181 4.5005
R65131 VINN.n300 VINN.n181 4.5005
R65132 VINN.n265 VINN.n181 4.5005
R65133 VINN.n302 VINN.n181 4.5005
R65134 VINN.n264 VINN.n181 4.5005
R65135 VINN.n304 VINN.n181 4.5005
R65136 VINN.n263 VINN.n181 4.5005
R65137 VINN.n306 VINN.n181 4.5005
R65138 VINN.n262 VINN.n181 4.5005
R65139 VINN.n308 VINN.n181 4.5005
R65140 VINN.n261 VINN.n181 4.5005
R65141 VINN.n310 VINN.n181 4.5005
R65142 VINN.n260 VINN.n181 4.5005
R65143 VINN.n312 VINN.n181 4.5005
R65144 VINN.n259 VINN.n181 4.5005
R65145 VINN.n314 VINN.n181 4.5005
R65146 VINN.n258 VINN.n181 4.5005
R65147 VINN.n316 VINN.n181 4.5005
R65148 VINN.n257 VINN.n181 4.5005
R65149 VINN.n318 VINN.n181 4.5005
R65150 VINN.n256 VINN.n181 4.5005
R65151 VINN.n320 VINN.n181 4.5005
R65152 VINN.n255 VINN.n181 4.5005
R65153 VINN.n322 VINN.n181 4.5005
R65154 VINN.n254 VINN.n181 4.5005
R65155 VINN.n324 VINN.n181 4.5005
R65156 VINN.n253 VINN.n181 4.5005
R65157 VINN.n326 VINN.n181 4.5005
R65158 VINN.n252 VINN.n181 4.5005
R65159 VINN.n328 VINN.n181 4.5005
R65160 VINN.n251 VINN.n181 4.5005
R65161 VINN.n330 VINN.n181 4.5005
R65162 VINN.n250 VINN.n181 4.5005
R65163 VINN.n332 VINN.n181 4.5005
R65164 VINN.n249 VINN.n181 4.5005
R65165 VINN.n334 VINN.n181 4.5005
R65166 VINN.n248 VINN.n181 4.5005
R65167 VINN.n336 VINN.n181 4.5005
R65168 VINN.n247 VINN.n181 4.5005
R65169 VINN.n338 VINN.n181 4.5005
R65170 VINN.n246 VINN.n181 4.5005
R65171 VINN.n340 VINN.n181 4.5005
R65172 VINN.n245 VINN.n181 4.5005
R65173 VINN.n342 VINN.n181 4.5005
R65174 VINN.n244 VINN.n181 4.5005
R65175 VINN.n344 VINN.n181 4.5005
R65176 VINN.n243 VINN.n181 4.5005
R65177 VINN.n346 VINN.n181 4.5005
R65178 VINN.n242 VINN.n181 4.5005
R65179 VINN.n348 VINN.n181 4.5005
R65180 VINN.n241 VINN.n181 4.5005
R65181 VINN.n350 VINN.n181 4.5005
R65182 VINN.n240 VINN.n181 4.5005
R65183 VINN.n352 VINN.n181 4.5005
R65184 VINN.n239 VINN.n181 4.5005
R65185 VINN.n354 VINN.n181 4.5005
R65186 VINN.n238 VINN.n181 4.5005
R65187 VINN.n356 VINN.n181 4.5005
R65188 VINN.n237 VINN.n181 4.5005
R65189 VINN.n358 VINN.n181 4.5005
R65190 VINN.n236 VINN.n181 4.5005
R65191 VINN.n360 VINN.n181 4.5005
R65192 VINN.n235 VINN.n181 4.5005
R65193 VINN.n362 VINN.n181 4.5005
R65194 VINN.n234 VINN.n181 4.5005
R65195 VINN.n364 VINN.n181 4.5005
R65196 VINN.n233 VINN.n181 4.5005
R65197 VINN.n366 VINN.n181 4.5005
R65198 VINN.n232 VINN.n181 4.5005
R65199 VINN.n368 VINN.n181 4.5005
R65200 VINN.n231 VINN.n181 4.5005
R65201 VINN.n370 VINN.n181 4.5005
R65202 VINN.n230 VINN.n181 4.5005
R65203 VINN.n372 VINN.n181 4.5005
R65204 VINN.n229 VINN.n181 4.5005
R65205 VINN.n374 VINN.n181 4.5005
R65206 VINN.n228 VINN.n181 4.5005
R65207 VINN.n376 VINN.n181 4.5005
R65208 VINN.n227 VINN.n181 4.5005
R65209 VINN.n378 VINN.n181 4.5005
R65210 VINN.n226 VINN.n181 4.5005
R65211 VINN.n380 VINN.n181 4.5005
R65212 VINN.n225 VINN.n181 4.5005
R65213 VINN.n382 VINN.n181 4.5005
R65214 VINN.n224 VINN.n181 4.5005
R65215 VINN.n384 VINN.n181 4.5005
R65216 VINN.n223 VINN.n181 4.5005
R65217 VINN.n386 VINN.n181 4.5005
R65218 VINN.n222 VINN.n181 4.5005
R65219 VINN.n388 VINN.n181 4.5005
R65220 VINN.n221 VINN.n181 4.5005
R65221 VINN.n390 VINN.n181 4.5005
R65222 VINN.n220 VINN.n181 4.5005
R65223 VINN.n392 VINN.n181 4.5005
R65224 VINN.n219 VINN.n181 4.5005
R65225 VINN.n394 VINN.n181 4.5005
R65226 VINN.n218 VINN.n181 4.5005
R65227 VINN.n396 VINN.n181 4.5005
R65228 VINN.n217 VINN.n181 4.5005
R65229 VINN.n398 VINN.n181 4.5005
R65230 VINN.n216 VINN.n181 4.5005
R65231 VINN.n400 VINN.n181 4.5005
R65232 VINN.n215 VINN.n181 4.5005
R65233 VINN.n654 VINN.n181 4.5005
R65234 VINN.n656 VINN.n181 4.5005
R65235 VINN.n181 VINN.n0 4.5005
R65236 VINN.n278 VINN.n119 4.5005
R65237 VINN.n276 VINN.n119 4.5005
R65238 VINN.n280 VINN.n119 4.5005
R65239 VINN.n275 VINN.n119 4.5005
R65240 VINN.n282 VINN.n119 4.5005
R65241 VINN.n274 VINN.n119 4.5005
R65242 VINN.n284 VINN.n119 4.5005
R65243 VINN.n273 VINN.n119 4.5005
R65244 VINN.n286 VINN.n119 4.5005
R65245 VINN.n272 VINN.n119 4.5005
R65246 VINN.n288 VINN.n119 4.5005
R65247 VINN.n271 VINN.n119 4.5005
R65248 VINN.n290 VINN.n119 4.5005
R65249 VINN.n270 VINN.n119 4.5005
R65250 VINN.n292 VINN.n119 4.5005
R65251 VINN.n269 VINN.n119 4.5005
R65252 VINN.n294 VINN.n119 4.5005
R65253 VINN.n268 VINN.n119 4.5005
R65254 VINN.n296 VINN.n119 4.5005
R65255 VINN.n267 VINN.n119 4.5005
R65256 VINN.n298 VINN.n119 4.5005
R65257 VINN.n266 VINN.n119 4.5005
R65258 VINN.n300 VINN.n119 4.5005
R65259 VINN.n265 VINN.n119 4.5005
R65260 VINN.n302 VINN.n119 4.5005
R65261 VINN.n264 VINN.n119 4.5005
R65262 VINN.n304 VINN.n119 4.5005
R65263 VINN.n263 VINN.n119 4.5005
R65264 VINN.n306 VINN.n119 4.5005
R65265 VINN.n262 VINN.n119 4.5005
R65266 VINN.n308 VINN.n119 4.5005
R65267 VINN.n261 VINN.n119 4.5005
R65268 VINN.n310 VINN.n119 4.5005
R65269 VINN.n260 VINN.n119 4.5005
R65270 VINN.n312 VINN.n119 4.5005
R65271 VINN.n259 VINN.n119 4.5005
R65272 VINN.n314 VINN.n119 4.5005
R65273 VINN.n258 VINN.n119 4.5005
R65274 VINN.n316 VINN.n119 4.5005
R65275 VINN.n257 VINN.n119 4.5005
R65276 VINN.n318 VINN.n119 4.5005
R65277 VINN.n256 VINN.n119 4.5005
R65278 VINN.n320 VINN.n119 4.5005
R65279 VINN.n255 VINN.n119 4.5005
R65280 VINN.n322 VINN.n119 4.5005
R65281 VINN.n254 VINN.n119 4.5005
R65282 VINN.n324 VINN.n119 4.5005
R65283 VINN.n253 VINN.n119 4.5005
R65284 VINN.n326 VINN.n119 4.5005
R65285 VINN.n252 VINN.n119 4.5005
R65286 VINN.n328 VINN.n119 4.5005
R65287 VINN.n251 VINN.n119 4.5005
R65288 VINN.n330 VINN.n119 4.5005
R65289 VINN.n250 VINN.n119 4.5005
R65290 VINN.n332 VINN.n119 4.5005
R65291 VINN.n249 VINN.n119 4.5005
R65292 VINN.n334 VINN.n119 4.5005
R65293 VINN.n248 VINN.n119 4.5005
R65294 VINN.n336 VINN.n119 4.5005
R65295 VINN.n247 VINN.n119 4.5005
R65296 VINN.n338 VINN.n119 4.5005
R65297 VINN.n246 VINN.n119 4.5005
R65298 VINN.n340 VINN.n119 4.5005
R65299 VINN.n245 VINN.n119 4.5005
R65300 VINN.n342 VINN.n119 4.5005
R65301 VINN.n244 VINN.n119 4.5005
R65302 VINN.n344 VINN.n119 4.5005
R65303 VINN.n243 VINN.n119 4.5005
R65304 VINN.n346 VINN.n119 4.5005
R65305 VINN.n242 VINN.n119 4.5005
R65306 VINN.n348 VINN.n119 4.5005
R65307 VINN.n241 VINN.n119 4.5005
R65308 VINN.n350 VINN.n119 4.5005
R65309 VINN.n240 VINN.n119 4.5005
R65310 VINN.n352 VINN.n119 4.5005
R65311 VINN.n239 VINN.n119 4.5005
R65312 VINN.n354 VINN.n119 4.5005
R65313 VINN.n238 VINN.n119 4.5005
R65314 VINN.n356 VINN.n119 4.5005
R65315 VINN.n237 VINN.n119 4.5005
R65316 VINN.n358 VINN.n119 4.5005
R65317 VINN.n236 VINN.n119 4.5005
R65318 VINN.n360 VINN.n119 4.5005
R65319 VINN.n235 VINN.n119 4.5005
R65320 VINN.n362 VINN.n119 4.5005
R65321 VINN.n234 VINN.n119 4.5005
R65322 VINN.n364 VINN.n119 4.5005
R65323 VINN.n233 VINN.n119 4.5005
R65324 VINN.n366 VINN.n119 4.5005
R65325 VINN.n232 VINN.n119 4.5005
R65326 VINN.n368 VINN.n119 4.5005
R65327 VINN.n231 VINN.n119 4.5005
R65328 VINN.n370 VINN.n119 4.5005
R65329 VINN.n230 VINN.n119 4.5005
R65330 VINN.n372 VINN.n119 4.5005
R65331 VINN.n229 VINN.n119 4.5005
R65332 VINN.n374 VINN.n119 4.5005
R65333 VINN.n228 VINN.n119 4.5005
R65334 VINN.n376 VINN.n119 4.5005
R65335 VINN.n227 VINN.n119 4.5005
R65336 VINN.n378 VINN.n119 4.5005
R65337 VINN.n226 VINN.n119 4.5005
R65338 VINN.n380 VINN.n119 4.5005
R65339 VINN.n225 VINN.n119 4.5005
R65340 VINN.n382 VINN.n119 4.5005
R65341 VINN.n224 VINN.n119 4.5005
R65342 VINN.n384 VINN.n119 4.5005
R65343 VINN.n223 VINN.n119 4.5005
R65344 VINN.n386 VINN.n119 4.5005
R65345 VINN.n222 VINN.n119 4.5005
R65346 VINN.n388 VINN.n119 4.5005
R65347 VINN.n221 VINN.n119 4.5005
R65348 VINN.n390 VINN.n119 4.5005
R65349 VINN.n220 VINN.n119 4.5005
R65350 VINN.n392 VINN.n119 4.5005
R65351 VINN.n219 VINN.n119 4.5005
R65352 VINN.n394 VINN.n119 4.5005
R65353 VINN.n218 VINN.n119 4.5005
R65354 VINN.n396 VINN.n119 4.5005
R65355 VINN.n217 VINN.n119 4.5005
R65356 VINN.n398 VINN.n119 4.5005
R65357 VINN.n216 VINN.n119 4.5005
R65358 VINN.n400 VINN.n119 4.5005
R65359 VINN.n215 VINN.n119 4.5005
R65360 VINN.n654 VINN.n119 4.5005
R65361 VINN.n656 VINN.n119 4.5005
R65362 VINN.n119 VINN.n0 4.5005
R65363 VINN.n278 VINN.n182 4.5005
R65364 VINN.n276 VINN.n182 4.5005
R65365 VINN.n280 VINN.n182 4.5005
R65366 VINN.n275 VINN.n182 4.5005
R65367 VINN.n282 VINN.n182 4.5005
R65368 VINN.n274 VINN.n182 4.5005
R65369 VINN.n284 VINN.n182 4.5005
R65370 VINN.n273 VINN.n182 4.5005
R65371 VINN.n286 VINN.n182 4.5005
R65372 VINN.n272 VINN.n182 4.5005
R65373 VINN.n288 VINN.n182 4.5005
R65374 VINN.n271 VINN.n182 4.5005
R65375 VINN.n290 VINN.n182 4.5005
R65376 VINN.n270 VINN.n182 4.5005
R65377 VINN.n292 VINN.n182 4.5005
R65378 VINN.n269 VINN.n182 4.5005
R65379 VINN.n294 VINN.n182 4.5005
R65380 VINN.n268 VINN.n182 4.5005
R65381 VINN.n296 VINN.n182 4.5005
R65382 VINN.n267 VINN.n182 4.5005
R65383 VINN.n298 VINN.n182 4.5005
R65384 VINN.n266 VINN.n182 4.5005
R65385 VINN.n300 VINN.n182 4.5005
R65386 VINN.n265 VINN.n182 4.5005
R65387 VINN.n302 VINN.n182 4.5005
R65388 VINN.n264 VINN.n182 4.5005
R65389 VINN.n304 VINN.n182 4.5005
R65390 VINN.n263 VINN.n182 4.5005
R65391 VINN.n306 VINN.n182 4.5005
R65392 VINN.n262 VINN.n182 4.5005
R65393 VINN.n308 VINN.n182 4.5005
R65394 VINN.n261 VINN.n182 4.5005
R65395 VINN.n310 VINN.n182 4.5005
R65396 VINN.n260 VINN.n182 4.5005
R65397 VINN.n312 VINN.n182 4.5005
R65398 VINN.n259 VINN.n182 4.5005
R65399 VINN.n314 VINN.n182 4.5005
R65400 VINN.n258 VINN.n182 4.5005
R65401 VINN.n316 VINN.n182 4.5005
R65402 VINN.n257 VINN.n182 4.5005
R65403 VINN.n318 VINN.n182 4.5005
R65404 VINN.n256 VINN.n182 4.5005
R65405 VINN.n320 VINN.n182 4.5005
R65406 VINN.n255 VINN.n182 4.5005
R65407 VINN.n322 VINN.n182 4.5005
R65408 VINN.n254 VINN.n182 4.5005
R65409 VINN.n324 VINN.n182 4.5005
R65410 VINN.n253 VINN.n182 4.5005
R65411 VINN.n326 VINN.n182 4.5005
R65412 VINN.n252 VINN.n182 4.5005
R65413 VINN.n328 VINN.n182 4.5005
R65414 VINN.n251 VINN.n182 4.5005
R65415 VINN.n330 VINN.n182 4.5005
R65416 VINN.n250 VINN.n182 4.5005
R65417 VINN.n332 VINN.n182 4.5005
R65418 VINN.n249 VINN.n182 4.5005
R65419 VINN.n334 VINN.n182 4.5005
R65420 VINN.n248 VINN.n182 4.5005
R65421 VINN.n336 VINN.n182 4.5005
R65422 VINN.n247 VINN.n182 4.5005
R65423 VINN.n338 VINN.n182 4.5005
R65424 VINN.n246 VINN.n182 4.5005
R65425 VINN.n340 VINN.n182 4.5005
R65426 VINN.n245 VINN.n182 4.5005
R65427 VINN.n342 VINN.n182 4.5005
R65428 VINN.n244 VINN.n182 4.5005
R65429 VINN.n344 VINN.n182 4.5005
R65430 VINN.n243 VINN.n182 4.5005
R65431 VINN.n346 VINN.n182 4.5005
R65432 VINN.n242 VINN.n182 4.5005
R65433 VINN.n348 VINN.n182 4.5005
R65434 VINN.n241 VINN.n182 4.5005
R65435 VINN.n350 VINN.n182 4.5005
R65436 VINN.n240 VINN.n182 4.5005
R65437 VINN.n352 VINN.n182 4.5005
R65438 VINN.n239 VINN.n182 4.5005
R65439 VINN.n354 VINN.n182 4.5005
R65440 VINN.n238 VINN.n182 4.5005
R65441 VINN.n356 VINN.n182 4.5005
R65442 VINN.n237 VINN.n182 4.5005
R65443 VINN.n358 VINN.n182 4.5005
R65444 VINN.n236 VINN.n182 4.5005
R65445 VINN.n360 VINN.n182 4.5005
R65446 VINN.n235 VINN.n182 4.5005
R65447 VINN.n362 VINN.n182 4.5005
R65448 VINN.n234 VINN.n182 4.5005
R65449 VINN.n364 VINN.n182 4.5005
R65450 VINN.n233 VINN.n182 4.5005
R65451 VINN.n366 VINN.n182 4.5005
R65452 VINN.n232 VINN.n182 4.5005
R65453 VINN.n368 VINN.n182 4.5005
R65454 VINN.n231 VINN.n182 4.5005
R65455 VINN.n370 VINN.n182 4.5005
R65456 VINN.n230 VINN.n182 4.5005
R65457 VINN.n372 VINN.n182 4.5005
R65458 VINN.n229 VINN.n182 4.5005
R65459 VINN.n374 VINN.n182 4.5005
R65460 VINN.n228 VINN.n182 4.5005
R65461 VINN.n376 VINN.n182 4.5005
R65462 VINN.n227 VINN.n182 4.5005
R65463 VINN.n378 VINN.n182 4.5005
R65464 VINN.n226 VINN.n182 4.5005
R65465 VINN.n380 VINN.n182 4.5005
R65466 VINN.n225 VINN.n182 4.5005
R65467 VINN.n382 VINN.n182 4.5005
R65468 VINN.n224 VINN.n182 4.5005
R65469 VINN.n384 VINN.n182 4.5005
R65470 VINN.n223 VINN.n182 4.5005
R65471 VINN.n386 VINN.n182 4.5005
R65472 VINN.n222 VINN.n182 4.5005
R65473 VINN.n388 VINN.n182 4.5005
R65474 VINN.n221 VINN.n182 4.5005
R65475 VINN.n390 VINN.n182 4.5005
R65476 VINN.n220 VINN.n182 4.5005
R65477 VINN.n392 VINN.n182 4.5005
R65478 VINN.n219 VINN.n182 4.5005
R65479 VINN.n394 VINN.n182 4.5005
R65480 VINN.n218 VINN.n182 4.5005
R65481 VINN.n396 VINN.n182 4.5005
R65482 VINN.n217 VINN.n182 4.5005
R65483 VINN.n398 VINN.n182 4.5005
R65484 VINN.n216 VINN.n182 4.5005
R65485 VINN.n400 VINN.n182 4.5005
R65486 VINN.n215 VINN.n182 4.5005
R65487 VINN.n654 VINN.n182 4.5005
R65488 VINN.n656 VINN.n182 4.5005
R65489 VINN.n182 VINN.n0 4.5005
R65490 VINN.n278 VINN.n118 4.5005
R65491 VINN.n276 VINN.n118 4.5005
R65492 VINN.n280 VINN.n118 4.5005
R65493 VINN.n275 VINN.n118 4.5005
R65494 VINN.n282 VINN.n118 4.5005
R65495 VINN.n274 VINN.n118 4.5005
R65496 VINN.n284 VINN.n118 4.5005
R65497 VINN.n273 VINN.n118 4.5005
R65498 VINN.n286 VINN.n118 4.5005
R65499 VINN.n272 VINN.n118 4.5005
R65500 VINN.n288 VINN.n118 4.5005
R65501 VINN.n271 VINN.n118 4.5005
R65502 VINN.n290 VINN.n118 4.5005
R65503 VINN.n270 VINN.n118 4.5005
R65504 VINN.n292 VINN.n118 4.5005
R65505 VINN.n269 VINN.n118 4.5005
R65506 VINN.n294 VINN.n118 4.5005
R65507 VINN.n268 VINN.n118 4.5005
R65508 VINN.n296 VINN.n118 4.5005
R65509 VINN.n267 VINN.n118 4.5005
R65510 VINN.n298 VINN.n118 4.5005
R65511 VINN.n266 VINN.n118 4.5005
R65512 VINN.n300 VINN.n118 4.5005
R65513 VINN.n265 VINN.n118 4.5005
R65514 VINN.n302 VINN.n118 4.5005
R65515 VINN.n264 VINN.n118 4.5005
R65516 VINN.n304 VINN.n118 4.5005
R65517 VINN.n263 VINN.n118 4.5005
R65518 VINN.n306 VINN.n118 4.5005
R65519 VINN.n262 VINN.n118 4.5005
R65520 VINN.n308 VINN.n118 4.5005
R65521 VINN.n261 VINN.n118 4.5005
R65522 VINN.n310 VINN.n118 4.5005
R65523 VINN.n260 VINN.n118 4.5005
R65524 VINN.n312 VINN.n118 4.5005
R65525 VINN.n259 VINN.n118 4.5005
R65526 VINN.n314 VINN.n118 4.5005
R65527 VINN.n258 VINN.n118 4.5005
R65528 VINN.n316 VINN.n118 4.5005
R65529 VINN.n257 VINN.n118 4.5005
R65530 VINN.n318 VINN.n118 4.5005
R65531 VINN.n256 VINN.n118 4.5005
R65532 VINN.n320 VINN.n118 4.5005
R65533 VINN.n255 VINN.n118 4.5005
R65534 VINN.n322 VINN.n118 4.5005
R65535 VINN.n254 VINN.n118 4.5005
R65536 VINN.n324 VINN.n118 4.5005
R65537 VINN.n253 VINN.n118 4.5005
R65538 VINN.n326 VINN.n118 4.5005
R65539 VINN.n252 VINN.n118 4.5005
R65540 VINN.n328 VINN.n118 4.5005
R65541 VINN.n251 VINN.n118 4.5005
R65542 VINN.n330 VINN.n118 4.5005
R65543 VINN.n250 VINN.n118 4.5005
R65544 VINN.n332 VINN.n118 4.5005
R65545 VINN.n249 VINN.n118 4.5005
R65546 VINN.n334 VINN.n118 4.5005
R65547 VINN.n248 VINN.n118 4.5005
R65548 VINN.n336 VINN.n118 4.5005
R65549 VINN.n247 VINN.n118 4.5005
R65550 VINN.n338 VINN.n118 4.5005
R65551 VINN.n246 VINN.n118 4.5005
R65552 VINN.n340 VINN.n118 4.5005
R65553 VINN.n245 VINN.n118 4.5005
R65554 VINN.n342 VINN.n118 4.5005
R65555 VINN.n244 VINN.n118 4.5005
R65556 VINN.n344 VINN.n118 4.5005
R65557 VINN.n243 VINN.n118 4.5005
R65558 VINN.n346 VINN.n118 4.5005
R65559 VINN.n242 VINN.n118 4.5005
R65560 VINN.n348 VINN.n118 4.5005
R65561 VINN.n241 VINN.n118 4.5005
R65562 VINN.n350 VINN.n118 4.5005
R65563 VINN.n240 VINN.n118 4.5005
R65564 VINN.n352 VINN.n118 4.5005
R65565 VINN.n239 VINN.n118 4.5005
R65566 VINN.n354 VINN.n118 4.5005
R65567 VINN.n238 VINN.n118 4.5005
R65568 VINN.n356 VINN.n118 4.5005
R65569 VINN.n237 VINN.n118 4.5005
R65570 VINN.n358 VINN.n118 4.5005
R65571 VINN.n236 VINN.n118 4.5005
R65572 VINN.n360 VINN.n118 4.5005
R65573 VINN.n235 VINN.n118 4.5005
R65574 VINN.n362 VINN.n118 4.5005
R65575 VINN.n234 VINN.n118 4.5005
R65576 VINN.n364 VINN.n118 4.5005
R65577 VINN.n233 VINN.n118 4.5005
R65578 VINN.n366 VINN.n118 4.5005
R65579 VINN.n232 VINN.n118 4.5005
R65580 VINN.n368 VINN.n118 4.5005
R65581 VINN.n231 VINN.n118 4.5005
R65582 VINN.n370 VINN.n118 4.5005
R65583 VINN.n230 VINN.n118 4.5005
R65584 VINN.n372 VINN.n118 4.5005
R65585 VINN.n229 VINN.n118 4.5005
R65586 VINN.n374 VINN.n118 4.5005
R65587 VINN.n228 VINN.n118 4.5005
R65588 VINN.n376 VINN.n118 4.5005
R65589 VINN.n227 VINN.n118 4.5005
R65590 VINN.n378 VINN.n118 4.5005
R65591 VINN.n226 VINN.n118 4.5005
R65592 VINN.n380 VINN.n118 4.5005
R65593 VINN.n225 VINN.n118 4.5005
R65594 VINN.n382 VINN.n118 4.5005
R65595 VINN.n224 VINN.n118 4.5005
R65596 VINN.n384 VINN.n118 4.5005
R65597 VINN.n223 VINN.n118 4.5005
R65598 VINN.n386 VINN.n118 4.5005
R65599 VINN.n222 VINN.n118 4.5005
R65600 VINN.n388 VINN.n118 4.5005
R65601 VINN.n221 VINN.n118 4.5005
R65602 VINN.n390 VINN.n118 4.5005
R65603 VINN.n220 VINN.n118 4.5005
R65604 VINN.n392 VINN.n118 4.5005
R65605 VINN.n219 VINN.n118 4.5005
R65606 VINN.n394 VINN.n118 4.5005
R65607 VINN.n218 VINN.n118 4.5005
R65608 VINN.n396 VINN.n118 4.5005
R65609 VINN.n217 VINN.n118 4.5005
R65610 VINN.n398 VINN.n118 4.5005
R65611 VINN.n216 VINN.n118 4.5005
R65612 VINN.n400 VINN.n118 4.5005
R65613 VINN.n215 VINN.n118 4.5005
R65614 VINN.n654 VINN.n118 4.5005
R65615 VINN.n656 VINN.n118 4.5005
R65616 VINN.n118 VINN.n0 4.5005
R65617 VINN.n278 VINN.n183 4.5005
R65618 VINN.n276 VINN.n183 4.5005
R65619 VINN.n280 VINN.n183 4.5005
R65620 VINN.n275 VINN.n183 4.5005
R65621 VINN.n282 VINN.n183 4.5005
R65622 VINN.n274 VINN.n183 4.5005
R65623 VINN.n284 VINN.n183 4.5005
R65624 VINN.n273 VINN.n183 4.5005
R65625 VINN.n286 VINN.n183 4.5005
R65626 VINN.n272 VINN.n183 4.5005
R65627 VINN.n288 VINN.n183 4.5005
R65628 VINN.n271 VINN.n183 4.5005
R65629 VINN.n290 VINN.n183 4.5005
R65630 VINN.n270 VINN.n183 4.5005
R65631 VINN.n292 VINN.n183 4.5005
R65632 VINN.n269 VINN.n183 4.5005
R65633 VINN.n294 VINN.n183 4.5005
R65634 VINN.n268 VINN.n183 4.5005
R65635 VINN.n296 VINN.n183 4.5005
R65636 VINN.n267 VINN.n183 4.5005
R65637 VINN.n298 VINN.n183 4.5005
R65638 VINN.n266 VINN.n183 4.5005
R65639 VINN.n300 VINN.n183 4.5005
R65640 VINN.n265 VINN.n183 4.5005
R65641 VINN.n302 VINN.n183 4.5005
R65642 VINN.n264 VINN.n183 4.5005
R65643 VINN.n304 VINN.n183 4.5005
R65644 VINN.n263 VINN.n183 4.5005
R65645 VINN.n306 VINN.n183 4.5005
R65646 VINN.n262 VINN.n183 4.5005
R65647 VINN.n308 VINN.n183 4.5005
R65648 VINN.n261 VINN.n183 4.5005
R65649 VINN.n310 VINN.n183 4.5005
R65650 VINN.n260 VINN.n183 4.5005
R65651 VINN.n312 VINN.n183 4.5005
R65652 VINN.n259 VINN.n183 4.5005
R65653 VINN.n314 VINN.n183 4.5005
R65654 VINN.n258 VINN.n183 4.5005
R65655 VINN.n316 VINN.n183 4.5005
R65656 VINN.n257 VINN.n183 4.5005
R65657 VINN.n318 VINN.n183 4.5005
R65658 VINN.n256 VINN.n183 4.5005
R65659 VINN.n320 VINN.n183 4.5005
R65660 VINN.n255 VINN.n183 4.5005
R65661 VINN.n322 VINN.n183 4.5005
R65662 VINN.n254 VINN.n183 4.5005
R65663 VINN.n324 VINN.n183 4.5005
R65664 VINN.n253 VINN.n183 4.5005
R65665 VINN.n326 VINN.n183 4.5005
R65666 VINN.n252 VINN.n183 4.5005
R65667 VINN.n328 VINN.n183 4.5005
R65668 VINN.n251 VINN.n183 4.5005
R65669 VINN.n330 VINN.n183 4.5005
R65670 VINN.n250 VINN.n183 4.5005
R65671 VINN.n332 VINN.n183 4.5005
R65672 VINN.n249 VINN.n183 4.5005
R65673 VINN.n334 VINN.n183 4.5005
R65674 VINN.n248 VINN.n183 4.5005
R65675 VINN.n336 VINN.n183 4.5005
R65676 VINN.n247 VINN.n183 4.5005
R65677 VINN.n338 VINN.n183 4.5005
R65678 VINN.n246 VINN.n183 4.5005
R65679 VINN.n340 VINN.n183 4.5005
R65680 VINN.n245 VINN.n183 4.5005
R65681 VINN.n342 VINN.n183 4.5005
R65682 VINN.n244 VINN.n183 4.5005
R65683 VINN.n344 VINN.n183 4.5005
R65684 VINN.n243 VINN.n183 4.5005
R65685 VINN.n346 VINN.n183 4.5005
R65686 VINN.n242 VINN.n183 4.5005
R65687 VINN.n348 VINN.n183 4.5005
R65688 VINN.n241 VINN.n183 4.5005
R65689 VINN.n350 VINN.n183 4.5005
R65690 VINN.n240 VINN.n183 4.5005
R65691 VINN.n352 VINN.n183 4.5005
R65692 VINN.n239 VINN.n183 4.5005
R65693 VINN.n354 VINN.n183 4.5005
R65694 VINN.n238 VINN.n183 4.5005
R65695 VINN.n356 VINN.n183 4.5005
R65696 VINN.n237 VINN.n183 4.5005
R65697 VINN.n358 VINN.n183 4.5005
R65698 VINN.n236 VINN.n183 4.5005
R65699 VINN.n360 VINN.n183 4.5005
R65700 VINN.n235 VINN.n183 4.5005
R65701 VINN.n362 VINN.n183 4.5005
R65702 VINN.n234 VINN.n183 4.5005
R65703 VINN.n364 VINN.n183 4.5005
R65704 VINN.n233 VINN.n183 4.5005
R65705 VINN.n366 VINN.n183 4.5005
R65706 VINN.n232 VINN.n183 4.5005
R65707 VINN.n368 VINN.n183 4.5005
R65708 VINN.n231 VINN.n183 4.5005
R65709 VINN.n370 VINN.n183 4.5005
R65710 VINN.n230 VINN.n183 4.5005
R65711 VINN.n372 VINN.n183 4.5005
R65712 VINN.n229 VINN.n183 4.5005
R65713 VINN.n374 VINN.n183 4.5005
R65714 VINN.n228 VINN.n183 4.5005
R65715 VINN.n376 VINN.n183 4.5005
R65716 VINN.n227 VINN.n183 4.5005
R65717 VINN.n378 VINN.n183 4.5005
R65718 VINN.n226 VINN.n183 4.5005
R65719 VINN.n380 VINN.n183 4.5005
R65720 VINN.n225 VINN.n183 4.5005
R65721 VINN.n382 VINN.n183 4.5005
R65722 VINN.n224 VINN.n183 4.5005
R65723 VINN.n384 VINN.n183 4.5005
R65724 VINN.n223 VINN.n183 4.5005
R65725 VINN.n386 VINN.n183 4.5005
R65726 VINN.n222 VINN.n183 4.5005
R65727 VINN.n388 VINN.n183 4.5005
R65728 VINN.n221 VINN.n183 4.5005
R65729 VINN.n390 VINN.n183 4.5005
R65730 VINN.n220 VINN.n183 4.5005
R65731 VINN.n392 VINN.n183 4.5005
R65732 VINN.n219 VINN.n183 4.5005
R65733 VINN.n394 VINN.n183 4.5005
R65734 VINN.n218 VINN.n183 4.5005
R65735 VINN.n396 VINN.n183 4.5005
R65736 VINN.n217 VINN.n183 4.5005
R65737 VINN.n398 VINN.n183 4.5005
R65738 VINN.n216 VINN.n183 4.5005
R65739 VINN.n400 VINN.n183 4.5005
R65740 VINN.n215 VINN.n183 4.5005
R65741 VINN.n654 VINN.n183 4.5005
R65742 VINN.n656 VINN.n183 4.5005
R65743 VINN.n183 VINN.n0 4.5005
R65744 VINN.n278 VINN.n117 4.5005
R65745 VINN.n276 VINN.n117 4.5005
R65746 VINN.n280 VINN.n117 4.5005
R65747 VINN.n275 VINN.n117 4.5005
R65748 VINN.n282 VINN.n117 4.5005
R65749 VINN.n274 VINN.n117 4.5005
R65750 VINN.n284 VINN.n117 4.5005
R65751 VINN.n273 VINN.n117 4.5005
R65752 VINN.n286 VINN.n117 4.5005
R65753 VINN.n272 VINN.n117 4.5005
R65754 VINN.n288 VINN.n117 4.5005
R65755 VINN.n271 VINN.n117 4.5005
R65756 VINN.n290 VINN.n117 4.5005
R65757 VINN.n270 VINN.n117 4.5005
R65758 VINN.n292 VINN.n117 4.5005
R65759 VINN.n269 VINN.n117 4.5005
R65760 VINN.n294 VINN.n117 4.5005
R65761 VINN.n268 VINN.n117 4.5005
R65762 VINN.n296 VINN.n117 4.5005
R65763 VINN.n267 VINN.n117 4.5005
R65764 VINN.n298 VINN.n117 4.5005
R65765 VINN.n266 VINN.n117 4.5005
R65766 VINN.n300 VINN.n117 4.5005
R65767 VINN.n265 VINN.n117 4.5005
R65768 VINN.n302 VINN.n117 4.5005
R65769 VINN.n264 VINN.n117 4.5005
R65770 VINN.n304 VINN.n117 4.5005
R65771 VINN.n263 VINN.n117 4.5005
R65772 VINN.n306 VINN.n117 4.5005
R65773 VINN.n262 VINN.n117 4.5005
R65774 VINN.n308 VINN.n117 4.5005
R65775 VINN.n261 VINN.n117 4.5005
R65776 VINN.n310 VINN.n117 4.5005
R65777 VINN.n260 VINN.n117 4.5005
R65778 VINN.n312 VINN.n117 4.5005
R65779 VINN.n259 VINN.n117 4.5005
R65780 VINN.n314 VINN.n117 4.5005
R65781 VINN.n258 VINN.n117 4.5005
R65782 VINN.n316 VINN.n117 4.5005
R65783 VINN.n257 VINN.n117 4.5005
R65784 VINN.n318 VINN.n117 4.5005
R65785 VINN.n256 VINN.n117 4.5005
R65786 VINN.n320 VINN.n117 4.5005
R65787 VINN.n255 VINN.n117 4.5005
R65788 VINN.n322 VINN.n117 4.5005
R65789 VINN.n254 VINN.n117 4.5005
R65790 VINN.n324 VINN.n117 4.5005
R65791 VINN.n253 VINN.n117 4.5005
R65792 VINN.n326 VINN.n117 4.5005
R65793 VINN.n252 VINN.n117 4.5005
R65794 VINN.n328 VINN.n117 4.5005
R65795 VINN.n251 VINN.n117 4.5005
R65796 VINN.n330 VINN.n117 4.5005
R65797 VINN.n250 VINN.n117 4.5005
R65798 VINN.n332 VINN.n117 4.5005
R65799 VINN.n249 VINN.n117 4.5005
R65800 VINN.n334 VINN.n117 4.5005
R65801 VINN.n248 VINN.n117 4.5005
R65802 VINN.n336 VINN.n117 4.5005
R65803 VINN.n247 VINN.n117 4.5005
R65804 VINN.n338 VINN.n117 4.5005
R65805 VINN.n246 VINN.n117 4.5005
R65806 VINN.n340 VINN.n117 4.5005
R65807 VINN.n245 VINN.n117 4.5005
R65808 VINN.n342 VINN.n117 4.5005
R65809 VINN.n244 VINN.n117 4.5005
R65810 VINN.n344 VINN.n117 4.5005
R65811 VINN.n243 VINN.n117 4.5005
R65812 VINN.n346 VINN.n117 4.5005
R65813 VINN.n242 VINN.n117 4.5005
R65814 VINN.n348 VINN.n117 4.5005
R65815 VINN.n241 VINN.n117 4.5005
R65816 VINN.n350 VINN.n117 4.5005
R65817 VINN.n240 VINN.n117 4.5005
R65818 VINN.n352 VINN.n117 4.5005
R65819 VINN.n239 VINN.n117 4.5005
R65820 VINN.n354 VINN.n117 4.5005
R65821 VINN.n238 VINN.n117 4.5005
R65822 VINN.n356 VINN.n117 4.5005
R65823 VINN.n237 VINN.n117 4.5005
R65824 VINN.n358 VINN.n117 4.5005
R65825 VINN.n236 VINN.n117 4.5005
R65826 VINN.n360 VINN.n117 4.5005
R65827 VINN.n235 VINN.n117 4.5005
R65828 VINN.n362 VINN.n117 4.5005
R65829 VINN.n234 VINN.n117 4.5005
R65830 VINN.n364 VINN.n117 4.5005
R65831 VINN.n233 VINN.n117 4.5005
R65832 VINN.n366 VINN.n117 4.5005
R65833 VINN.n232 VINN.n117 4.5005
R65834 VINN.n368 VINN.n117 4.5005
R65835 VINN.n231 VINN.n117 4.5005
R65836 VINN.n370 VINN.n117 4.5005
R65837 VINN.n230 VINN.n117 4.5005
R65838 VINN.n372 VINN.n117 4.5005
R65839 VINN.n229 VINN.n117 4.5005
R65840 VINN.n374 VINN.n117 4.5005
R65841 VINN.n228 VINN.n117 4.5005
R65842 VINN.n376 VINN.n117 4.5005
R65843 VINN.n227 VINN.n117 4.5005
R65844 VINN.n378 VINN.n117 4.5005
R65845 VINN.n226 VINN.n117 4.5005
R65846 VINN.n380 VINN.n117 4.5005
R65847 VINN.n225 VINN.n117 4.5005
R65848 VINN.n382 VINN.n117 4.5005
R65849 VINN.n224 VINN.n117 4.5005
R65850 VINN.n384 VINN.n117 4.5005
R65851 VINN.n223 VINN.n117 4.5005
R65852 VINN.n386 VINN.n117 4.5005
R65853 VINN.n222 VINN.n117 4.5005
R65854 VINN.n388 VINN.n117 4.5005
R65855 VINN.n221 VINN.n117 4.5005
R65856 VINN.n390 VINN.n117 4.5005
R65857 VINN.n220 VINN.n117 4.5005
R65858 VINN.n392 VINN.n117 4.5005
R65859 VINN.n219 VINN.n117 4.5005
R65860 VINN.n394 VINN.n117 4.5005
R65861 VINN.n218 VINN.n117 4.5005
R65862 VINN.n396 VINN.n117 4.5005
R65863 VINN.n217 VINN.n117 4.5005
R65864 VINN.n398 VINN.n117 4.5005
R65865 VINN.n216 VINN.n117 4.5005
R65866 VINN.n400 VINN.n117 4.5005
R65867 VINN.n215 VINN.n117 4.5005
R65868 VINN.n654 VINN.n117 4.5005
R65869 VINN.n656 VINN.n117 4.5005
R65870 VINN.n117 VINN.n0 4.5005
R65871 VINN.n278 VINN.n184 4.5005
R65872 VINN.n276 VINN.n184 4.5005
R65873 VINN.n280 VINN.n184 4.5005
R65874 VINN.n275 VINN.n184 4.5005
R65875 VINN.n282 VINN.n184 4.5005
R65876 VINN.n274 VINN.n184 4.5005
R65877 VINN.n284 VINN.n184 4.5005
R65878 VINN.n273 VINN.n184 4.5005
R65879 VINN.n286 VINN.n184 4.5005
R65880 VINN.n272 VINN.n184 4.5005
R65881 VINN.n288 VINN.n184 4.5005
R65882 VINN.n271 VINN.n184 4.5005
R65883 VINN.n290 VINN.n184 4.5005
R65884 VINN.n270 VINN.n184 4.5005
R65885 VINN.n292 VINN.n184 4.5005
R65886 VINN.n269 VINN.n184 4.5005
R65887 VINN.n294 VINN.n184 4.5005
R65888 VINN.n268 VINN.n184 4.5005
R65889 VINN.n296 VINN.n184 4.5005
R65890 VINN.n267 VINN.n184 4.5005
R65891 VINN.n298 VINN.n184 4.5005
R65892 VINN.n266 VINN.n184 4.5005
R65893 VINN.n300 VINN.n184 4.5005
R65894 VINN.n265 VINN.n184 4.5005
R65895 VINN.n302 VINN.n184 4.5005
R65896 VINN.n264 VINN.n184 4.5005
R65897 VINN.n304 VINN.n184 4.5005
R65898 VINN.n263 VINN.n184 4.5005
R65899 VINN.n306 VINN.n184 4.5005
R65900 VINN.n262 VINN.n184 4.5005
R65901 VINN.n308 VINN.n184 4.5005
R65902 VINN.n261 VINN.n184 4.5005
R65903 VINN.n310 VINN.n184 4.5005
R65904 VINN.n260 VINN.n184 4.5005
R65905 VINN.n312 VINN.n184 4.5005
R65906 VINN.n259 VINN.n184 4.5005
R65907 VINN.n314 VINN.n184 4.5005
R65908 VINN.n258 VINN.n184 4.5005
R65909 VINN.n316 VINN.n184 4.5005
R65910 VINN.n257 VINN.n184 4.5005
R65911 VINN.n318 VINN.n184 4.5005
R65912 VINN.n256 VINN.n184 4.5005
R65913 VINN.n320 VINN.n184 4.5005
R65914 VINN.n255 VINN.n184 4.5005
R65915 VINN.n322 VINN.n184 4.5005
R65916 VINN.n254 VINN.n184 4.5005
R65917 VINN.n324 VINN.n184 4.5005
R65918 VINN.n253 VINN.n184 4.5005
R65919 VINN.n326 VINN.n184 4.5005
R65920 VINN.n252 VINN.n184 4.5005
R65921 VINN.n328 VINN.n184 4.5005
R65922 VINN.n251 VINN.n184 4.5005
R65923 VINN.n330 VINN.n184 4.5005
R65924 VINN.n250 VINN.n184 4.5005
R65925 VINN.n332 VINN.n184 4.5005
R65926 VINN.n249 VINN.n184 4.5005
R65927 VINN.n334 VINN.n184 4.5005
R65928 VINN.n248 VINN.n184 4.5005
R65929 VINN.n336 VINN.n184 4.5005
R65930 VINN.n247 VINN.n184 4.5005
R65931 VINN.n338 VINN.n184 4.5005
R65932 VINN.n246 VINN.n184 4.5005
R65933 VINN.n340 VINN.n184 4.5005
R65934 VINN.n245 VINN.n184 4.5005
R65935 VINN.n342 VINN.n184 4.5005
R65936 VINN.n244 VINN.n184 4.5005
R65937 VINN.n344 VINN.n184 4.5005
R65938 VINN.n243 VINN.n184 4.5005
R65939 VINN.n346 VINN.n184 4.5005
R65940 VINN.n242 VINN.n184 4.5005
R65941 VINN.n348 VINN.n184 4.5005
R65942 VINN.n241 VINN.n184 4.5005
R65943 VINN.n350 VINN.n184 4.5005
R65944 VINN.n240 VINN.n184 4.5005
R65945 VINN.n352 VINN.n184 4.5005
R65946 VINN.n239 VINN.n184 4.5005
R65947 VINN.n354 VINN.n184 4.5005
R65948 VINN.n238 VINN.n184 4.5005
R65949 VINN.n356 VINN.n184 4.5005
R65950 VINN.n237 VINN.n184 4.5005
R65951 VINN.n358 VINN.n184 4.5005
R65952 VINN.n236 VINN.n184 4.5005
R65953 VINN.n360 VINN.n184 4.5005
R65954 VINN.n235 VINN.n184 4.5005
R65955 VINN.n362 VINN.n184 4.5005
R65956 VINN.n234 VINN.n184 4.5005
R65957 VINN.n364 VINN.n184 4.5005
R65958 VINN.n233 VINN.n184 4.5005
R65959 VINN.n366 VINN.n184 4.5005
R65960 VINN.n232 VINN.n184 4.5005
R65961 VINN.n368 VINN.n184 4.5005
R65962 VINN.n231 VINN.n184 4.5005
R65963 VINN.n370 VINN.n184 4.5005
R65964 VINN.n230 VINN.n184 4.5005
R65965 VINN.n372 VINN.n184 4.5005
R65966 VINN.n229 VINN.n184 4.5005
R65967 VINN.n374 VINN.n184 4.5005
R65968 VINN.n228 VINN.n184 4.5005
R65969 VINN.n376 VINN.n184 4.5005
R65970 VINN.n227 VINN.n184 4.5005
R65971 VINN.n378 VINN.n184 4.5005
R65972 VINN.n226 VINN.n184 4.5005
R65973 VINN.n380 VINN.n184 4.5005
R65974 VINN.n225 VINN.n184 4.5005
R65975 VINN.n382 VINN.n184 4.5005
R65976 VINN.n224 VINN.n184 4.5005
R65977 VINN.n384 VINN.n184 4.5005
R65978 VINN.n223 VINN.n184 4.5005
R65979 VINN.n386 VINN.n184 4.5005
R65980 VINN.n222 VINN.n184 4.5005
R65981 VINN.n388 VINN.n184 4.5005
R65982 VINN.n221 VINN.n184 4.5005
R65983 VINN.n390 VINN.n184 4.5005
R65984 VINN.n220 VINN.n184 4.5005
R65985 VINN.n392 VINN.n184 4.5005
R65986 VINN.n219 VINN.n184 4.5005
R65987 VINN.n394 VINN.n184 4.5005
R65988 VINN.n218 VINN.n184 4.5005
R65989 VINN.n396 VINN.n184 4.5005
R65990 VINN.n217 VINN.n184 4.5005
R65991 VINN.n398 VINN.n184 4.5005
R65992 VINN.n216 VINN.n184 4.5005
R65993 VINN.n400 VINN.n184 4.5005
R65994 VINN.n215 VINN.n184 4.5005
R65995 VINN.n654 VINN.n184 4.5005
R65996 VINN.n656 VINN.n184 4.5005
R65997 VINN.n184 VINN.n0 4.5005
R65998 VINN.n278 VINN.n116 4.5005
R65999 VINN.n276 VINN.n116 4.5005
R66000 VINN.n280 VINN.n116 4.5005
R66001 VINN.n275 VINN.n116 4.5005
R66002 VINN.n282 VINN.n116 4.5005
R66003 VINN.n274 VINN.n116 4.5005
R66004 VINN.n284 VINN.n116 4.5005
R66005 VINN.n273 VINN.n116 4.5005
R66006 VINN.n286 VINN.n116 4.5005
R66007 VINN.n272 VINN.n116 4.5005
R66008 VINN.n288 VINN.n116 4.5005
R66009 VINN.n271 VINN.n116 4.5005
R66010 VINN.n290 VINN.n116 4.5005
R66011 VINN.n270 VINN.n116 4.5005
R66012 VINN.n292 VINN.n116 4.5005
R66013 VINN.n269 VINN.n116 4.5005
R66014 VINN.n294 VINN.n116 4.5005
R66015 VINN.n268 VINN.n116 4.5005
R66016 VINN.n296 VINN.n116 4.5005
R66017 VINN.n267 VINN.n116 4.5005
R66018 VINN.n298 VINN.n116 4.5005
R66019 VINN.n266 VINN.n116 4.5005
R66020 VINN.n300 VINN.n116 4.5005
R66021 VINN.n265 VINN.n116 4.5005
R66022 VINN.n302 VINN.n116 4.5005
R66023 VINN.n264 VINN.n116 4.5005
R66024 VINN.n304 VINN.n116 4.5005
R66025 VINN.n263 VINN.n116 4.5005
R66026 VINN.n306 VINN.n116 4.5005
R66027 VINN.n262 VINN.n116 4.5005
R66028 VINN.n308 VINN.n116 4.5005
R66029 VINN.n261 VINN.n116 4.5005
R66030 VINN.n310 VINN.n116 4.5005
R66031 VINN.n260 VINN.n116 4.5005
R66032 VINN.n312 VINN.n116 4.5005
R66033 VINN.n259 VINN.n116 4.5005
R66034 VINN.n314 VINN.n116 4.5005
R66035 VINN.n258 VINN.n116 4.5005
R66036 VINN.n316 VINN.n116 4.5005
R66037 VINN.n257 VINN.n116 4.5005
R66038 VINN.n318 VINN.n116 4.5005
R66039 VINN.n256 VINN.n116 4.5005
R66040 VINN.n320 VINN.n116 4.5005
R66041 VINN.n255 VINN.n116 4.5005
R66042 VINN.n322 VINN.n116 4.5005
R66043 VINN.n254 VINN.n116 4.5005
R66044 VINN.n324 VINN.n116 4.5005
R66045 VINN.n253 VINN.n116 4.5005
R66046 VINN.n326 VINN.n116 4.5005
R66047 VINN.n252 VINN.n116 4.5005
R66048 VINN.n328 VINN.n116 4.5005
R66049 VINN.n251 VINN.n116 4.5005
R66050 VINN.n330 VINN.n116 4.5005
R66051 VINN.n250 VINN.n116 4.5005
R66052 VINN.n332 VINN.n116 4.5005
R66053 VINN.n249 VINN.n116 4.5005
R66054 VINN.n334 VINN.n116 4.5005
R66055 VINN.n248 VINN.n116 4.5005
R66056 VINN.n336 VINN.n116 4.5005
R66057 VINN.n247 VINN.n116 4.5005
R66058 VINN.n338 VINN.n116 4.5005
R66059 VINN.n246 VINN.n116 4.5005
R66060 VINN.n340 VINN.n116 4.5005
R66061 VINN.n245 VINN.n116 4.5005
R66062 VINN.n342 VINN.n116 4.5005
R66063 VINN.n244 VINN.n116 4.5005
R66064 VINN.n344 VINN.n116 4.5005
R66065 VINN.n243 VINN.n116 4.5005
R66066 VINN.n346 VINN.n116 4.5005
R66067 VINN.n242 VINN.n116 4.5005
R66068 VINN.n348 VINN.n116 4.5005
R66069 VINN.n241 VINN.n116 4.5005
R66070 VINN.n350 VINN.n116 4.5005
R66071 VINN.n240 VINN.n116 4.5005
R66072 VINN.n352 VINN.n116 4.5005
R66073 VINN.n239 VINN.n116 4.5005
R66074 VINN.n354 VINN.n116 4.5005
R66075 VINN.n238 VINN.n116 4.5005
R66076 VINN.n356 VINN.n116 4.5005
R66077 VINN.n237 VINN.n116 4.5005
R66078 VINN.n358 VINN.n116 4.5005
R66079 VINN.n236 VINN.n116 4.5005
R66080 VINN.n360 VINN.n116 4.5005
R66081 VINN.n235 VINN.n116 4.5005
R66082 VINN.n362 VINN.n116 4.5005
R66083 VINN.n234 VINN.n116 4.5005
R66084 VINN.n364 VINN.n116 4.5005
R66085 VINN.n233 VINN.n116 4.5005
R66086 VINN.n366 VINN.n116 4.5005
R66087 VINN.n232 VINN.n116 4.5005
R66088 VINN.n368 VINN.n116 4.5005
R66089 VINN.n231 VINN.n116 4.5005
R66090 VINN.n370 VINN.n116 4.5005
R66091 VINN.n230 VINN.n116 4.5005
R66092 VINN.n372 VINN.n116 4.5005
R66093 VINN.n229 VINN.n116 4.5005
R66094 VINN.n374 VINN.n116 4.5005
R66095 VINN.n228 VINN.n116 4.5005
R66096 VINN.n376 VINN.n116 4.5005
R66097 VINN.n227 VINN.n116 4.5005
R66098 VINN.n378 VINN.n116 4.5005
R66099 VINN.n226 VINN.n116 4.5005
R66100 VINN.n380 VINN.n116 4.5005
R66101 VINN.n225 VINN.n116 4.5005
R66102 VINN.n382 VINN.n116 4.5005
R66103 VINN.n224 VINN.n116 4.5005
R66104 VINN.n384 VINN.n116 4.5005
R66105 VINN.n223 VINN.n116 4.5005
R66106 VINN.n386 VINN.n116 4.5005
R66107 VINN.n222 VINN.n116 4.5005
R66108 VINN.n388 VINN.n116 4.5005
R66109 VINN.n221 VINN.n116 4.5005
R66110 VINN.n390 VINN.n116 4.5005
R66111 VINN.n220 VINN.n116 4.5005
R66112 VINN.n392 VINN.n116 4.5005
R66113 VINN.n219 VINN.n116 4.5005
R66114 VINN.n394 VINN.n116 4.5005
R66115 VINN.n218 VINN.n116 4.5005
R66116 VINN.n396 VINN.n116 4.5005
R66117 VINN.n217 VINN.n116 4.5005
R66118 VINN.n398 VINN.n116 4.5005
R66119 VINN.n216 VINN.n116 4.5005
R66120 VINN.n400 VINN.n116 4.5005
R66121 VINN.n215 VINN.n116 4.5005
R66122 VINN.n654 VINN.n116 4.5005
R66123 VINN.n656 VINN.n116 4.5005
R66124 VINN.n116 VINN.n0 4.5005
R66125 VINN.n278 VINN.n185 4.5005
R66126 VINN.n276 VINN.n185 4.5005
R66127 VINN.n280 VINN.n185 4.5005
R66128 VINN.n275 VINN.n185 4.5005
R66129 VINN.n282 VINN.n185 4.5005
R66130 VINN.n274 VINN.n185 4.5005
R66131 VINN.n284 VINN.n185 4.5005
R66132 VINN.n273 VINN.n185 4.5005
R66133 VINN.n286 VINN.n185 4.5005
R66134 VINN.n272 VINN.n185 4.5005
R66135 VINN.n288 VINN.n185 4.5005
R66136 VINN.n271 VINN.n185 4.5005
R66137 VINN.n290 VINN.n185 4.5005
R66138 VINN.n270 VINN.n185 4.5005
R66139 VINN.n292 VINN.n185 4.5005
R66140 VINN.n269 VINN.n185 4.5005
R66141 VINN.n294 VINN.n185 4.5005
R66142 VINN.n268 VINN.n185 4.5005
R66143 VINN.n296 VINN.n185 4.5005
R66144 VINN.n267 VINN.n185 4.5005
R66145 VINN.n298 VINN.n185 4.5005
R66146 VINN.n266 VINN.n185 4.5005
R66147 VINN.n300 VINN.n185 4.5005
R66148 VINN.n265 VINN.n185 4.5005
R66149 VINN.n302 VINN.n185 4.5005
R66150 VINN.n264 VINN.n185 4.5005
R66151 VINN.n304 VINN.n185 4.5005
R66152 VINN.n263 VINN.n185 4.5005
R66153 VINN.n306 VINN.n185 4.5005
R66154 VINN.n262 VINN.n185 4.5005
R66155 VINN.n308 VINN.n185 4.5005
R66156 VINN.n261 VINN.n185 4.5005
R66157 VINN.n310 VINN.n185 4.5005
R66158 VINN.n260 VINN.n185 4.5005
R66159 VINN.n312 VINN.n185 4.5005
R66160 VINN.n259 VINN.n185 4.5005
R66161 VINN.n314 VINN.n185 4.5005
R66162 VINN.n258 VINN.n185 4.5005
R66163 VINN.n316 VINN.n185 4.5005
R66164 VINN.n257 VINN.n185 4.5005
R66165 VINN.n318 VINN.n185 4.5005
R66166 VINN.n256 VINN.n185 4.5005
R66167 VINN.n320 VINN.n185 4.5005
R66168 VINN.n255 VINN.n185 4.5005
R66169 VINN.n322 VINN.n185 4.5005
R66170 VINN.n254 VINN.n185 4.5005
R66171 VINN.n324 VINN.n185 4.5005
R66172 VINN.n253 VINN.n185 4.5005
R66173 VINN.n326 VINN.n185 4.5005
R66174 VINN.n252 VINN.n185 4.5005
R66175 VINN.n328 VINN.n185 4.5005
R66176 VINN.n251 VINN.n185 4.5005
R66177 VINN.n330 VINN.n185 4.5005
R66178 VINN.n250 VINN.n185 4.5005
R66179 VINN.n332 VINN.n185 4.5005
R66180 VINN.n249 VINN.n185 4.5005
R66181 VINN.n334 VINN.n185 4.5005
R66182 VINN.n248 VINN.n185 4.5005
R66183 VINN.n336 VINN.n185 4.5005
R66184 VINN.n247 VINN.n185 4.5005
R66185 VINN.n338 VINN.n185 4.5005
R66186 VINN.n246 VINN.n185 4.5005
R66187 VINN.n340 VINN.n185 4.5005
R66188 VINN.n245 VINN.n185 4.5005
R66189 VINN.n342 VINN.n185 4.5005
R66190 VINN.n244 VINN.n185 4.5005
R66191 VINN.n344 VINN.n185 4.5005
R66192 VINN.n243 VINN.n185 4.5005
R66193 VINN.n346 VINN.n185 4.5005
R66194 VINN.n242 VINN.n185 4.5005
R66195 VINN.n348 VINN.n185 4.5005
R66196 VINN.n241 VINN.n185 4.5005
R66197 VINN.n350 VINN.n185 4.5005
R66198 VINN.n240 VINN.n185 4.5005
R66199 VINN.n352 VINN.n185 4.5005
R66200 VINN.n239 VINN.n185 4.5005
R66201 VINN.n354 VINN.n185 4.5005
R66202 VINN.n238 VINN.n185 4.5005
R66203 VINN.n356 VINN.n185 4.5005
R66204 VINN.n237 VINN.n185 4.5005
R66205 VINN.n358 VINN.n185 4.5005
R66206 VINN.n236 VINN.n185 4.5005
R66207 VINN.n360 VINN.n185 4.5005
R66208 VINN.n235 VINN.n185 4.5005
R66209 VINN.n362 VINN.n185 4.5005
R66210 VINN.n234 VINN.n185 4.5005
R66211 VINN.n364 VINN.n185 4.5005
R66212 VINN.n233 VINN.n185 4.5005
R66213 VINN.n366 VINN.n185 4.5005
R66214 VINN.n232 VINN.n185 4.5005
R66215 VINN.n368 VINN.n185 4.5005
R66216 VINN.n231 VINN.n185 4.5005
R66217 VINN.n370 VINN.n185 4.5005
R66218 VINN.n230 VINN.n185 4.5005
R66219 VINN.n372 VINN.n185 4.5005
R66220 VINN.n229 VINN.n185 4.5005
R66221 VINN.n374 VINN.n185 4.5005
R66222 VINN.n228 VINN.n185 4.5005
R66223 VINN.n376 VINN.n185 4.5005
R66224 VINN.n227 VINN.n185 4.5005
R66225 VINN.n378 VINN.n185 4.5005
R66226 VINN.n226 VINN.n185 4.5005
R66227 VINN.n380 VINN.n185 4.5005
R66228 VINN.n225 VINN.n185 4.5005
R66229 VINN.n382 VINN.n185 4.5005
R66230 VINN.n224 VINN.n185 4.5005
R66231 VINN.n384 VINN.n185 4.5005
R66232 VINN.n223 VINN.n185 4.5005
R66233 VINN.n386 VINN.n185 4.5005
R66234 VINN.n222 VINN.n185 4.5005
R66235 VINN.n388 VINN.n185 4.5005
R66236 VINN.n221 VINN.n185 4.5005
R66237 VINN.n390 VINN.n185 4.5005
R66238 VINN.n220 VINN.n185 4.5005
R66239 VINN.n392 VINN.n185 4.5005
R66240 VINN.n219 VINN.n185 4.5005
R66241 VINN.n394 VINN.n185 4.5005
R66242 VINN.n218 VINN.n185 4.5005
R66243 VINN.n396 VINN.n185 4.5005
R66244 VINN.n217 VINN.n185 4.5005
R66245 VINN.n398 VINN.n185 4.5005
R66246 VINN.n216 VINN.n185 4.5005
R66247 VINN.n400 VINN.n185 4.5005
R66248 VINN.n215 VINN.n185 4.5005
R66249 VINN.n654 VINN.n185 4.5005
R66250 VINN.n656 VINN.n185 4.5005
R66251 VINN.n185 VINN.n0 4.5005
R66252 VINN.n278 VINN.n115 4.5005
R66253 VINN.n276 VINN.n115 4.5005
R66254 VINN.n280 VINN.n115 4.5005
R66255 VINN.n275 VINN.n115 4.5005
R66256 VINN.n282 VINN.n115 4.5005
R66257 VINN.n274 VINN.n115 4.5005
R66258 VINN.n284 VINN.n115 4.5005
R66259 VINN.n273 VINN.n115 4.5005
R66260 VINN.n286 VINN.n115 4.5005
R66261 VINN.n272 VINN.n115 4.5005
R66262 VINN.n288 VINN.n115 4.5005
R66263 VINN.n271 VINN.n115 4.5005
R66264 VINN.n290 VINN.n115 4.5005
R66265 VINN.n270 VINN.n115 4.5005
R66266 VINN.n292 VINN.n115 4.5005
R66267 VINN.n269 VINN.n115 4.5005
R66268 VINN.n294 VINN.n115 4.5005
R66269 VINN.n268 VINN.n115 4.5005
R66270 VINN.n296 VINN.n115 4.5005
R66271 VINN.n267 VINN.n115 4.5005
R66272 VINN.n298 VINN.n115 4.5005
R66273 VINN.n266 VINN.n115 4.5005
R66274 VINN.n300 VINN.n115 4.5005
R66275 VINN.n265 VINN.n115 4.5005
R66276 VINN.n302 VINN.n115 4.5005
R66277 VINN.n264 VINN.n115 4.5005
R66278 VINN.n304 VINN.n115 4.5005
R66279 VINN.n263 VINN.n115 4.5005
R66280 VINN.n306 VINN.n115 4.5005
R66281 VINN.n262 VINN.n115 4.5005
R66282 VINN.n308 VINN.n115 4.5005
R66283 VINN.n261 VINN.n115 4.5005
R66284 VINN.n310 VINN.n115 4.5005
R66285 VINN.n260 VINN.n115 4.5005
R66286 VINN.n312 VINN.n115 4.5005
R66287 VINN.n259 VINN.n115 4.5005
R66288 VINN.n314 VINN.n115 4.5005
R66289 VINN.n258 VINN.n115 4.5005
R66290 VINN.n316 VINN.n115 4.5005
R66291 VINN.n257 VINN.n115 4.5005
R66292 VINN.n318 VINN.n115 4.5005
R66293 VINN.n256 VINN.n115 4.5005
R66294 VINN.n320 VINN.n115 4.5005
R66295 VINN.n255 VINN.n115 4.5005
R66296 VINN.n322 VINN.n115 4.5005
R66297 VINN.n254 VINN.n115 4.5005
R66298 VINN.n324 VINN.n115 4.5005
R66299 VINN.n253 VINN.n115 4.5005
R66300 VINN.n326 VINN.n115 4.5005
R66301 VINN.n252 VINN.n115 4.5005
R66302 VINN.n328 VINN.n115 4.5005
R66303 VINN.n251 VINN.n115 4.5005
R66304 VINN.n330 VINN.n115 4.5005
R66305 VINN.n250 VINN.n115 4.5005
R66306 VINN.n332 VINN.n115 4.5005
R66307 VINN.n249 VINN.n115 4.5005
R66308 VINN.n334 VINN.n115 4.5005
R66309 VINN.n248 VINN.n115 4.5005
R66310 VINN.n336 VINN.n115 4.5005
R66311 VINN.n247 VINN.n115 4.5005
R66312 VINN.n338 VINN.n115 4.5005
R66313 VINN.n246 VINN.n115 4.5005
R66314 VINN.n340 VINN.n115 4.5005
R66315 VINN.n245 VINN.n115 4.5005
R66316 VINN.n342 VINN.n115 4.5005
R66317 VINN.n244 VINN.n115 4.5005
R66318 VINN.n344 VINN.n115 4.5005
R66319 VINN.n243 VINN.n115 4.5005
R66320 VINN.n346 VINN.n115 4.5005
R66321 VINN.n242 VINN.n115 4.5005
R66322 VINN.n348 VINN.n115 4.5005
R66323 VINN.n241 VINN.n115 4.5005
R66324 VINN.n350 VINN.n115 4.5005
R66325 VINN.n240 VINN.n115 4.5005
R66326 VINN.n352 VINN.n115 4.5005
R66327 VINN.n239 VINN.n115 4.5005
R66328 VINN.n354 VINN.n115 4.5005
R66329 VINN.n238 VINN.n115 4.5005
R66330 VINN.n356 VINN.n115 4.5005
R66331 VINN.n237 VINN.n115 4.5005
R66332 VINN.n358 VINN.n115 4.5005
R66333 VINN.n236 VINN.n115 4.5005
R66334 VINN.n360 VINN.n115 4.5005
R66335 VINN.n235 VINN.n115 4.5005
R66336 VINN.n362 VINN.n115 4.5005
R66337 VINN.n234 VINN.n115 4.5005
R66338 VINN.n364 VINN.n115 4.5005
R66339 VINN.n233 VINN.n115 4.5005
R66340 VINN.n366 VINN.n115 4.5005
R66341 VINN.n232 VINN.n115 4.5005
R66342 VINN.n368 VINN.n115 4.5005
R66343 VINN.n231 VINN.n115 4.5005
R66344 VINN.n370 VINN.n115 4.5005
R66345 VINN.n230 VINN.n115 4.5005
R66346 VINN.n372 VINN.n115 4.5005
R66347 VINN.n229 VINN.n115 4.5005
R66348 VINN.n374 VINN.n115 4.5005
R66349 VINN.n228 VINN.n115 4.5005
R66350 VINN.n376 VINN.n115 4.5005
R66351 VINN.n227 VINN.n115 4.5005
R66352 VINN.n378 VINN.n115 4.5005
R66353 VINN.n226 VINN.n115 4.5005
R66354 VINN.n380 VINN.n115 4.5005
R66355 VINN.n225 VINN.n115 4.5005
R66356 VINN.n382 VINN.n115 4.5005
R66357 VINN.n224 VINN.n115 4.5005
R66358 VINN.n384 VINN.n115 4.5005
R66359 VINN.n223 VINN.n115 4.5005
R66360 VINN.n386 VINN.n115 4.5005
R66361 VINN.n222 VINN.n115 4.5005
R66362 VINN.n388 VINN.n115 4.5005
R66363 VINN.n221 VINN.n115 4.5005
R66364 VINN.n390 VINN.n115 4.5005
R66365 VINN.n220 VINN.n115 4.5005
R66366 VINN.n392 VINN.n115 4.5005
R66367 VINN.n219 VINN.n115 4.5005
R66368 VINN.n394 VINN.n115 4.5005
R66369 VINN.n218 VINN.n115 4.5005
R66370 VINN.n396 VINN.n115 4.5005
R66371 VINN.n217 VINN.n115 4.5005
R66372 VINN.n398 VINN.n115 4.5005
R66373 VINN.n216 VINN.n115 4.5005
R66374 VINN.n400 VINN.n115 4.5005
R66375 VINN.n215 VINN.n115 4.5005
R66376 VINN.n654 VINN.n115 4.5005
R66377 VINN.n656 VINN.n115 4.5005
R66378 VINN.n115 VINN.n0 4.5005
R66379 VINN.n278 VINN.n186 4.5005
R66380 VINN.n276 VINN.n186 4.5005
R66381 VINN.n280 VINN.n186 4.5005
R66382 VINN.n275 VINN.n186 4.5005
R66383 VINN.n282 VINN.n186 4.5005
R66384 VINN.n274 VINN.n186 4.5005
R66385 VINN.n284 VINN.n186 4.5005
R66386 VINN.n273 VINN.n186 4.5005
R66387 VINN.n286 VINN.n186 4.5005
R66388 VINN.n272 VINN.n186 4.5005
R66389 VINN.n288 VINN.n186 4.5005
R66390 VINN.n271 VINN.n186 4.5005
R66391 VINN.n290 VINN.n186 4.5005
R66392 VINN.n270 VINN.n186 4.5005
R66393 VINN.n292 VINN.n186 4.5005
R66394 VINN.n269 VINN.n186 4.5005
R66395 VINN.n294 VINN.n186 4.5005
R66396 VINN.n268 VINN.n186 4.5005
R66397 VINN.n296 VINN.n186 4.5005
R66398 VINN.n267 VINN.n186 4.5005
R66399 VINN.n298 VINN.n186 4.5005
R66400 VINN.n266 VINN.n186 4.5005
R66401 VINN.n300 VINN.n186 4.5005
R66402 VINN.n265 VINN.n186 4.5005
R66403 VINN.n302 VINN.n186 4.5005
R66404 VINN.n264 VINN.n186 4.5005
R66405 VINN.n304 VINN.n186 4.5005
R66406 VINN.n263 VINN.n186 4.5005
R66407 VINN.n306 VINN.n186 4.5005
R66408 VINN.n262 VINN.n186 4.5005
R66409 VINN.n308 VINN.n186 4.5005
R66410 VINN.n261 VINN.n186 4.5005
R66411 VINN.n310 VINN.n186 4.5005
R66412 VINN.n260 VINN.n186 4.5005
R66413 VINN.n312 VINN.n186 4.5005
R66414 VINN.n259 VINN.n186 4.5005
R66415 VINN.n314 VINN.n186 4.5005
R66416 VINN.n258 VINN.n186 4.5005
R66417 VINN.n316 VINN.n186 4.5005
R66418 VINN.n257 VINN.n186 4.5005
R66419 VINN.n318 VINN.n186 4.5005
R66420 VINN.n256 VINN.n186 4.5005
R66421 VINN.n320 VINN.n186 4.5005
R66422 VINN.n255 VINN.n186 4.5005
R66423 VINN.n322 VINN.n186 4.5005
R66424 VINN.n254 VINN.n186 4.5005
R66425 VINN.n324 VINN.n186 4.5005
R66426 VINN.n253 VINN.n186 4.5005
R66427 VINN.n326 VINN.n186 4.5005
R66428 VINN.n252 VINN.n186 4.5005
R66429 VINN.n328 VINN.n186 4.5005
R66430 VINN.n251 VINN.n186 4.5005
R66431 VINN.n330 VINN.n186 4.5005
R66432 VINN.n250 VINN.n186 4.5005
R66433 VINN.n332 VINN.n186 4.5005
R66434 VINN.n249 VINN.n186 4.5005
R66435 VINN.n334 VINN.n186 4.5005
R66436 VINN.n248 VINN.n186 4.5005
R66437 VINN.n336 VINN.n186 4.5005
R66438 VINN.n247 VINN.n186 4.5005
R66439 VINN.n338 VINN.n186 4.5005
R66440 VINN.n246 VINN.n186 4.5005
R66441 VINN.n340 VINN.n186 4.5005
R66442 VINN.n245 VINN.n186 4.5005
R66443 VINN.n342 VINN.n186 4.5005
R66444 VINN.n244 VINN.n186 4.5005
R66445 VINN.n344 VINN.n186 4.5005
R66446 VINN.n243 VINN.n186 4.5005
R66447 VINN.n346 VINN.n186 4.5005
R66448 VINN.n242 VINN.n186 4.5005
R66449 VINN.n348 VINN.n186 4.5005
R66450 VINN.n241 VINN.n186 4.5005
R66451 VINN.n350 VINN.n186 4.5005
R66452 VINN.n240 VINN.n186 4.5005
R66453 VINN.n352 VINN.n186 4.5005
R66454 VINN.n239 VINN.n186 4.5005
R66455 VINN.n354 VINN.n186 4.5005
R66456 VINN.n238 VINN.n186 4.5005
R66457 VINN.n356 VINN.n186 4.5005
R66458 VINN.n237 VINN.n186 4.5005
R66459 VINN.n358 VINN.n186 4.5005
R66460 VINN.n236 VINN.n186 4.5005
R66461 VINN.n360 VINN.n186 4.5005
R66462 VINN.n235 VINN.n186 4.5005
R66463 VINN.n362 VINN.n186 4.5005
R66464 VINN.n234 VINN.n186 4.5005
R66465 VINN.n364 VINN.n186 4.5005
R66466 VINN.n233 VINN.n186 4.5005
R66467 VINN.n366 VINN.n186 4.5005
R66468 VINN.n232 VINN.n186 4.5005
R66469 VINN.n368 VINN.n186 4.5005
R66470 VINN.n231 VINN.n186 4.5005
R66471 VINN.n370 VINN.n186 4.5005
R66472 VINN.n230 VINN.n186 4.5005
R66473 VINN.n372 VINN.n186 4.5005
R66474 VINN.n229 VINN.n186 4.5005
R66475 VINN.n374 VINN.n186 4.5005
R66476 VINN.n228 VINN.n186 4.5005
R66477 VINN.n376 VINN.n186 4.5005
R66478 VINN.n227 VINN.n186 4.5005
R66479 VINN.n378 VINN.n186 4.5005
R66480 VINN.n226 VINN.n186 4.5005
R66481 VINN.n380 VINN.n186 4.5005
R66482 VINN.n225 VINN.n186 4.5005
R66483 VINN.n382 VINN.n186 4.5005
R66484 VINN.n224 VINN.n186 4.5005
R66485 VINN.n384 VINN.n186 4.5005
R66486 VINN.n223 VINN.n186 4.5005
R66487 VINN.n386 VINN.n186 4.5005
R66488 VINN.n222 VINN.n186 4.5005
R66489 VINN.n388 VINN.n186 4.5005
R66490 VINN.n221 VINN.n186 4.5005
R66491 VINN.n390 VINN.n186 4.5005
R66492 VINN.n220 VINN.n186 4.5005
R66493 VINN.n392 VINN.n186 4.5005
R66494 VINN.n219 VINN.n186 4.5005
R66495 VINN.n394 VINN.n186 4.5005
R66496 VINN.n218 VINN.n186 4.5005
R66497 VINN.n396 VINN.n186 4.5005
R66498 VINN.n217 VINN.n186 4.5005
R66499 VINN.n398 VINN.n186 4.5005
R66500 VINN.n216 VINN.n186 4.5005
R66501 VINN.n400 VINN.n186 4.5005
R66502 VINN.n215 VINN.n186 4.5005
R66503 VINN.n654 VINN.n186 4.5005
R66504 VINN.n656 VINN.n186 4.5005
R66505 VINN.n186 VINN.n0 4.5005
R66506 VINN.n278 VINN.n114 4.5005
R66507 VINN.n276 VINN.n114 4.5005
R66508 VINN.n280 VINN.n114 4.5005
R66509 VINN.n275 VINN.n114 4.5005
R66510 VINN.n282 VINN.n114 4.5005
R66511 VINN.n274 VINN.n114 4.5005
R66512 VINN.n284 VINN.n114 4.5005
R66513 VINN.n273 VINN.n114 4.5005
R66514 VINN.n286 VINN.n114 4.5005
R66515 VINN.n272 VINN.n114 4.5005
R66516 VINN.n288 VINN.n114 4.5005
R66517 VINN.n271 VINN.n114 4.5005
R66518 VINN.n290 VINN.n114 4.5005
R66519 VINN.n270 VINN.n114 4.5005
R66520 VINN.n292 VINN.n114 4.5005
R66521 VINN.n269 VINN.n114 4.5005
R66522 VINN.n294 VINN.n114 4.5005
R66523 VINN.n268 VINN.n114 4.5005
R66524 VINN.n296 VINN.n114 4.5005
R66525 VINN.n267 VINN.n114 4.5005
R66526 VINN.n298 VINN.n114 4.5005
R66527 VINN.n266 VINN.n114 4.5005
R66528 VINN.n300 VINN.n114 4.5005
R66529 VINN.n265 VINN.n114 4.5005
R66530 VINN.n302 VINN.n114 4.5005
R66531 VINN.n264 VINN.n114 4.5005
R66532 VINN.n304 VINN.n114 4.5005
R66533 VINN.n263 VINN.n114 4.5005
R66534 VINN.n306 VINN.n114 4.5005
R66535 VINN.n262 VINN.n114 4.5005
R66536 VINN.n308 VINN.n114 4.5005
R66537 VINN.n261 VINN.n114 4.5005
R66538 VINN.n310 VINN.n114 4.5005
R66539 VINN.n260 VINN.n114 4.5005
R66540 VINN.n312 VINN.n114 4.5005
R66541 VINN.n259 VINN.n114 4.5005
R66542 VINN.n314 VINN.n114 4.5005
R66543 VINN.n258 VINN.n114 4.5005
R66544 VINN.n316 VINN.n114 4.5005
R66545 VINN.n257 VINN.n114 4.5005
R66546 VINN.n318 VINN.n114 4.5005
R66547 VINN.n256 VINN.n114 4.5005
R66548 VINN.n320 VINN.n114 4.5005
R66549 VINN.n255 VINN.n114 4.5005
R66550 VINN.n322 VINN.n114 4.5005
R66551 VINN.n254 VINN.n114 4.5005
R66552 VINN.n324 VINN.n114 4.5005
R66553 VINN.n253 VINN.n114 4.5005
R66554 VINN.n326 VINN.n114 4.5005
R66555 VINN.n252 VINN.n114 4.5005
R66556 VINN.n328 VINN.n114 4.5005
R66557 VINN.n251 VINN.n114 4.5005
R66558 VINN.n330 VINN.n114 4.5005
R66559 VINN.n250 VINN.n114 4.5005
R66560 VINN.n332 VINN.n114 4.5005
R66561 VINN.n249 VINN.n114 4.5005
R66562 VINN.n334 VINN.n114 4.5005
R66563 VINN.n248 VINN.n114 4.5005
R66564 VINN.n336 VINN.n114 4.5005
R66565 VINN.n247 VINN.n114 4.5005
R66566 VINN.n338 VINN.n114 4.5005
R66567 VINN.n246 VINN.n114 4.5005
R66568 VINN.n340 VINN.n114 4.5005
R66569 VINN.n245 VINN.n114 4.5005
R66570 VINN.n342 VINN.n114 4.5005
R66571 VINN.n244 VINN.n114 4.5005
R66572 VINN.n344 VINN.n114 4.5005
R66573 VINN.n243 VINN.n114 4.5005
R66574 VINN.n346 VINN.n114 4.5005
R66575 VINN.n242 VINN.n114 4.5005
R66576 VINN.n348 VINN.n114 4.5005
R66577 VINN.n241 VINN.n114 4.5005
R66578 VINN.n350 VINN.n114 4.5005
R66579 VINN.n240 VINN.n114 4.5005
R66580 VINN.n352 VINN.n114 4.5005
R66581 VINN.n239 VINN.n114 4.5005
R66582 VINN.n354 VINN.n114 4.5005
R66583 VINN.n238 VINN.n114 4.5005
R66584 VINN.n356 VINN.n114 4.5005
R66585 VINN.n237 VINN.n114 4.5005
R66586 VINN.n358 VINN.n114 4.5005
R66587 VINN.n236 VINN.n114 4.5005
R66588 VINN.n360 VINN.n114 4.5005
R66589 VINN.n235 VINN.n114 4.5005
R66590 VINN.n362 VINN.n114 4.5005
R66591 VINN.n234 VINN.n114 4.5005
R66592 VINN.n364 VINN.n114 4.5005
R66593 VINN.n233 VINN.n114 4.5005
R66594 VINN.n366 VINN.n114 4.5005
R66595 VINN.n232 VINN.n114 4.5005
R66596 VINN.n368 VINN.n114 4.5005
R66597 VINN.n231 VINN.n114 4.5005
R66598 VINN.n370 VINN.n114 4.5005
R66599 VINN.n230 VINN.n114 4.5005
R66600 VINN.n372 VINN.n114 4.5005
R66601 VINN.n229 VINN.n114 4.5005
R66602 VINN.n374 VINN.n114 4.5005
R66603 VINN.n228 VINN.n114 4.5005
R66604 VINN.n376 VINN.n114 4.5005
R66605 VINN.n227 VINN.n114 4.5005
R66606 VINN.n378 VINN.n114 4.5005
R66607 VINN.n226 VINN.n114 4.5005
R66608 VINN.n380 VINN.n114 4.5005
R66609 VINN.n225 VINN.n114 4.5005
R66610 VINN.n382 VINN.n114 4.5005
R66611 VINN.n224 VINN.n114 4.5005
R66612 VINN.n384 VINN.n114 4.5005
R66613 VINN.n223 VINN.n114 4.5005
R66614 VINN.n386 VINN.n114 4.5005
R66615 VINN.n222 VINN.n114 4.5005
R66616 VINN.n388 VINN.n114 4.5005
R66617 VINN.n221 VINN.n114 4.5005
R66618 VINN.n390 VINN.n114 4.5005
R66619 VINN.n220 VINN.n114 4.5005
R66620 VINN.n392 VINN.n114 4.5005
R66621 VINN.n219 VINN.n114 4.5005
R66622 VINN.n394 VINN.n114 4.5005
R66623 VINN.n218 VINN.n114 4.5005
R66624 VINN.n396 VINN.n114 4.5005
R66625 VINN.n217 VINN.n114 4.5005
R66626 VINN.n398 VINN.n114 4.5005
R66627 VINN.n216 VINN.n114 4.5005
R66628 VINN.n400 VINN.n114 4.5005
R66629 VINN.n215 VINN.n114 4.5005
R66630 VINN.n654 VINN.n114 4.5005
R66631 VINN.n656 VINN.n114 4.5005
R66632 VINN.n114 VINN.n0 4.5005
R66633 VINN.n278 VINN.n187 4.5005
R66634 VINN.n276 VINN.n187 4.5005
R66635 VINN.n280 VINN.n187 4.5005
R66636 VINN.n275 VINN.n187 4.5005
R66637 VINN.n282 VINN.n187 4.5005
R66638 VINN.n274 VINN.n187 4.5005
R66639 VINN.n284 VINN.n187 4.5005
R66640 VINN.n273 VINN.n187 4.5005
R66641 VINN.n286 VINN.n187 4.5005
R66642 VINN.n272 VINN.n187 4.5005
R66643 VINN.n288 VINN.n187 4.5005
R66644 VINN.n271 VINN.n187 4.5005
R66645 VINN.n290 VINN.n187 4.5005
R66646 VINN.n270 VINN.n187 4.5005
R66647 VINN.n292 VINN.n187 4.5005
R66648 VINN.n269 VINN.n187 4.5005
R66649 VINN.n294 VINN.n187 4.5005
R66650 VINN.n268 VINN.n187 4.5005
R66651 VINN.n296 VINN.n187 4.5005
R66652 VINN.n267 VINN.n187 4.5005
R66653 VINN.n298 VINN.n187 4.5005
R66654 VINN.n266 VINN.n187 4.5005
R66655 VINN.n300 VINN.n187 4.5005
R66656 VINN.n265 VINN.n187 4.5005
R66657 VINN.n302 VINN.n187 4.5005
R66658 VINN.n264 VINN.n187 4.5005
R66659 VINN.n304 VINN.n187 4.5005
R66660 VINN.n263 VINN.n187 4.5005
R66661 VINN.n306 VINN.n187 4.5005
R66662 VINN.n262 VINN.n187 4.5005
R66663 VINN.n308 VINN.n187 4.5005
R66664 VINN.n261 VINN.n187 4.5005
R66665 VINN.n310 VINN.n187 4.5005
R66666 VINN.n260 VINN.n187 4.5005
R66667 VINN.n312 VINN.n187 4.5005
R66668 VINN.n259 VINN.n187 4.5005
R66669 VINN.n314 VINN.n187 4.5005
R66670 VINN.n258 VINN.n187 4.5005
R66671 VINN.n316 VINN.n187 4.5005
R66672 VINN.n257 VINN.n187 4.5005
R66673 VINN.n318 VINN.n187 4.5005
R66674 VINN.n256 VINN.n187 4.5005
R66675 VINN.n320 VINN.n187 4.5005
R66676 VINN.n255 VINN.n187 4.5005
R66677 VINN.n322 VINN.n187 4.5005
R66678 VINN.n254 VINN.n187 4.5005
R66679 VINN.n324 VINN.n187 4.5005
R66680 VINN.n253 VINN.n187 4.5005
R66681 VINN.n326 VINN.n187 4.5005
R66682 VINN.n252 VINN.n187 4.5005
R66683 VINN.n328 VINN.n187 4.5005
R66684 VINN.n251 VINN.n187 4.5005
R66685 VINN.n330 VINN.n187 4.5005
R66686 VINN.n250 VINN.n187 4.5005
R66687 VINN.n332 VINN.n187 4.5005
R66688 VINN.n249 VINN.n187 4.5005
R66689 VINN.n334 VINN.n187 4.5005
R66690 VINN.n248 VINN.n187 4.5005
R66691 VINN.n336 VINN.n187 4.5005
R66692 VINN.n247 VINN.n187 4.5005
R66693 VINN.n338 VINN.n187 4.5005
R66694 VINN.n246 VINN.n187 4.5005
R66695 VINN.n340 VINN.n187 4.5005
R66696 VINN.n245 VINN.n187 4.5005
R66697 VINN.n342 VINN.n187 4.5005
R66698 VINN.n244 VINN.n187 4.5005
R66699 VINN.n344 VINN.n187 4.5005
R66700 VINN.n243 VINN.n187 4.5005
R66701 VINN.n346 VINN.n187 4.5005
R66702 VINN.n242 VINN.n187 4.5005
R66703 VINN.n348 VINN.n187 4.5005
R66704 VINN.n241 VINN.n187 4.5005
R66705 VINN.n350 VINN.n187 4.5005
R66706 VINN.n240 VINN.n187 4.5005
R66707 VINN.n352 VINN.n187 4.5005
R66708 VINN.n239 VINN.n187 4.5005
R66709 VINN.n354 VINN.n187 4.5005
R66710 VINN.n238 VINN.n187 4.5005
R66711 VINN.n356 VINN.n187 4.5005
R66712 VINN.n237 VINN.n187 4.5005
R66713 VINN.n358 VINN.n187 4.5005
R66714 VINN.n236 VINN.n187 4.5005
R66715 VINN.n360 VINN.n187 4.5005
R66716 VINN.n235 VINN.n187 4.5005
R66717 VINN.n362 VINN.n187 4.5005
R66718 VINN.n234 VINN.n187 4.5005
R66719 VINN.n364 VINN.n187 4.5005
R66720 VINN.n233 VINN.n187 4.5005
R66721 VINN.n366 VINN.n187 4.5005
R66722 VINN.n232 VINN.n187 4.5005
R66723 VINN.n368 VINN.n187 4.5005
R66724 VINN.n231 VINN.n187 4.5005
R66725 VINN.n370 VINN.n187 4.5005
R66726 VINN.n230 VINN.n187 4.5005
R66727 VINN.n372 VINN.n187 4.5005
R66728 VINN.n229 VINN.n187 4.5005
R66729 VINN.n374 VINN.n187 4.5005
R66730 VINN.n228 VINN.n187 4.5005
R66731 VINN.n376 VINN.n187 4.5005
R66732 VINN.n227 VINN.n187 4.5005
R66733 VINN.n378 VINN.n187 4.5005
R66734 VINN.n226 VINN.n187 4.5005
R66735 VINN.n380 VINN.n187 4.5005
R66736 VINN.n225 VINN.n187 4.5005
R66737 VINN.n382 VINN.n187 4.5005
R66738 VINN.n224 VINN.n187 4.5005
R66739 VINN.n384 VINN.n187 4.5005
R66740 VINN.n223 VINN.n187 4.5005
R66741 VINN.n386 VINN.n187 4.5005
R66742 VINN.n222 VINN.n187 4.5005
R66743 VINN.n388 VINN.n187 4.5005
R66744 VINN.n221 VINN.n187 4.5005
R66745 VINN.n390 VINN.n187 4.5005
R66746 VINN.n220 VINN.n187 4.5005
R66747 VINN.n392 VINN.n187 4.5005
R66748 VINN.n219 VINN.n187 4.5005
R66749 VINN.n394 VINN.n187 4.5005
R66750 VINN.n218 VINN.n187 4.5005
R66751 VINN.n396 VINN.n187 4.5005
R66752 VINN.n217 VINN.n187 4.5005
R66753 VINN.n398 VINN.n187 4.5005
R66754 VINN.n216 VINN.n187 4.5005
R66755 VINN.n400 VINN.n187 4.5005
R66756 VINN.n215 VINN.n187 4.5005
R66757 VINN.n654 VINN.n187 4.5005
R66758 VINN.n656 VINN.n187 4.5005
R66759 VINN.n187 VINN.n0 4.5005
R66760 VINN.n278 VINN.n113 4.5005
R66761 VINN.n276 VINN.n113 4.5005
R66762 VINN.n280 VINN.n113 4.5005
R66763 VINN.n275 VINN.n113 4.5005
R66764 VINN.n282 VINN.n113 4.5005
R66765 VINN.n274 VINN.n113 4.5005
R66766 VINN.n284 VINN.n113 4.5005
R66767 VINN.n273 VINN.n113 4.5005
R66768 VINN.n286 VINN.n113 4.5005
R66769 VINN.n272 VINN.n113 4.5005
R66770 VINN.n288 VINN.n113 4.5005
R66771 VINN.n271 VINN.n113 4.5005
R66772 VINN.n290 VINN.n113 4.5005
R66773 VINN.n270 VINN.n113 4.5005
R66774 VINN.n292 VINN.n113 4.5005
R66775 VINN.n269 VINN.n113 4.5005
R66776 VINN.n294 VINN.n113 4.5005
R66777 VINN.n268 VINN.n113 4.5005
R66778 VINN.n296 VINN.n113 4.5005
R66779 VINN.n267 VINN.n113 4.5005
R66780 VINN.n298 VINN.n113 4.5005
R66781 VINN.n266 VINN.n113 4.5005
R66782 VINN.n300 VINN.n113 4.5005
R66783 VINN.n265 VINN.n113 4.5005
R66784 VINN.n302 VINN.n113 4.5005
R66785 VINN.n264 VINN.n113 4.5005
R66786 VINN.n304 VINN.n113 4.5005
R66787 VINN.n263 VINN.n113 4.5005
R66788 VINN.n306 VINN.n113 4.5005
R66789 VINN.n262 VINN.n113 4.5005
R66790 VINN.n308 VINN.n113 4.5005
R66791 VINN.n261 VINN.n113 4.5005
R66792 VINN.n310 VINN.n113 4.5005
R66793 VINN.n260 VINN.n113 4.5005
R66794 VINN.n312 VINN.n113 4.5005
R66795 VINN.n259 VINN.n113 4.5005
R66796 VINN.n314 VINN.n113 4.5005
R66797 VINN.n258 VINN.n113 4.5005
R66798 VINN.n316 VINN.n113 4.5005
R66799 VINN.n257 VINN.n113 4.5005
R66800 VINN.n318 VINN.n113 4.5005
R66801 VINN.n256 VINN.n113 4.5005
R66802 VINN.n320 VINN.n113 4.5005
R66803 VINN.n255 VINN.n113 4.5005
R66804 VINN.n322 VINN.n113 4.5005
R66805 VINN.n254 VINN.n113 4.5005
R66806 VINN.n324 VINN.n113 4.5005
R66807 VINN.n253 VINN.n113 4.5005
R66808 VINN.n326 VINN.n113 4.5005
R66809 VINN.n252 VINN.n113 4.5005
R66810 VINN.n328 VINN.n113 4.5005
R66811 VINN.n251 VINN.n113 4.5005
R66812 VINN.n330 VINN.n113 4.5005
R66813 VINN.n250 VINN.n113 4.5005
R66814 VINN.n332 VINN.n113 4.5005
R66815 VINN.n249 VINN.n113 4.5005
R66816 VINN.n334 VINN.n113 4.5005
R66817 VINN.n248 VINN.n113 4.5005
R66818 VINN.n336 VINN.n113 4.5005
R66819 VINN.n247 VINN.n113 4.5005
R66820 VINN.n338 VINN.n113 4.5005
R66821 VINN.n246 VINN.n113 4.5005
R66822 VINN.n340 VINN.n113 4.5005
R66823 VINN.n245 VINN.n113 4.5005
R66824 VINN.n342 VINN.n113 4.5005
R66825 VINN.n244 VINN.n113 4.5005
R66826 VINN.n344 VINN.n113 4.5005
R66827 VINN.n243 VINN.n113 4.5005
R66828 VINN.n346 VINN.n113 4.5005
R66829 VINN.n242 VINN.n113 4.5005
R66830 VINN.n348 VINN.n113 4.5005
R66831 VINN.n241 VINN.n113 4.5005
R66832 VINN.n350 VINN.n113 4.5005
R66833 VINN.n240 VINN.n113 4.5005
R66834 VINN.n352 VINN.n113 4.5005
R66835 VINN.n239 VINN.n113 4.5005
R66836 VINN.n354 VINN.n113 4.5005
R66837 VINN.n238 VINN.n113 4.5005
R66838 VINN.n356 VINN.n113 4.5005
R66839 VINN.n237 VINN.n113 4.5005
R66840 VINN.n358 VINN.n113 4.5005
R66841 VINN.n236 VINN.n113 4.5005
R66842 VINN.n360 VINN.n113 4.5005
R66843 VINN.n235 VINN.n113 4.5005
R66844 VINN.n362 VINN.n113 4.5005
R66845 VINN.n234 VINN.n113 4.5005
R66846 VINN.n364 VINN.n113 4.5005
R66847 VINN.n233 VINN.n113 4.5005
R66848 VINN.n366 VINN.n113 4.5005
R66849 VINN.n232 VINN.n113 4.5005
R66850 VINN.n368 VINN.n113 4.5005
R66851 VINN.n231 VINN.n113 4.5005
R66852 VINN.n370 VINN.n113 4.5005
R66853 VINN.n230 VINN.n113 4.5005
R66854 VINN.n372 VINN.n113 4.5005
R66855 VINN.n229 VINN.n113 4.5005
R66856 VINN.n374 VINN.n113 4.5005
R66857 VINN.n228 VINN.n113 4.5005
R66858 VINN.n376 VINN.n113 4.5005
R66859 VINN.n227 VINN.n113 4.5005
R66860 VINN.n378 VINN.n113 4.5005
R66861 VINN.n226 VINN.n113 4.5005
R66862 VINN.n380 VINN.n113 4.5005
R66863 VINN.n225 VINN.n113 4.5005
R66864 VINN.n382 VINN.n113 4.5005
R66865 VINN.n224 VINN.n113 4.5005
R66866 VINN.n384 VINN.n113 4.5005
R66867 VINN.n223 VINN.n113 4.5005
R66868 VINN.n386 VINN.n113 4.5005
R66869 VINN.n222 VINN.n113 4.5005
R66870 VINN.n388 VINN.n113 4.5005
R66871 VINN.n221 VINN.n113 4.5005
R66872 VINN.n390 VINN.n113 4.5005
R66873 VINN.n220 VINN.n113 4.5005
R66874 VINN.n392 VINN.n113 4.5005
R66875 VINN.n219 VINN.n113 4.5005
R66876 VINN.n394 VINN.n113 4.5005
R66877 VINN.n218 VINN.n113 4.5005
R66878 VINN.n396 VINN.n113 4.5005
R66879 VINN.n217 VINN.n113 4.5005
R66880 VINN.n398 VINN.n113 4.5005
R66881 VINN.n216 VINN.n113 4.5005
R66882 VINN.n400 VINN.n113 4.5005
R66883 VINN.n215 VINN.n113 4.5005
R66884 VINN.n654 VINN.n113 4.5005
R66885 VINN.n656 VINN.n113 4.5005
R66886 VINN.n113 VINN.n0 4.5005
R66887 VINN.n278 VINN.n188 4.5005
R66888 VINN.n276 VINN.n188 4.5005
R66889 VINN.n280 VINN.n188 4.5005
R66890 VINN.n275 VINN.n188 4.5005
R66891 VINN.n282 VINN.n188 4.5005
R66892 VINN.n274 VINN.n188 4.5005
R66893 VINN.n284 VINN.n188 4.5005
R66894 VINN.n273 VINN.n188 4.5005
R66895 VINN.n286 VINN.n188 4.5005
R66896 VINN.n272 VINN.n188 4.5005
R66897 VINN.n288 VINN.n188 4.5005
R66898 VINN.n271 VINN.n188 4.5005
R66899 VINN.n290 VINN.n188 4.5005
R66900 VINN.n270 VINN.n188 4.5005
R66901 VINN.n292 VINN.n188 4.5005
R66902 VINN.n269 VINN.n188 4.5005
R66903 VINN.n294 VINN.n188 4.5005
R66904 VINN.n268 VINN.n188 4.5005
R66905 VINN.n296 VINN.n188 4.5005
R66906 VINN.n267 VINN.n188 4.5005
R66907 VINN.n298 VINN.n188 4.5005
R66908 VINN.n266 VINN.n188 4.5005
R66909 VINN.n300 VINN.n188 4.5005
R66910 VINN.n265 VINN.n188 4.5005
R66911 VINN.n302 VINN.n188 4.5005
R66912 VINN.n264 VINN.n188 4.5005
R66913 VINN.n304 VINN.n188 4.5005
R66914 VINN.n263 VINN.n188 4.5005
R66915 VINN.n306 VINN.n188 4.5005
R66916 VINN.n262 VINN.n188 4.5005
R66917 VINN.n308 VINN.n188 4.5005
R66918 VINN.n261 VINN.n188 4.5005
R66919 VINN.n310 VINN.n188 4.5005
R66920 VINN.n260 VINN.n188 4.5005
R66921 VINN.n312 VINN.n188 4.5005
R66922 VINN.n259 VINN.n188 4.5005
R66923 VINN.n314 VINN.n188 4.5005
R66924 VINN.n258 VINN.n188 4.5005
R66925 VINN.n316 VINN.n188 4.5005
R66926 VINN.n257 VINN.n188 4.5005
R66927 VINN.n318 VINN.n188 4.5005
R66928 VINN.n256 VINN.n188 4.5005
R66929 VINN.n320 VINN.n188 4.5005
R66930 VINN.n255 VINN.n188 4.5005
R66931 VINN.n322 VINN.n188 4.5005
R66932 VINN.n254 VINN.n188 4.5005
R66933 VINN.n324 VINN.n188 4.5005
R66934 VINN.n253 VINN.n188 4.5005
R66935 VINN.n326 VINN.n188 4.5005
R66936 VINN.n252 VINN.n188 4.5005
R66937 VINN.n328 VINN.n188 4.5005
R66938 VINN.n251 VINN.n188 4.5005
R66939 VINN.n330 VINN.n188 4.5005
R66940 VINN.n250 VINN.n188 4.5005
R66941 VINN.n332 VINN.n188 4.5005
R66942 VINN.n249 VINN.n188 4.5005
R66943 VINN.n334 VINN.n188 4.5005
R66944 VINN.n248 VINN.n188 4.5005
R66945 VINN.n336 VINN.n188 4.5005
R66946 VINN.n247 VINN.n188 4.5005
R66947 VINN.n338 VINN.n188 4.5005
R66948 VINN.n246 VINN.n188 4.5005
R66949 VINN.n340 VINN.n188 4.5005
R66950 VINN.n245 VINN.n188 4.5005
R66951 VINN.n342 VINN.n188 4.5005
R66952 VINN.n244 VINN.n188 4.5005
R66953 VINN.n344 VINN.n188 4.5005
R66954 VINN.n243 VINN.n188 4.5005
R66955 VINN.n346 VINN.n188 4.5005
R66956 VINN.n242 VINN.n188 4.5005
R66957 VINN.n348 VINN.n188 4.5005
R66958 VINN.n241 VINN.n188 4.5005
R66959 VINN.n350 VINN.n188 4.5005
R66960 VINN.n240 VINN.n188 4.5005
R66961 VINN.n352 VINN.n188 4.5005
R66962 VINN.n239 VINN.n188 4.5005
R66963 VINN.n354 VINN.n188 4.5005
R66964 VINN.n238 VINN.n188 4.5005
R66965 VINN.n356 VINN.n188 4.5005
R66966 VINN.n237 VINN.n188 4.5005
R66967 VINN.n358 VINN.n188 4.5005
R66968 VINN.n236 VINN.n188 4.5005
R66969 VINN.n360 VINN.n188 4.5005
R66970 VINN.n235 VINN.n188 4.5005
R66971 VINN.n362 VINN.n188 4.5005
R66972 VINN.n234 VINN.n188 4.5005
R66973 VINN.n364 VINN.n188 4.5005
R66974 VINN.n233 VINN.n188 4.5005
R66975 VINN.n366 VINN.n188 4.5005
R66976 VINN.n232 VINN.n188 4.5005
R66977 VINN.n368 VINN.n188 4.5005
R66978 VINN.n231 VINN.n188 4.5005
R66979 VINN.n370 VINN.n188 4.5005
R66980 VINN.n230 VINN.n188 4.5005
R66981 VINN.n372 VINN.n188 4.5005
R66982 VINN.n229 VINN.n188 4.5005
R66983 VINN.n374 VINN.n188 4.5005
R66984 VINN.n228 VINN.n188 4.5005
R66985 VINN.n376 VINN.n188 4.5005
R66986 VINN.n227 VINN.n188 4.5005
R66987 VINN.n378 VINN.n188 4.5005
R66988 VINN.n226 VINN.n188 4.5005
R66989 VINN.n380 VINN.n188 4.5005
R66990 VINN.n225 VINN.n188 4.5005
R66991 VINN.n382 VINN.n188 4.5005
R66992 VINN.n224 VINN.n188 4.5005
R66993 VINN.n384 VINN.n188 4.5005
R66994 VINN.n223 VINN.n188 4.5005
R66995 VINN.n386 VINN.n188 4.5005
R66996 VINN.n222 VINN.n188 4.5005
R66997 VINN.n388 VINN.n188 4.5005
R66998 VINN.n221 VINN.n188 4.5005
R66999 VINN.n390 VINN.n188 4.5005
R67000 VINN.n220 VINN.n188 4.5005
R67001 VINN.n392 VINN.n188 4.5005
R67002 VINN.n219 VINN.n188 4.5005
R67003 VINN.n394 VINN.n188 4.5005
R67004 VINN.n218 VINN.n188 4.5005
R67005 VINN.n396 VINN.n188 4.5005
R67006 VINN.n217 VINN.n188 4.5005
R67007 VINN.n398 VINN.n188 4.5005
R67008 VINN.n216 VINN.n188 4.5005
R67009 VINN.n400 VINN.n188 4.5005
R67010 VINN.n215 VINN.n188 4.5005
R67011 VINN.n654 VINN.n188 4.5005
R67012 VINN.n656 VINN.n188 4.5005
R67013 VINN.n188 VINN.n0 4.5005
R67014 VINN.n278 VINN.n112 4.5005
R67015 VINN.n276 VINN.n112 4.5005
R67016 VINN.n280 VINN.n112 4.5005
R67017 VINN.n275 VINN.n112 4.5005
R67018 VINN.n282 VINN.n112 4.5005
R67019 VINN.n274 VINN.n112 4.5005
R67020 VINN.n284 VINN.n112 4.5005
R67021 VINN.n273 VINN.n112 4.5005
R67022 VINN.n286 VINN.n112 4.5005
R67023 VINN.n272 VINN.n112 4.5005
R67024 VINN.n288 VINN.n112 4.5005
R67025 VINN.n271 VINN.n112 4.5005
R67026 VINN.n290 VINN.n112 4.5005
R67027 VINN.n270 VINN.n112 4.5005
R67028 VINN.n292 VINN.n112 4.5005
R67029 VINN.n269 VINN.n112 4.5005
R67030 VINN.n294 VINN.n112 4.5005
R67031 VINN.n268 VINN.n112 4.5005
R67032 VINN.n296 VINN.n112 4.5005
R67033 VINN.n267 VINN.n112 4.5005
R67034 VINN.n298 VINN.n112 4.5005
R67035 VINN.n266 VINN.n112 4.5005
R67036 VINN.n300 VINN.n112 4.5005
R67037 VINN.n265 VINN.n112 4.5005
R67038 VINN.n302 VINN.n112 4.5005
R67039 VINN.n264 VINN.n112 4.5005
R67040 VINN.n304 VINN.n112 4.5005
R67041 VINN.n263 VINN.n112 4.5005
R67042 VINN.n306 VINN.n112 4.5005
R67043 VINN.n262 VINN.n112 4.5005
R67044 VINN.n308 VINN.n112 4.5005
R67045 VINN.n261 VINN.n112 4.5005
R67046 VINN.n310 VINN.n112 4.5005
R67047 VINN.n260 VINN.n112 4.5005
R67048 VINN.n312 VINN.n112 4.5005
R67049 VINN.n259 VINN.n112 4.5005
R67050 VINN.n314 VINN.n112 4.5005
R67051 VINN.n258 VINN.n112 4.5005
R67052 VINN.n316 VINN.n112 4.5005
R67053 VINN.n257 VINN.n112 4.5005
R67054 VINN.n318 VINN.n112 4.5005
R67055 VINN.n256 VINN.n112 4.5005
R67056 VINN.n320 VINN.n112 4.5005
R67057 VINN.n255 VINN.n112 4.5005
R67058 VINN.n322 VINN.n112 4.5005
R67059 VINN.n254 VINN.n112 4.5005
R67060 VINN.n324 VINN.n112 4.5005
R67061 VINN.n253 VINN.n112 4.5005
R67062 VINN.n326 VINN.n112 4.5005
R67063 VINN.n252 VINN.n112 4.5005
R67064 VINN.n328 VINN.n112 4.5005
R67065 VINN.n251 VINN.n112 4.5005
R67066 VINN.n330 VINN.n112 4.5005
R67067 VINN.n250 VINN.n112 4.5005
R67068 VINN.n332 VINN.n112 4.5005
R67069 VINN.n249 VINN.n112 4.5005
R67070 VINN.n334 VINN.n112 4.5005
R67071 VINN.n248 VINN.n112 4.5005
R67072 VINN.n336 VINN.n112 4.5005
R67073 VINN.n247 VINN.n112 4.5005
R67074 VINN.n338 VINN.n112 4.5005
R67075 VINN.n246 VINN.n112 4.5005
R67076 VINN.n340 VINN.n112 4.5005
R67077 VINN.n245 VINN.n112 4.5005
R67078 VINN.n342 VINN.n112 4.5005
R67079 VINN.n244 VINN.n112 4.5005
R67080 VINN.n344 VINN.n112 4.5005
R67081 VINN.n243 VINN.n112 4.5005
R67082 VINN.n346 VINN.n112 4.5005
R67083 VINN.n242 VINN.n112 4.5005
R67084 VINN.n348 VINN.n112 4.5005
R67085 VINN.n241 VINN.n112 4.5005
R67086 VINN.n350 VINN.n112 4.5005
R67087 VINN.n240 VINN.n112 4.5005
R67088 VINN.n352 VINN.n112 4.5005
R67089 VINN.n239 VINN.n112 4.5005
R67090 VINN.n354 VINN.n112 4.5005
R67091 VINN.n238 VINN.n112 4.5005
R67092 VINN.n356 VINN.n112 4.5005
R67093 VINN.n237 VINN.n112 4.5005
R67094 VINN.n358 VINN.n112 4.5005
R67095 VINN.n236 VINN.n112 4.5005
R67096 VINN.n360 VINN.n112 4.5005
R67097 VINN.n235 VINN.n112 4.5005
R67098 VINN.n362 VINN.n112 4.5005
R67099 VINN.n234 VINN.n112 4.5005
R67100 VINN.n364 VINN.n112 4.5005
R67101 VINN.n233 VINN.n112 4.5005
R67102 VINN.n366 VINN.n112 4.5005
R67103 VINN.n232 VINN.n112 4.5005
R67104 VINN.n368 VINN.n112 4.5005
R67105 VINN.n231 VINN.n112 4.5005
R67106 VINN.n370 VINN.n112 4.5005
R67107 VINN.n230 VINN.n112 4.5005
R67108 VINN.n372 VINN.n112 4.5005
R67109 VINN.n229 VINN.n112 4.5005
R67110 VINN.n374 VINN.n112 4.5005
R67111 VINN.n228 VINN.n112 4.5005
R67112 VINN.n376 VINN.n112 4.5005
R67113 VINN.n227 VINN.n112 4.5005
R67114 VINN.n378 VINN.n112 4.5005
R67115 VINN.n226 VINN.n112 4.5005
R67116 VINN.n380 VINN.n112 4.5005
R67117 VINN.n225 VINN.n112 4.5005
R67118 VINN.n382 VINN.n112 4.5005
R67119 VINN.n224 VINN.n112 4.5005
R67120 VINN.n384 VINN.n112 4.5005
R67121 VINN.n223 VINN.n112 4.5005
R67122 VINN.n386 VINN.n112 4.5005
R67123 VINN.n222 VINN.n112 4.5005
R67124 VINN.n388 VINN.n112 4.5005
R67125 VINN.n221 VINN.n112 4.5005
R67126 VINN.n390 VINN.n112 4.5005
R67127 VINN.n220 VINN.n112 4.5005
R67128 VINN.n392 VINN.n112 4.5005
R67129 VINN.n219 VINN.n112 4.5005
R67130 VINN.n394 VINN.n112 4.5005
R67131 VINN.n218 VINN.n112 4.5005
R67132 VINN.n396 VINN.n112 4.5005
R67133 VINN.n217 VINN.n112 4.5005
R67134 VINN.n398 VINN.n112 4.5005
R67135 VINN.n216 VINN.n112 4.5005
R67136 VINN.n400 VINN.n112 4.5005
R67137 VINN.n215 VINN.n112 4.5005
R67138 VINN.n654 VINN.n112 4.5005
R67139 VINN.n656 VINN.n112 4.5005
R67140 VINN.n112 VINN.n0 4.5005
R67141 VINN.n278 VINN.n189 4.5005
R67142 VINN.n276 VINN.n189 4.5005
R67143 VINN.n280 VINN.n189 4.5005
R67144 VINN.n275 VINN.n189 4.5005
R67145 VINN.n282 VINN.n189 4.5005
R67146 VINN.n274 VINN.n189 4.5005
R67147 VINN.n284 VINN.n189 4.5005
R67148 VINN.n273 VINN.n189 4.5005
R67149 VINN.n286 VINN.n189 4.5005
R67150 VINN.n272 VINN.n189 4.5005
R67151 VINN.n288 VINN.n189 4.5005
R67152 VINN.n271 VINN.n189 4.5005
R67153 VINN.n290 VINN.n189 4.5005
R67154 VINN.n270 VINN.n189 4.5005
R67155 VINN.n292 VINN.n189 4.5005
R67156 VINN.n269 VINN.n189 4.5005
R67157 VINN.n294 VINN.n189 4.5005
R67158 VINN.n268 VINN.n189 4.5005
R67159 VINN.n296 VINN.n189 4.5005
R67160 VINN.n267 VINN.n189 4.5005
R67161 VINN.n298 VINN.n189 4.5005
R67162 VINN.n266 VINN.n189 4.5005
R67163 VINN.n300 VINN.n189 4.5005
R67164 VINN.n265 VINN.n189 4.5005
R67165 VINN.n302 VINN.n189 4.5005
R67166 VINN.n264 VINN.n189 4.5005
R67167 VINN.n304 VINN.n189 4.5005
R67168 VINN.n263 VINN.n189 4.5005
R67169 VINN.n306 VINN.n189 4.5005
R67170 VINN.n262 VINN.n189 4.5005
R67171 VINN.n308 VINN.n189 4.5005
R67172 VINN.n261 VINN.n189 4.5005
R67173 VINN.n310 VINN.n189 4.5005
R67174 VINN.n260 VINN.n189 4.5005
R67175 VINN.n312 VINN.n189 4.5005
R67176 VINN.n259 VINN.n189 4.5005
R67177 VINN.n314 VINN.n189 4.5005
R67178 VINN.n258 VINN.n189 4.5005
R67179 VINN.n316 VINN.n189 4.5005
R67180 VINN.n257 VINN.n189 4.5005
R67181 VINN.n318 VINN.n189 4.5005
R67182 VINN.n256 VINN.n189 4.5005
R67183 VINN.n320 VINN.n189 4.5005
R67184 VINN.n255 VINN.n189 4.5005
R67185 VINN.n322 VINN.n189 4.5005
R67186 VINN.n254 VINN.n189 4.5005
R67187 VINN.n324 VINN.n189 4.5005
R67188 VINN.n253 VINN.n189 4.5005
R67189 VINN.n326 VINN.n189 4.5005
R67190 VINN.n252 VINN.n189 4.5005
R67191 VINN.n328 VINN.n189 4.5005
R67192 VINN.n251 VINN.n189 4.5005
R67193 VINN.n330 VINN.n189 4.5005
R67194 VINN.n250 VINN.n189 4.5005
R67195 VINN.n332 VINN.n189 4.5005
R67196 VINN.n249 VINN.n189 4.5005
R67197 VINN.n334 VINN.n189 4.5005
R67198 VINN.n248 VINN.n189 4.5005
R67199 VINN.n336 VINN.n189 4.5005
R67200 VINN.n247 VINN.n189 4.5005
R67201 VINN.n338 VINN.n189 4.5005
R67202 VINN.n246 VINN.n189 4.5005
R67203 VINN.n340 VINN.n189 4.5005
R67204 VINN.n245 VINN.n189 4.5005
R67205 VINN.n342 VINN.n189 4.5005
R67206 VINN.n244 VINN.n189 4.5005
R67207 VINN.n344 VINN.n189 4.5005
R67208 VINN.n243 VINN.n189 4.5005
R67209 VINN.n346 VINN.n189 4.5005
R67210 VINN.n242 VINN.n189 4.5005
R67211 VINN.n348 VINN.n189 4.5005
R67212 VINN.n241 VINN.n189 4.5005
R67213 VINN.n350 VINN.n189 4.5005
R67214 VINN.n240 VINN.n189 4.5005
R67215 VINN.n352 VINN.n189 4.5005
R67216 VINN.n239 VINN.n189 4.5005
R67217 VINN.n354 VINN.n189 4.5005
R67218 VINN.n238 VINN.n189 4.5005
R67219 VINN.n356 VINN.n189 4.5005
R67220 VINN.n237 VINN.n189 4.5005
R67221 VINN.n358 VINN.n189 4.5005
R67222 VINN.n236 VINN.n189 4.5005
R67223 VINN.n360 VINN.n189 4.5005
R67224 VINN.n235 VINN.n189 4.5005
R67225 VINN.n362 VINN.n189 4.5005
R67226 VINN.n234 VINN.n189 4.5005
R67227 VINN.n364 VINN.n189 4.5005
R67228 VINN.n233 VINN.n189 4.5005
R67229 VINN.n366 VINN.n189 4.5005
R67230 VINN.n232 VINN.n189 4.5005
R67231 VINN.n368 VINN.n189 4.5005
R67232 VINN.n231 VINN.n189 4.5005
R67233 VINN.n370 VINN.n189 4.5005
R67234 VINN.n230 VINN.n189 4.5005
R67235 VINN.n372 VINN.n189 4.5005
R67236 VINN.n229 VINN.n189 4.5005
R67237 VINN.n374 VINN.n189 4.5005
R67238 VINN.n228 VINN.n189 4.5005
R67239 VINN.n376 VINN.n189 4.5005
R67240 VINN.n227 VINN.n189 4.5005
R67241 VINN.n378 VINN.n189 4.5005
R67242 VINN.n226 VINN.n189 4.5005
R67243 VINN.n380 VINN.n189 4.5005
R67244 VINN.n225 VINN.n189 4.5005
R67245 VINN.n382 VINN.n189 4.5005
R67246 VINN.n224 VINN.n189 4.5005
R67247 VINN.n384 VINN.n189 4.5005
R67248 VINN.n223 VINN.n189 4.5005
R67249 VINN.n386 VINN.n189 4.5005
R67250 VINN.n222 VINN.n189 4.5005
R67251 VINN.n388 VINN.n189 4.5005
R67252 VINN.n221 VINN.n189 4.5005
R67253 VINN.n390 VINN.n189 4.5005
R67254 VINN.n220 VINN.n189 4.5005
R67255 VINN.n392 VINN.n189 4.5005
R67256 VINN.n219 VINN.n189 4.5005
R67257 VINN.n394 VINN.n189 4.5005
R67258 VINN.n218 VINN.n189 4.5005
R67259 VINN.n396 VINN.n189 4.5005
R67260 VINN.n217 VINN.n189 4.5005
R67261 VINN.n398 VINN.n189 4.5005
R67262 VINN.n216 VINN.n189 4.5005
R67263 VINN.n400 VINN.n189 4.5005
R67264 VINN.n215 VINN.n189 4.5005
R67265 VINN.n654 VINN.n189 4.5005
R67266 VINN.n656 VINN.n189 4.5005
R67267 VINN.n189 VINN.n0 4.5005
R67268 VINN.n278 VINN.n111 4.5005
R67269 VINN.n276 VINN.n111 4.5005
R67270 VINN.n280 VINN.n111 4.5005
R67271 VINN.n275 VINN.n111 4.5005
R67272 VINN.n282 VINN.n111 4.5005
R67273 VINN.n274 VINN.n111 4.5005
R67274 VINN.n284 VINN.n111 4.5005
R67275 VINN.n273 VINN.n111 4.5005
R67276 VINN.n286 VINN.n111 4.5005
R67277 VINN.n272 VINN.n111 4.5005
R67278 VINN.n288 VINN.n111 4.5005
R67279 VINN.n271 VINN.n111 4.5005
R67280 VINN.n290 VINN.n111 4.5005
R67281 VINN.n270 VINN.n111 4.5005
R67282 VINN.n292 VINN.n111 4.5005
R67283 VINN.n269 VINN.n111 4.5005
R67284 VINN.n294 VINN.n111 4.5005
R67285 VINN.n268 VINN.n111 4.5005
R67286 VINN.n296 VINN.n111 4.5005
R67287 VINN.n267 VINN.n111 4.5005
R67288 VINN.n298 VINN.n111 4.5005
R67289 VINN.n266 VINN.n111 4.5005
R67290 VINN.n300 VINN.n111 4.5005
R67291 VINN.n265 VINN.n111 4.5005
R67292 VINN.n302 VINN.n111 4.5005
R67293 VINN.n264 VINN.n111 4.5005
R67294 VINN.n304 VINN.n111 4.5005
R67295 VINN.n263 VINN.n111 4.5005
R67296 VINN.n306 VINN.n111 4.5005
R67297 VINN.n262 VINN.n111 4.5005
R67298 VINN.n308 VINN.n111 4.5005
R67299 VINN.n261 VINN.n111 4.5005
R67300 VINN.n310 VINN.n111 4.5005
R67301 VINN.n260 VINN.n111 4.5005
R67302 VINN.n312 VINN.n111 4.5005
R67303 VINN.n259 VINN.n111 4.5005
R67304 VINN.n314 VINN.n111 4.5005
R67305 VINN.n258 VINN.n111 4.5005
R67306 VINN.n316 VINN.n111 4.5005
R67307 VINN.n257 VINN.n111 4.5005
R67308 VINN.n318 VINN.n111 4.5005
R67309 VINN.n256 VINN.n111 4.5005
R67310 VINN.n320 VINN.n111 4.5005
R67311 VINN.n255 VINN.n111 4.5005
R67312 VINN.n322 VINN.n111 4.5005
R67313 VINN.n254 VINN.n111 4.5005
R67314 VINN.n324 VINN.n111 4.5005
R67315 VINN.n253 VINN.n111 4.5005
R67316 VINN.n326 VINN.n111 4.5005
R67317 VINN.n252 VINN.n111 4.5005
R67318 VINN.n328 VINN.n111 4.5005
R67319 VINN.n251 VINN.n111 4.5005
R67320 VINN.n330 VINN.n111 4.5005
R67321 VINN.n250 VINN.n111 4.5005
R67322 VINN.n332 VINN.n111 4.5005
R67323 VINN.n249 VINN.n111 4.5005
R67324 VINN.n334 VINN.n111 4.5005
R67325 VINN.n248 VINN.n111 4.5005
R67326 VINN.n336 VINN.n111 4.5005
R67327 VINN.n247 VINN.n111 4.5005
R67328 VINN.n338 VINN.n111 4.5005
R67329 VINN.n246 VINN.n111 4.5005
R67330 VINN.n340 VINN.n111 4.5005
R67331 VINN.n245 VINN.n111 4.5005
R67332 VINN.n342 VINN.n111 4.5005
R67333 VINN.n244 VINN.n111 4.5005
R67334 VINN.n344 VINN.n111 4.5005
R67335 VINN.n243 VINN.n111 4.5005
R67336 VINN.n346 VINN.n111 4.5005
R67337 VINN.n242 VINN.n111 4.5005
R67338 VINN.n348 VINN.n111 4.5005
R67339 VINN.n241 VINN.n111 4.5005
R67340 VINN.n350 VINN.n111 4.5005
R67341 VINN.n240 VINN.n111 4.5005
R67342 VINN.n352 VINN.n111 4.5005
R67343 VINN.n239 VINN.n111 4.5005
R67344 VINN.n354 VINN.n111 4.5005
R67345 VINN.n238 VINN.n111 4.5005
R67346 VINN.n356 VINN.n111 4.5005
R67347 VINN.n237 VINN.n111 4.5005
R67348 VINN.n358 VINN.n111 4.5005
R67349 VINN.n236 VINN.n111 4.5005
R67350 VINN.n360 VINN.n111 4.5005
R67351 VINN.n235 VINN.n111 4.5005
R67352 VINN.n362 VINN.n111 4.5005
R67353 VINN.n234 VINN.n111 4.5005
R67354 VINN.n364 VINN.n111 4.5005
R67355 VINN.n233 VINN.n111 4.5005
R67356 VINN.n366 VINN.n111 4.5005
R67357 VINN.n232 VINN.n111 4.5005
R67358 VINN.n368 VINN.n111 4.5005
R67359 VINN.n231 VINN.n111 4.5005
R67360 VINN.n370 VINN.n111 4.5005
R67361 VINN.n230 VINN.n111 4.5005
R67362 VINN.n372 VINN.n111 4.5005
R67363 VINN.n229 VINN.n111 4.5005
R67364 VINN.n374 VINN.n111 4.5005
R67365 VINN.n228 VINN.n111 4.5005
R67366 VINN.n376 VINN.n111 4.5005
R67367 VINN.n227 VINN.n111 4.5005
R67368 VINN.n378 VINN.n111 4.5005
R67369 VINN.n226 VINN.n111 4.5005
R67370 VINN.n380 VINN.n111 4.5005
R67371 VINN.n225 VINN.n111 4.5005
R67372 VINN.n382 VINN.n111 4.5005
R67373 VINN.n224 VINN.n111 4.5005
R67374 VINN.n384 VINN.n111 4.5005
R67375 VINN.n223 VINN.n111 4.5005
R67376 VINN.n386 VINN.n111 4.5005
R67377 VINN.n222 VINN.n111 4.5005
R67378 VINN.n388 VINN.n111 4.5005
R67379 VINN.n221 VINN.n111 4.5005
R67380 VINN.n390 VINN.n111 4.5005
R67381 VINN.n220 VINN.n111 4.5005
R67382 VINN.n392 VINN.n111 4.5005
R67383 VINN.n219 VINN.n111 4.5005
R67384 VINN.n394 VINN.n111 4.5005
R67385 VINN.n218 VINN.n111 4.5005
R67386 VINN.n396 VINN.n111 4.5005
R67387 VINN.n217 VINN.n111 4.5005
R67388 VINN.n398 VINN.n111 4.5005
R67389 VINN.n216 VINN.n111 4.5005
R67390 VINN.n400 VINN.n111 4.5005
R67391 VINN.n215 VINN.n111 4.5005
R67392 VINN.n654 VINN.n111 4.5005
R67393 VINN.n656 VINN.n111 4.5005
R67394 VINN.n111 VINN.n0 4.5005
R67395 VINN.n278 VINN.n190 4.5005
R67396 VINN.n276 VINN.n190 4.5005
R67397 VINN.n280 VINN.n190 4.5005
R67398 VINN.n275 VINN.n190 4.5005
R67399 VINN.n282 VINN.n190 4.5005
R67400 VINN.n274 VINN.n190 4.5005
R67401 VINN.n284 VINN.n190 4.5005
R67402 VINN.n273 VINN.n190 4.5005
R67403 VINN.n286 VINN.n190 4.5005
R67404 VINN.n272 VINN.n190 4.5005
R67405 VINN.n288 VINN.n190 4.5005
R67406 VINN.n271 VINN.n190 4.5005
R67407 VINN.n290 VINN.n190 4.5005
R67408 VINN.n270 VINN.n190 4.5005
R67409 VINN.n292 VINN.n190 4.5005
R67410 VINN.n269 VINN.n190 4.5005
R67411 VINN.n294 VINN.n190 4.5005
R67412 VINN.n268 VINN.n190 4.5005
R67413 VINN.n296 VINN.n190 4.5005
R67414 VINN.n267 VINN.n190 4.5005
R67415 VINN.n298 VINN.n190 4.5005
R67416 VINN.n266 VINN.n190 4.5005
R67417 VINN.n300 VINN.n190 4.5005
R67418 VINN.n265 VINN.n190 4.5005
R67419 VINN.n302 VINN.n190 4.5005
R67420 VINN.n264 VINN.n190 4.5005
R67421 VINN.n304 VINN.n190 4.5005
R67422 VINN.n263 VINN.n190 4.5005
R67423 VINN.n306 VINN.n190 4.5005
R67424 VINN.n262 VINN.n190 4.5005
R67425 VINN.n308 VINN.n190 4.5005
R67426 VINN.n261 VINN.n190 4.5005
R67427 VINN.n310 VINN.n190 4.5005
R67428 VINN.n260 VINN.n190 4.5005
R67429 VINN.n312 VINN.n190 4.5005
R67430 VINN.n259 VINN.n190 4.5005
R67431 VINN.n314 VINN.n190 4.5005
R67432 VINN.n258 VINN.n190 4.5005
R67433 VINN.n316 VINN.n190 4.5005
R67434 VINN.n257 VINN.n190 4.5005
R67435 VINN.n318 VINN.n190 4.5005
R67436 VINN.n256 VINN.n190 4.5005
R67437 VINN.n320 VINN.n190 4.5005
R67438 VINN.n255 VINN.n190 4.5005
R67439 VINN.n322 VINN.n190 4.5005
R67440 VINN.n254 VINN.n190 4.5005
R67441 VINN.n324 VINN.n190 4.5005
R67442 VINN.n253 VINN.n190 4.5005
R67443 VINN.n326 VINN.n190 4.5005
R67444 VINN.n252 VINN.n190 4.5005
R67445 VINN.n328 VINN.n190 4.5005
R67446 VINN.n251 VINN.n190 4.5005
R67447 VINN.n330 VINN.n190 4.5005
R67448 VINN.n250 VINN.n190 4.5005
R67449 VINN.n332 VINN.n190 4.5005
R67450 VINN.n249 VINN.n190 4.5005
R67451 VINN.n334 VINN.n190 4.5005
R67452 VINN.n248 VINN.n190 4.5005
R67453 VINN.n336 VINN.n190 4.5005
R67454 VINN.n247 VINN.n190 4.5005
R67455 VINN.n338 VINN.n190 4.5005
R67456 VINN.n246 VINN.n190 4.5005
R67457 VINN.n340 VINN.n190 4.5005
R67458 VINN.n245 VINN.n190 4.5005
R67459 VINN.n342 VINN.n190 4.5005
R67460 VINN.n244 VINN.n190 4.5005
R67461 VINN.n344 VINN.n190 4.5005
R67462 VINN.n243 VINN.n190 4.5005
R67463 VINN.n346 VINN.n190 4.5005
R67464 VINN.n242 VINN.n190 4.5005
R67465 VINN.n348 VINN.n190 4.5005
R67466 VINN.n241 VINN.n190 4.5005
R67467 VINN.n350 VINN.n190 4.5005
R67468 VINN.n240 VINN.n190 4.5005
R67469 VINN.n352 VINN.n190 4.5005
R67470 VINN.n239 VINN.n190 4.5005
R67471 VINN.n354 VINN.n190 4.5005
R67472 VINN.n238 VINN.n190 4.5005
R67473 VINN.n356 VINN.n190 4.5005
R67474 VINN.n237 VINN.n190 4.5005
R67475 VINN.n358 VINN.n190 4.5005
R67476 VINN.n236 VINN.n190 4.5005
R67477 VINN.n360 VINN.n190 4.5005
R67478 VINN.n235 VINN.n190 4.5005
R67479 VINN.n362 VINN.n190 4.5005
R67480 VINN.n234 VINN.n190 4.5005
R67481 VINN.n364 VINN.n190 4.5005
R67482 VINN.n233 VINN.n190 4.5005
R67483 VINN.n366 VINN.n190 4.5005
R67484 VINN.n232 VINN.n190 4.5005
R67485 VINN.n368 VINN.n190 4.5005
R67486 VINN.n231 VINN.n190 4.5005
R67487 VINN.n370 VINN.n190 4.5005
R67488 VINN.n230 VINN.n190 4.5005
R67489 VINN.n372 VINN.n190 4.5005
R67490 VINN.n229 VINN.n190 4.5005
R67491 VINN.n374 VINN.n190 4.5005
R67492 VINN.n228 VINN.n190 4.5005
R67493 VINN.n376 VINN.n190 4.5005
R67494 VINN.n227 VINN.n190 4.5005
R67495 VINN.n378 VINN.n190 4.5005
R67496 VINN.n226 VINN.n190 4.5005
R67497 VINN.n380 VINN.n190 4.5005
R67498 VINN.n225 VINN.n190 4.5005
R67499 VINN.n382 VINN.n190 4.5005
R67500 VINN.n224 VINN.n190 4.5005
R67501 VINN.n384 VINN.n190 4.5005
R67502 VINN.n223 VINN.n190 4.5005
R67503 VINN.n386 VINN.n190 4.5005
R67504 VINN.n222 VINN.n190 4.5005
R67505 VINN.n388 VINN.n190 4.5005
R67506 VINN.n221 VINN.n190 4.5005
R67507 VINN.n390 VINN.n190 4.5005
R67508 VINN.n220 VINN.n190 4.5005
R67509 VINN.n392 VINN.n190 4.5005
R67510 VINN.n219 VINN.n190 4.5005
R67511 VINN.n394 VINN.n190 4.5005
R67512 VINN.n218 VINN.n190 4.5005
R67513 VINN.n396 VINN.n190 4.5005
R67514 VINN.n217 VINN.n190 4.5005
R67515 VINN.n398 VINN.n190 4.5005
R67516 VINN.n216 VINN.n190 4.5005
R67517 VINN.n400 VINN.n190 4.5005
R67518 VINN.n215 VINN.n190 4.5005
R67519 VINN.n654 VINN.n190 4.5005
R67520 VINN.n656 VINN.n190 4.5005
R67521 VINN.n190 VINN.n0 4.5005
R67522 VINN.n278 VINN.n110 4.5005
R67523 VINN.n276 VINN.n110 4.5005
R67524 VINN.n280 VINN.n110 4.5005
R67525 VINN.n275 VINN.n110 4.5005
R67526 VINN.n282 VINN.n110 4.5005
R67527 VINN.n274 VINN.n110 4.5005
R67528 VINN.n284 VINN.n110 4.5005
R67529 VINN.n273 VINN.n110 4.5005
R67530 VINN.n286 VINN.n110 4.5005
R67531 VINN.n272 VINN.n110 4.5005
R67532 VINN.n288 VINN.n110 4.5005
R67533 VINN.n271 VINN.n110 4.5005
R67534 VINN.n290 VINN.n110 4.5005
R67535 VINN.n270 VINN.n110 4.5005
R67536 VINN.n292 VINN.n110 4.5005
R67537 VINN.n269 VINN.n110 4.5005
R67538 VINN.n294 VINN.n110 4.5005
R67539 VINN.n268 VINN.n110 4.5005
R67540 VINN.n296 VINN.n110 4.5005
R67541 VINN.n267 VINN.n110 4.5005
R67542 VINN.n298 VINN.n110 4.5005
R67543 VINN.n266 VINN.n110 4.5005
R67544 VINN.n300 VINN.n110 4.5005
R67545 VINN.n265 VINN.n110 4.5005
R67546 VINN.n302 VINN.n110 4.5005
R67547 VINN.n264 VINN.n110 4.5005
R67548 VINN.n304 VINN.n110 4.5005
R67549 VINN.n263 VINN.n110 4.5005
R67550 VINN.n306 VINN.n110 4.5005
R67551 VINN.n262 VINN.n110 4.5005
R67552 VINN.n308 VINN.n110 4.5005
R67553 VINN.n261 VINN.n110 4.5005
R67554 VINN.n310 VINN.n110 4.5005
R67555 VINN.n260 VINN.n110 4.5005
R67556 VINN.n312 VINN.n110 4.5005
R67557 VINN.n259 VINN.n110 4.5005
R67558 VINN.n314 VINN.n110 4.5005
R67559 VINN.n258 VINN.n110 4.5005
R67560 VINN.n316 VINN.n110 4.5005
R67561 VINN.n257 VINN.n110 4.5005
R67562 VINN.n318 VINN.n110 4.5005
R67563 VINN.n256 VINN.n110 4.5005
R67564 VINN.n320 VINN.n110 4.5005
R67565 VINN.n255 VINN.n110 4.5005
R67566 VINN.n322 VINN.n110 4.5005
R67567 VINN.n254 VINN.n110 4.5005
R67568 VINN.n324 VINN.n110 4.5005
R67569 VINN.n253 VINN.n110 4.5005
R67570 VINN.n326 VINN.n110 4.5005
R67571 VINN.n252 VINN.n110 4.5005
R67572 VINN.n328 VINN.n110 4.5005
R67573 VINN.n251 VINN.n110 4.5005
R67574 VINN.n330 VINN.n110 4.5005
R67575 VINN.n250 VINN.n110 4.5005
R67576 VINN.n332 VINN.n110 4.5005
R67577 VINN.n249 VINN.n110 4.5005
R67578 VINN.n334 VINN.n110 4.5005
R67579 VINN.n248 VINN.n110 4.5005
R67580 VINN.n336 VINN.n110 4.5005
R67581 VINN.n247 VINN.n110 4.5005
R67582 VINN.n338 VINN.n110 4.5005
R67583 VINN.n246 VINN.n110 4.5005
R67584 VINN.n340 VINN.n110 4.5005
R67585 VINN.n245 VINN.n110 4.5005
R67586 VINN.n342 VINN.n110 4.5005
R67587 VINN.n244 VINN.n110 4.5005
R67588 VINN.n344 VINN.n110 4.5005
R67589 VINN.n243 VINN.n110 4.5005
R67590 VINN.n346 VINN.n110 4.5005
R67591 VINN.n242 VINN.n110 4.5005
R67592 VINN.n348 VINN.n110 4.5005
R67593 VINN.n241 VINN.n110 4.5005
R67594 VINN.n350 VINN.n110 4.5005
R67595 VINN.n240 VINN.n110 4.5005
R67596 VINN.n352 VINN.n110 4.5005
R67597 VINN.n239 VINN.n110 4.5005
R67598 VINN.n354 VINN.n110 4.5005
R67599 VINN.n238 VINN.n110 4.5005
R67600 VINN.n356 VINN.n110 4.5005
R67601 VINN.n237 VINN.n110 4.5005
R67602 VINN.n358 VINN.n110 4.5005
R67603 VINN.n236 VINN.n110 4.5005
R67604 VINN.n360 VINN.n110 4.5005
R67605 VINN.n235 VINN.n110 4.5005
R67606 VINN.n362 VINN.n110 4.5005
R67607 VINN.n234 VINN.n110 4.5005
R67608 VINN.n364 VINN.n110 4.5005
R67609 VINN.n233 VINN.n110 4.5005
R67610 VINN.n366 VINN.n110 4.5005
R67611 VINN.n232 VINN.n110 4.5005
R67612 VINN.n368 VINN.n110 4.5005
R67613 VINN.n231 VINN.n110 4.5005
R67614 VINN.n370 VINN.n110 4.5005
R67615 VINN.n230 VINN.n110 4.5005
R67616 VINN.n372 VINN.n110 4.5005
R67617 VINN.n229 VINN.n110 4.5005
R67618 VINN.n374 VINN.n110 4.5005
R67619 VINN.n228 VINN.n110 4.5005
R67620 VINN.n376 VINN.n110 4.5005
R67621 VINN.n227 VINN.n110 4.5005
R67622 VINN.n378 VINN.n110 4.5005
R67623 VINN.n226 VINN.n110 4.5005
R67624 VINN.n380 VINN.n110 4.5005
R67625 VINN.n225 VINN.n110 4.5005
R67626 VINN.n382 VINN.n110 4.5005
R67627 VINN.n224 VINN.n110 4.5005
R67628 VINN.n384 VINN.n110 4.5005
R67629 VINN.n223 VINN.n110 4.5005
R67630 VINN.n386 VINN.n110 4.5005
R67631 VINN.n222 VINN.n110 4.5005
R67632 VINN.n388 VINN.n110 4.5005
R67633 VINN.n221 VINN.n110 4.5005
R67634 VINN.n390 VINN.n110 4.5005
R67635 VINN.n220 VINN.n110 4.5005
R67636 VINN.n392 VINN.n110 4.5005
R67637 VINN.n219 VINN.n110 4.5005
R67638 VINN.n394 VINN.n110 4.5005
R67639 VINN.n218 VINN.n110 4.5005
R67640 VINN.n396 VINN.n110 4.5005
R67641 VINN.n217 VINN.n110 4.5005
R67642 VINN.n398 VINN.n110 4.5005
R67643 VINN.n216 VINN.n110 4.5005
R67644 VINN.n400 VINN.n110 4.5005
R67645 VINN.n215 VINN.n110 4.5005
R67646 VINN.n654 VINN.n110 4.5005
R67647 VINN.n656 VINN.n110 4.5005
R67648 VINN.n110 VINN.n0 4.5005
R67649 VINN.n278 VINN.n191 4.5005
R67650 VINN.n276 VINN.n191 4.5005
R67651 VINN.n280 VINN.n191 4.5005
R67652 VINN.n275 VINN.n191 4.5005
R67653 VINN.n282 VINN.n191 4.5005
R67654 VINN.n274 VINN.n191 4.5005
R67655 VINN.n284 VINN.n191 4.5005
R67656 VINN.n273 VINN.n191 4.5005
R67657 VINN.n286 VINN.n191 4.5005
R67658 VINN.n272 VINN.n191 4.5005
R67659 VINN.n288 VINN.n191 4.5005
R67660 VINN.n271 VINN.n191 4.5005
R67661 VINN.n290 VINN.n191 4.5005
R67662 VINN.n270 VINN.n191 4.5005
R67663 VINN.n292 VINN.n191 4.5005
R67664 VINN.n269 VINN.n191 4.5005
R67665 VINN.n294 VINN.n191 4.5005
R67666 VINN.n268 VINN.n191 4.5005
R67667 VINN.n296 VINN.n191 4.5005
R67668 VINN.n267 VINN.n191 4.5005
R67669 VINN.n298 VINN.n191 4.5005
R67670 VINN.n266 VINN.n191 4.5005
R67671 VINN.n300 VINN.n191 4.5005
R67672 VINN.n265 VINN.n191 4.5005
R67673 VINN.n302 VINN.n191 4.5005
R67674 VINN.n264 VINN.n191 4.5005
R67675 VINN.n304 VINN.n191 4.5005
R67676 VINN.n263 VINN.n191 4.5005
R67677 VINN.n306 VINN.n191 4.5005
R67678 VINN.n262 VINN.n191 4.5005
R67679 VINN.n308 VINN.n191 4.5005
R67680 VINN.n261 VINN.n191 4.5005
R67681 VINN.n310 VINN.n191 4.5005
R67682 VINN.n260 VINN.n191 4.5005
R67683 VINN.n312 VINN.n191 4.5005
R67684 VINN.n259 VINN.n191 4.5005
R67685 VINN.n314 VINN.n191 4.5005
R67686 VINN.n258 VINN.n191 4.5005
R67687 VINN.n316 VINN.n191 4.5005
R67688 VINN.n257 VINN.n191 4.5005
R67689 VINN.n318 VINN.n191 4.5005
R67690 VINN.n256 VINN.n191 4.5005
R67691 VINN.n320 VINN.n191 4.5005
R67692 VINN.n255 VINN.n191 4.5005
R67693 VINN.n322 VINN.n191 4.5005
R67694 VINN.n254 VINN.n191 4.5005
R67695 VINN.n324 VINN.n191 4.5005
R67696 VINN.n253 VINN.n191 4.5005
R67697 VINN.n326 VINN.n191 4.5005
R67698 VINN.n252 VINN.n191 4.5005
R67699 VINN.n328 VINN.n191 4.5005
R67700 VINN.n251 VINN.n191 4.5005
R67701 VINN.n330 VINN.n191 4.5005
R67702 VINN.n250 VINN.n191 4.5005
R67703 VINN.n332 VINN.n191 4.5005
R67704 VINN.n249 VINN.n191 4.5005
R67705 VINN.n334 VINN.n191 4.5005
R67706 VINN.n248 VINN.n191 4.5005
R67707 VINN.n336 VINN.n191 4.5005
R67708 VINN.n247 VINN.n191 4.5005
R67709 VINN.n338 VINN.n191 4.5005
R67710 VINN.n246 VINN.n191 4.5005
R67711 VINN.n340 VINN.n191 4.5005
R67712 VINN.n245 VINN.n191 4.5005
R67713 VINN.n342 VINN.n191 4.5005
R67714 VINN.n244 VINN.n191 4.5005
R67715 VINN.n344 VINN.n191 4.5005
R67716 VINN.n243 VINN.n191 4.5005
R67717 VINN.n346 VINN.n191 4.5005
R67718 VINN.n242 VINN.n191 4.5005
R67719 VINN.n348 VINN.n191 4.5005
R67720 VINN.n241 VINN.n191 4.5005
R67721 VINN.n350 VINN.n191 4.5005
R67722 VINN.n240 VINN.n191 4.5005
R67723 VINN.n352 VINN.n191 4.5005
R67724 VINN.n239 VINN.n191 4.5005
R67725 VINN.n354 VINN.n191 4.5005
R67726 VINN.n238 VINN.n191 4.5005
R67727 VINN.n356 VINN.n191 4.5005
R67728 VINN.n237 VINN.n191 4.5005
R67729 VINN.n358 VINN.n191 4.5005
R67730 VINN.n236 VINN.n191 4.5005
R67731 VINN.n360 VINN.n191 4.5005
R67732 VINN.n235 VINN.n191 4.5005
R67733 VINN.n362 VINN.n191 4.5005
R67734 VINN.n234 VINN.n191 4.5005
R67735 VINN.n364 VINN.n191 4.5005
R67736 VINN.n233 VINN.n191 4.5005
R67737 VINN.n366 VINN.n191 4.5005
R67738 VINN.n232 VINN.n191 4.5005
R67739 VINN.n368 VINN.n191 4.5005
R67740 VINN.n231 VINN.n191 4.5005
R67741 VINN.n370 VINN.n191 4.5005
R67742 VINN.n230 VINN.n191 4.5005
R67743 VINN.n372 VINN.n191 4.5005
R67744 VINN.n229 VINN.n191 4.5005
R67745 VINN.n374 VINN.n191 4.5005
R67746 VINN.n228 VINN.n191 4.5005
R67747 VINN.n376 VINN.n191 4.5005
R67748 VINN.n227 VINN.n191 4.5005
R67749 VINN.n378 VINN.n191 4.5005
R67750 VINN.n226 VINN.n191 4.5005
R67751 VINN.n380 VINN.n191 4.5005
R67752 VINN.n225 VINN.n191 4.5005
R67753 VINN.n382 VINN.n191 4.5005
R67754 VINN.n224 VINN.n191 4.5005
R67755 VINN.n384 VINN.n191 4.5005
R67756 VINN.n223 VINN.n191 4.5005
R67757 VINN.n386 VINN.n191 4.5005
R67758 VINN.n222 VINN.n191 4.5005
R67759 VINN.n388 VINN.n191 4.5005
R67760 VINN.n221 VINN.n191 4.5005
R67761 VINN.n390 VINN.n191 4.5005
R67762 VINN.n220 VINN.n191 4.5005
R67763 VINN.n392 VINN.n191 4.5005
R67764 VINN.n219 VINN.n191 4.5005
R67765 VINN.n394 VINN.n191 4.5005
R67766 VINN.n218 VINN.n191 4.5005
R67767 VINN.n396 VINN.n191 4.5005
R67768 VINN.n217 VINN.n191 4.5005
R67769 VINN.n398 VINN.n191 4.5005
R67770 VINN.n216 VINN.n191 4.5005
R67771 VINN.n400 VINN.n191 4.5005
R67772 VINN.n215 VINN.n191 4.5005
R67773 VINN.n654 VINN.n191 4.5005
R67774 VINN.n656 VINN.n191 4.5005
R67775 VINN.n191 VINN.n0 4.5005
R67776 VINN.n278 VINN.n109 4.5005
R67777 VINN.n276 VINN.n109 4.5005
R67778 VINN.n280 VINN.n109 4.5005
R67779 VINN.n275 VINN.n109 4.5005
R67780 VINN.n282 VINN.n109 4.5005
R67781 VINN.n274 VINN.n109 4.5005
R67782 VINN.n284 VINN.n109 4.5005
R67783 VINN.n273 VINN.n109 4.5005
R67784 VINN.n286 VINN.n109 4.5005
R67785 VINN.n272 VINN.n109 4.5005
R67786 VINN.n288 VINN.n109 4.5005
R67787 VINN.n271 VINN.n109 4.5005
R67788 VINN.n290 VINN.n109 4.5005
R67789 VINN.n270 VINN.n109 4.5005
R67790 VINN.n292 VINN.n109 4.5005
R67791 VINN.n269 VINN.n109 4.5005
R67792 VINN.n294 VINN.n109 4.5005
R67793 VINN.n268 VINN.n109 4.5005
R67794 VINN.n296 VINN.n109 4.5005
R67795 VINN.n267 VINN.n109 4.5005
R67796 VINN.n298 VINN.n109 4.5005
R67797 VINN.n266 VINN.n109 4.5005
R67798 VINN.n300 VINN.n109 4.5005
R67799 VINN.n265 VINN.n109 4.5005
R67800 VINN.n302 VINN.n109 4.5005
R67801 VINN.n264 VINN.n109 4.5005
R67802 VINN.n304 VINN.n109 4.5005
R67803 VINN.n263 VINN.n109 4.5005
R67804 VINN.n306 VINN.n109 4.5005
R67805 VINN.n262 VINN.n109 4.5005
R67806 VINN.n308 VINN.n109 4.5005
R67807 VINN.n261 VINN.n109 4.5005
R67808 VINN.n310 VINN.n109 4.5005
R67809 VINN.n260 VINN.n109 4.5005
R67810 VINN.n312 VINN.n109 4.5005
R67811 VINN.n259 VINN.n109 4.5005
R67812 VINN.n314 VINN.n109 4.5005
R67813 VINN.n258 VINN.n109 4.5005
R67814 VINN.n316 VINN.n109 4.5005
R67815 VINN.n257 VINN.n109 4.5005
R67816 VINN.n318 VINN.n109 4.5005
R67817 VINN.n256 VINN.n109 4.5005
R67818 VINN.n320 VINN.n109 4.5005
R67819 VINN.n255 VINN.n109 4.5005
R67820 VINN.n322 VINN.n109 4.5005
R67821 VINN.n254 VINN.n109 4.5005
R67822 VINN.n324 VINN.n109 4.5005
R67823 VINN.n253 VINN.n109 4.5005
R67824 VINN.n326 VINN.n109 4.5005
R67825 VINN.n252 VINN.n109 4.5005
R67826 VINN.n328 VINN.n109 4.5005
R67827 VINN.n251 VINN.n109 4.5005
R67828 VINN.n330 VINN.n109 4.5005
R67829 VINN.n250 VINN.n109 4.5005
R67830 VINN.n332 VINN.n109 4.5005
R67831 VINN.n249 VINN.n109 4.5005
R67832 VINN.n334 VINN.n109 4.5005
R67833 VINN.n248 VINN.n109 4.5005
R67834 VINN.n336 VINN.n109 4.5005
R67835 VINN.n247 VINN.n109 4.5005
R67836 VINN.n338 VINN.n109 4.5005
R67837 VINN.n246 VINN.n109 4.5005
R67838 VINN.n340 VINN.n109 4.5005
R67839 VINN.n245 VINN.n109 4.5005
R67840 VINN.n342 VINN.n109 4.5005
R67841 VINN.n244 VINN.n109 4.5005
R67842 VINN.n344 VINN.n109 4.5005
R67843 VINN.n243 VINN.n109 4.5005
R67844 VINN.n346 VINN.n109 4.5005
R67845 VINN.n242 VINN.n109 4.5005
R67846 VINN.n348 VINN.n109 4.5005
R67847 VINN.n241 VINN.n109 4.5005
R67848 VINN.n350 VINN.n109 4.5005
R67849 VINN.n240 VINN.n109 4.5005
R67850 VINN.n352 VINN.n109 4.5005
R67851 VINN.n239 VINN.n109 4.5005
R67852 VINN.n354 VINN.n109 4.5005
R67853 VINN.n238 VINN.n109 4.5005
R67854 VINN.n356 VINN.n109 4.5005
R67855 VINN.n237 VINN.n109 4.5005
R67856 VINN.n358 VINN.n109 4.5005
R67857 VINN.n236 VINN.n109 4.5005
R67858 VINN.n360 VINN.n109 4.5005
R67859 VINN.n235 VINN.n109 4.5005
R67860 VINN.n362 VINN.n109 4.5005
R67861 VINN.n234 VINN.n109 4.5005
R67862 VINN.n364 VINN.n109 4.5005
R67863 VINN.n233 VINN.n109 4.5005
R67864 VINN.n366 VINN.n109 4.5005
R67865 VINN.n232 VINN.n109 4.5005
R67866 VINN.n368 VINN.n109 4.5005
R67867 VINN.n231 VINN.n109 4.5005
R67868 VINN.n370 VINN.n109 4.5005
R67869 VINN.n230 VINN.n109 4.5005
R67870 VINN.n372 VINN.n109 4.5005
R67871 VINN.n229 VINN.n109 4.5005
R67872 VINN.n374 VINN.n109 4.5005
R67873 VINN.n228 VINN.n109 4.5005
R67874 VINN.n376 VINN.n109 4.5005
R67875 VINN.n227 VINN.n109 4.5005
R67876 VINN.n378 VINN.n109 4.5005
R67877 VINN.n226 VINN.n109 4.5005
R67878 VINN.n380 VINN.n109 4.5005
R67879 VINN.n225 VINN.n109 4.5005
R67880 VINN.n382 VINN.n109 4.5005
R67881 VINN.n224 VINN.n109 4.5005
R67882 VINN.n384 VINN.n109 4.5005
R67883 VINN.n223 VINN.n109 4.5005
R67884 VINN.n386 VINN.n109 4.5005
R67885 VINN.n222 VINN.n109 4.5005
R67886 VINN.n388 VINN.n109 4.5005
R67887 VINN.n221 VINN.n109 4.5005
R67888 VINN.n390 VINN.n109 4.5005
R67889 VINN.n220 VINN.n109 4.5005
R67890 VINN.n392 VINN.n109 4.5005
R67891 VINN.n219 VINN.n109 4.5005
R67892 VINN.n394 VINN.n109 4.5005
R67893 VINN.n218 VINN.n109 4.5005
R67894 VINN.n396 VINN.n109 4.5005
R67895 VINN.n217 VINN.n109 4.5005
R67896 VINN.n398 VINN.n109 4.5005
R67897 VINN.n216 VINN.n109 4.5005
R67898 VINN.n400 VINN.n109 4.5005
R67899 VINN.n215 VINN.n109 4.5005
R67900 VINN.n654 VINN.n109 4.5005
R67901 VINN.n656 VINN.n109 4.5005
R67902 VINN.n109 VINN.n0 4.5005
R67903 VINN.n278 VINN.n192 4.5005
R67904 VINN.n276 VINN.n192 4.5005
R67905 VINN.n280 VINN.n192 4.5005
R67906 VINN.n275 VINN.n192 4.5005
R67907 VINN.n282 VINN.n192 4.5005
R67908 VINN.n274 VINN.n192 4.5005
R67909 VINN.n284 VINN.n192 4.5005
R67910 VINN.n273 VINN.n192 4.5005
R67911 VINN.n286 VINN.n192 4.5005
R67912 VINN.n272 VINN.n192 4.5005
R67913 VINN.n288 VINN.n192 4.5005
R67914 VINN.n271 VINN.n192 4.5005
R67915 VINN.n290 VINN.n192 4.5005
R67916 VINN.n270 VINN.n192 4.5005
R67917 VINN.n292 VINN.n192 4.5005
R67918 VINN.n269 VINN.n192 4.5005
R67919 VINN.n294 VINN.n192 4.5005
R67920 VINN.n268 VINN.n192 4.5005
R67921 VINN.n296 VINN.n192 4.5005
R67922 VINN.n267 VINN.n192 4.5005
R67923 VINN.n298 VINN.n192 4.5005
R67924 VINN.n266 VINN.n192 4.5005
R67925 VINN.n300 VINN.n192 4.5005
R67926 VINN.n265 VINN.n192 4.5005
R67927 VINN.n302 VINN.n192 4.5005
R67928 VINN.n264 VINN.n192 4.5005
R67929 VINN.n304 VINN.n192 4.5005
R67930 VINN.n263 VINN.n192 4.5005
R67931 VINN.n306 VINN.n192 4.5005
R67932 VINN.n262 VINN.n192 4.5005
R67933 VINN.n308 VINN.n192 4.5005
R67934 VINN.n261 VINN.n192 4.5005
R67935 VINN.n310 VINN.n192 4.5005
R67936 VINN.n260 VINN.n192 4.5005
R67937 VINN.n312 VINN.n192 4.5005
R67938 VINN.n259 VINN.n192 4.5005
R67939 VINN.n314 VINN.n192 4.5005
R67940 VINN.n258 VINN.n192 4.5005
R67941 VINN.n316 VINN.n192 4.5005
R67942 VINN.n257 VINN.n192 4.5005
R67943 VINN.n318 VINN.n192 4.5005
R67944 VINN.n256 VINN.n192 4.5005
R67945 VINN.n320 VINN.n192 4.5005
R67946 VINN.n255 VINN.n192 4.5005
R67947 VINN.n322 VINN.n192 4.5005
R67948 VINN.n254 VINN.n192 4.5005
R67949 VINN.n324 VINN.n192 4.5005
R67950 VINN.n253 VINN.n192 4.5005
R67951 VINN.n326 VINN.n192 4.5005
R67952 VINN.n252 VINN.n192 4.5005
R67953 VINN.n328 VINN.n192 4.5005
R67954 VINN.n251 VINN.n192 4.5005
R67955 VINN.n330 VINN.n192 4.5005
R67956 VINN.n250 VINN.n192 4.5005
R67957 VINN.n332 VINN.n192 4.5005
R67958 VINN.n249 VINN.n192 4.5005
R67959 VINN.n334 VINN.n192 4.5005
R67960 VINN.n248 VINN.n192 4.5005
R67961 VINN.n336 VINN.n192 4.5005
R67962 VINN.n247 VINN.n192 4.5005
R67963 VINN.n338 VINN.n192 4.5005
R67964 VINN.n246 VINN.n192 4.5005
R67965 VINN.n340 VINN.n192 4.5005
R67966 VINN.n245 VINN.n192 4.5005
R67967 VINN.n342 VINN.n192 4.5005
R67968 VINN.n244 VINN.n192 4.5005
R67969 VINN.n344 VINN.n192 4.5005
R67970 VINN.n243 VINN.n192 4.5005
R67971 VINN.n346 VINN.n192 4.5005
R67972 VINN.n242 VINN.n192 4.5005
R67973 VINN.n348 VINN.n192 4.5005
R67974 VINN.n241 VINN.n192 4.5005
R67975 VINN.n350 VINN.n192 4.5005
R67976 VINN.n240 VINN.n192 4.5005
R67977 VINN.n352 VINN.n192 4.5005
R67978 VINN.n239 VINN.n192 4.5005
R67979 VINN.n354 VINN.n192 4.5005
R67980 VINN.n238 VINN.n192 4.5005
R67981 VINN.n356 VINN.n192 4.5005
R67982 VINN.n237 VINN.n192 4.5005
R67983 VINN.n358 VINN.n192 4.5005
R67984 VINN.n236 VINN.n192 4.5005
R67985 VINN.n360 VINN.n192 4.5005
R67986 VINN.n235 VINN.n192 4.5005
R67987 VINN.n362 VINN.n192 4.5005
R67988 VINN.n234 VINN.n192 4.5005
R67989 VINN.n364 VINN.n192 4.5005
R67990 VINN.n233 VINN.n192 4.5005
R67991 VINN.n366 VINN.n192 4.5005
R67992 VINN.n232 VINN.n192 4.5005
R67993 VINN.n368 VINN.n192 4.5005
R67994 VINN.n231 VINN.n192 4.5005
R67995 VINN.n370 VINN.n192 4.5005
R67996 VINN.n230 VINN.n192 4.5005
R67997 VINN.n372 VINN.n192 4.5005
R67998 VINN.n229 VINN.n192 4.5005
R67999 VINN.n374 VINN.n192 4.5005
R68000 VINN.n228 VINN.n192 4.5005
R68001 VINN.n376 VINN.n192 4.5005
R68002 VINN.n227 VINN.n192 4.5005
R68003 VINN.n378 VINN.n192 4.5005
R68004 VINN.n226 VINN.n192 4.5005
R68005 VINN.n380 VINN.n192 4.5005
R68006 VINN.n225 VINN.n192 4.5005
R68007 VINN.n382 VINN.n192 4.5005
R68008 VINN.n224 VINN.n192 4.5005
R68009 VINN.n384 VINN.n192 4.5005
R68010 VINN.n223 VINN.n192 4.5005
R68011 VINN.n386 VINN.n192 4.5005
R68012 VINN.n222 VINN.n192 4.5005
R68013 VINN.n388 VINN.n192 4.5005
R68014 VINN.n221 VINN.n192 4.5005
R68015 VINN.n390 VINN.n192 4.5005
R68016 VINN.n220 VINN.n192 4.5005
R68017 VINN.n392 VINN.n192 4.5005
R68018 VINN.n219 VINN.n192 4.5005
R68019 VINN.n394 VINN.n192 4.5005
R68020 VINN.n218 VINN.n192 4.5005
R68021 VINN.n396 VINN.n192 4.5005
R68022 VINN.n217 VINN.n192 4.5005
R68023 VINN.n398 VINN.n192 4.5005
R68024 VINN.n216 VINN.n192 4.5005
R68025 VINN.n400 VINN.n192 4.5005
R68026 VINN.n215 VINN.n192 4.5005
R68027 VINN.n654 VINN.n192 4.5005
R68028 VINN.n656 VINN.n192 4.5005
R68029 VINN.n192 VINN.n0 4.5005
R68030 VINN.n278 VINN.n108 4.5005
R68031 VINN.n276 VINN.n108 4.5005
R68032 VINN.n280 VINN.n108 4.5005
R68033 VINN.n275 VINN.n108 4.5005
R68034 VINN.n282 VINN.n108 4.5005
R68035 VINN.n274 VINN.n108 4.5005
R68036 VINN.n284 VINN.n108 4.5005
R68037 VINN.n273 VINN.n108 4.5005
R68038 VINN.n286 VINN.n108 4.5005
R68039 VINN.n272 VINN.n108 4.5005
R68040 VINN.n288 VINN.n108 4.5005
R68041 VINN.n271 VINN.n108 4.5005
R68042 VINN.n290 VINN.n108 4.5005
R68043 VINN.n270 VINN.n108 4.5005
R68044 VINN.n292 VINN.n108 4.5005
R68045 VINN.n269 VINN.n108 4.5005
R68046 VINN.n294 VINN.n108 4.5005
R68047 VINN.n268 VINN.n108 4.5005
R68048 VINN.n296 VINN.n108 4.5005
R68049 VINN.n267 VINN.n108 4.5005
R68050 VINN.n298 VINN.n108 4.5005
R68051 VINN.n266 VINN.n108 4.5005
R68052 VINN.n300 VINN.n108 4.5005
R68053 VINN.n265 VINN.n108 4.5005
R68054 VINN.n302 VINN.n108 4.5005
R68055 VINN.n264 VINN.n108 4.5005
R68056 VINN.n304 VINN.n108 4.5005
R68057 VINN.n263 VINN.n108 4.5005
R68058 VINN.n306 VINN.n108 4.5005
R68059 VINN.n262 VINN.n108 4.5005
R68060 VINN.n308 VINN.n108 4.5005
R68061 VINN.n261 VINN.n108 4.5005
R68062 VINN.n310 VINN.n108 4.5005
R68063 VINN.n260 VINN.n108 4.5005
R68064 VINN.n312 VINN.n108 4.5005
R68065 VINN.n259 VINN.n108 4.5005
R68066 VINN.n314 VINN.n108 4.5005
R68067 VINN.n258 VINN.n108 4.5005
R68068 VINN.n316 VINN.n108 4.5005
R68069 VINN.n257 VINN.n108 4.5005
R68070 VINN.n318 VINN.n108 4.5005
R68071 VINN.n256 VINN.n108 4.5005
R68072 VINN.n320 VINN.n108 4.5005
R68073 VINN.n255 VINN.n108 4.5005
R68074 VINN.n322 VINN.n108 4.5005
R68075 VINN.n254 VINN.n108 4.5005
R68076 VINN.n324 VINN.n108 4.5005
R68077 VINN.n253 VINN.n108 4.5005
R68078 VINN.n326 VINN.n108 4.5005
R68079 VINN.n252 VINN.n108 4.5005
R68080 VINN.n328 VINN.n108 4.5005
R68081 VINN.n251 VINN.n108 4.5005
R68082 VINN.n330 VINN.n108 4.5005
R68083 VINN.n250 VINN.n108 4.5005
R68084 VINN.n332 VINN.n108 4.5005
R68085 VINN.n249 VINN.n108 4.5005
R68086 VINN.n334 VINN.n108 4.5005
R68087 VINN.n248 VINN.n108 4.5005
R68088 VINN.n336 VINN.n108 4.5005
R68089 VINN.n247 VINN.n108 4.5005
R68090 VINN.n338 VINN.n108 4.5005
R68091 VINN.n246 VINN.n108 4.5005
R68092 VINN.n340 VINN.n108 4.5005
R68093 VINN.n245 VINN.n108 4.5005
R68094 VINN.n342 VINN.n108 4.5005
R68095 VINN.n244 VINN.n108 4.5005
R68096 VINN.n344 VINN.n108 4.5005
R68097 VINN.n243 VINN.n108 4.5005
R68098 VINN.n346 VINN.n108 4.5005
R68099 VINN.n242 VINN.n108 4.5005
R68100 VINN.n348 VINN.n108 4.5005
R68101 VINN.n241 VINN.n108 4.5005
R68102 VINN.n350 VINN.n108 4.5005
R68103 VINN.n240 VINN.n108 4.5005
R68104 VINN.n352 VINN.n108 4.5005
R68105 VINN.n239 VINN.n108 4.5005
R68106 VINN.n354 VINN.n108 4.5005
R68107 VINN.n238 VINN.n108 4.5005
R68108 VINN.n356 VINN.n108 4.5005
R68109 VINN.n237 VINN.n108 4.5005
R68110 VINN.n358 VINN.n108 4.5005
R68111 VINN.n236 VINN.n108 4.5005
R68112 VINN.n360 VINN.n108 4.5005
R68113 VINN.n235 VINN.n108 4.5005
R68114 VINN.n362 VINN.n108 4.5005
R68115 VINN.n234 VINN.n108 4.5005
R68116 VINN.n364 VINN.n108 4.5005
R68117 VINN.n233 VINN.n108 4.5005
R68118 VINN.n366 VINN.n108 4.5005
R68119 VINN.n232 VINN.n108 4.5005
R68120 VINN.n368 VINN.n108 4.5005
R68121 VINN.n231 VINN.n108 4.5005
R68122 VINN.n370 VINN.n108 4.5005
R68123 VINN.n230 VINN.n108 4.5005
R68124 VINN.n372 VINN.n108 4.5005
R68125 VINN.n229 VINN.n108 4.5005
R68126 VINN.n374 VINN.n108 4.5005
R68127 VINN.n228 VINN.n108 4.5005
R68128 VINN.n376 VINN.n108 4.5005
R68129 VINN.n227 VINN.n108 4.5005
R68130 VINN.n378 VINN.n108 4.5005
R68131 VINN.n226 VINN.n108 4.5005
R68132 VINN.n380 VINN.n108 4.5005
R68133 VINN.n225 VINN.n108 4.5005
R68134 VINN.n382 VINN.n108 4.5005
R68135 VINN.n224 VINN.n108 4.5005
R68136 VINN.n384 VINN.n108 4.5005
R68137 VINN.n223 VINN.n108 4.5005
R68138 VINN.n386 VINN.n108 4.5005
R68139 VINN.n222 VINN.n108 4.5005
R68140 VINN.n388 VINN.n108 4.5005
R68141 VINN.n221 VINN.n108 4.5005
R68142 VINN.n390 VINN.n108 4.5005
R68143 VINN.n220 VINN.n108 4.5005
R68144 VINN.n392 VINN.n108 4.5005
R68145 VINN.n219 VINN.n108 4.5005
R68146 VINN.n394 VINN.n108 4.5005
R68147 VINN.n218 VINN.n108 4.5005
R68148 VINN.n396 VINN.n108 4.5005
R68149 VINN.n217 VINN.n108 4.5005
R68150 VINN.n398 VINN.n108 4.5005
R68151 VINN.n216 VINN.n108 4.5005
R68152 VINN.n400 VINN.n108 4.5005
R68153 VINN.n215 VINN.n108 4.5005
R68154 VINN.n654 VINN.n108 4.5005
R68155 VINN.n656 VINN.n108 4.5005
R68156 VINN.n108 VINN.n0 4.5005
R68157 VINN.n278 VINN.n193 4.5005
R68158 VINN.n276 VINN.n193 4.5005
R68159 VINN.n280 VINN.n193 4.5005
R68160 VINN.n275 VINN.n193 4.5005
R68161 VINN.n282 VINN.n193 4.5005
R68162 VINN.n274 VINN.n193 4.5005
R68163 VINN.n284 VINN.n193 4.5005
R68164 VINN.n273 VINN.n193 4.5005
R68165 VINN.n286 VINN.n193 4.5005
R68166 VINN.n272 VINN.n193 4.5005
R68167 VINN.n288 VINN.n193 4.5005
R68168 VINN.n271 VINN.n193 4.5005
R68169 VINN.n290 VINN.n193 4.5005
R68170 VINN.n270 VINN.n193 4.5005
R68171 VINN.n292 VINN.n193 4.5005
R68172 VINN.n269 VINN.n193 4.5005
R68173 VINN.n294 VINN.n193 4.5005
R68174 VINN.n268 VINN.n193 4.5005
R68175 VINN.n296 VINN.n193 4.5005
R68176 VINN.n267 VINN.n193 4.5005
R68177 VINN.n298 VINN.n193 4.5005
R68178 VINN.n266 VINN.n193 4.5005
R68179 VINN.n300 VINN.n193 4.5005
R68180 VINN.n265 VINN.n193 4.5005
R68181 VINN.n302 VINN.n193 4.5005
R68182 VINN.n264 VINN.n193 4.5005
R68183 VINN.n304 VINN.n193 4.5005
R68184 VINN.n263 VINN.n193 4.5005
R68185 VINN.n306 VINN.n193 4.5005
R68186 VINN.n262 VINN.n193 4.5005
R68187 VINN.n308 VINN.n193 4.5005
R68188 VINN.n261 VINN.n193 4.5005
R68189 VINN.n310 VINN.n193 4.5005
R68190 VINN.n260 VINN.n193 4.5005
R68191 VINN.n312 VINN.n193 4.5005
R68192 VINN.n259 VINN.n193 4.5005
R68193 VINN.n314 VINN.n193 4.5005
R68194 VINN.n258 VINN.n193 4.5005
R68195 VINN.n316 VINN.n193 4.5005
R68196 VINN.n257 VINN.n193 4.5005
R68197 VINN.n318 VINN.n193 4.5005
R68198 VINN.n256 VINN.n193 4.5005
R68199 VINN.n320 VINN.n193 4.5005
R68200 VINN.n255 VINN.n193 4.5005
R68201 VINN.n322 VINN.n193 4.5005
R68202 VINN.n254 VINN.n193 4.5005
R68203 VINN.n324 VINN.n193 4.5005
R68204 VINN.n253 VINN.n193 4.5005
R68205 VINN.n326 VINN.n193 4.5005
R68206 VINN.n252 VINN.n193 4.5005
R68207 VINN.n328 VINN.n193 4.5005
R68208 VINN.n251 VINN.n193 4.5005
R68209 VINN.n330 VINN.n193 4.5005
R68210 VINN.n250 VINN.n193 4.5005
R68211 VINN.n332 VINN.n193 4.5005
R68212 VINN.n249 VINN.n193 4.5005
R68213 VINN.n334 VINN.n193 4.5005
R68214 VINN.n248 VINN.n193 4.5005
R68215 VINN.n336 VINN.n193 4.5005
R68216 VINN.n247 VINN.n193 4.5005
R68217 VINN.n338 VINN.n193 4.5005
R68218 VINN.n246 VINN.n193 4.5005
R68219 VINN.n340 VINN.n193 4.5005
R68220 VINN.n245 VINN.n193 4.5005
R68221 VINN.n342 VINN.n193 4.5005
R68222 VINN.n244 VINN.n193 4.5005
R68223 VINN.n344 VINN.n193 4.5005
R68224 VINN.n243 VINN.n193 4.5005
R68225 VINN.n346 VINN.n193 4.5005
R68226 VINN.n242 VINN.n193 4.5005
R68227 VINN.n348 VINN.n193 4.5005
R68228 VINN.n241 VINN.n193 4.5005
R68229 VINN.n350 VINN.n193 4.5005
R68230 VINN.n240 VINN.n193 4.5005
R68231 VINN.n352 VINN.n193 4.5005
R68232 VINN.n239 VINN.n193 4.5005
R68233 VINN.n354 VINN.n193 4.5005
R68234 VINN.n238 VINN.n193 4.5005
R68235 VINN.n356 VINN.n193 4.5005
R68236 VINN.n237 VINN.n193 4.5005
R68237 VINN.n358 VINN.n193 4.5005
R68238 VINN.n236 VINN.n193 4.5005
R68239 VINN.n360 VINN.n193 4.5005
R68240 VINN.n235 VINN.n193 4.5005
R68241 VINN.n362 VINN.n193 4.5005
R68242 VINN.n234 VINN.n193 4.5005
R68243 VINN.n364 VINN.n193 4.5005
R68244 VINN.n233 VINN.n193 4.5005
R68245 VINN.n366 VINN.n193 4.5005
R68246 VINN.n232 VINN.n193 4.5005
R68247 VINN.n368 VINN.n193 4.5005
R68248 VINN.n231 VINN.n193 4.5005
R68249 VINN.n370 VINN.n193 4.5005
R68250 VINN.n230 VINN.n193 4.5005
R68251 VINN.n372 VINN.n193 4.5005
R68252 VINN.n229 VINN.n193 4.5005
R68253 VINN.n374 VINN.n193 4.5005
R68254 VINN.n228 VINN.n193 4.5005
R68255 VINN.n376 VINN.n193 4.5005
R68256 VINN.n227 VINN.n193 4.5005
R68257 VINN.n378 VINN.n193 4.5005
R68258 VINN.n226 VINN.n193 4.5005
R68259 VINN.n380 VINN.n193 4.5005
R68260 VINN.n225 VINN.n193 4.5005
R68261 VINN.n382 VINN.n193 4.5005
R68262 VINN.n224 VINN.n193 4.5005
R68263 VINN.n384 VINN.n193 4.5005
R68264 VINN.n223 VINN.n193 4.5005
R68265 VINN.n386 VINN.n193 4.5005
R68266 VINN.n222 VINN.n193 4.5005
R68267 VINN.n388 VINN.n193 4.5005
R68268 VINN.n221 VINN.n193 4.5005
R68269 VINN.n390 VINN.n193 4.5005
R68270 VINN.n220 VINN.n193 4.5005
R68271 VINN.n392 VINN.n193 4.5005
R68272 VINN.n219 VINN.n193 4.5005
R68273 VINN.n394 VINN.n193 4.5005
R68274 VINN.n218 VINN.n193 4.5005
R68275 VINN.n396 VINN.n193 4.5005
R68276 VINN.n217 VINN.n193 4.5005
R68277 VINN.n398 VINN.n193 4.5005
R68278 VINN.n216 VINN.n193 4.5005
R68279 VINN.n400 VINN.n193 4.5005
R68280 VINN.n215 VINN.n193 4.5005
R68281 VINN.n654 VINN.n193 4.5005
R68282 VINN.n656 VINN.n193 4.5005
R68283 VINN.n193 VINN.n0 4.5005
R68284 VINN.n278 VINN.n107 4.5005
R68285 VINN.n276 VINN.n107 4.5005
R68286 VINN.n280 VINN.n107 4.5005
R68287 VINN.n275 VINN.n107 4.5005
R68288 VINN.n282 VINN.n107 4.5005
R68289 VINN.n274 VINN.n107 4.5005
R68290 VINN.n284 VINN.n107 4.5005
R68291 VINN.n273 VINN.n107 4.5005
R68292 VINN.n286 VINN.n107 4.5005
R68293 VINN.n272 VINN.n107 4.5005
R68294 VINN.n288 VINN.n107 4.5005
R68295 VINN.n271 VINN.n107 4.5005
R68296 VINN.n290 VINN.n107 4.5005
R68297 VINN.n270 VINN.n107 4.5005
R68298 VINN.n292 VINN.n107 4.5005
R68299 VINN.n269 VINN.n107 4.5005
R68300 VINN.n294 VINN.n107 4.5005
R68301 VINN.n268 VINN.n107 4.5005
R68302 VINN.n296 VINN.n107 4.5005
R68303 VINN.n267 VINN.n107 4.5005
R68304 VINN.n298 VINN.n107 4.5005
R68305 VINN.n266 VINN.n107 4.5005
R68306 VINN.n300 VINN.n107 4.5005
R68307 VINN.n265 VINN.n107 4.5005
R68308 VINN.n302 VINN.n107 4.5005
R68309 VINN.n264 VINN.n107 4.5005
R68310 VINN.n304 VINN.n107 4.5005
R68311 VINN.n263 VINN.n107 4.5005
R68312 VINN.n306 VINN.n107 4.5005
R68313 VINN.n262 VINN.n107 4.5005
R68314 VINN.n308 VINN.n107 4.5005
R68315 VINN.n261 VINN.n107 4.5005
R68316 VINN.n310 VINN.n107 4.5005
R68317 VINN.n260 VINN.n107 4.5005
R68318 VINN.n312 VINN.n107 4.5005
R68319 VINN.n259 VINN.n107 4.5005
R68320 VINN.n314 VINN.n107 4.5005
R68321 VINN.n258 VINN.n107 4.5005
R68322 VINN.n316 VINN.n107 4.5005
R68323 VINN.n257 VINN.n107 4.5005
R68324 VINN.n318 VINN.n107 4.5005
R68325 VINN.n256 VINN.n107 4.5005
R68326 VINN.n320 VINN.n107 4.5005
R68327 VINN.n255 VINN.n107 4.5005
R68328 VINN.n322 VINN.n107 4.5005
R68329 VINN.n254 VINN.n107 4.5005
R68330 VINN.n324 VINN.n107 4.5005
R68331 VINN.n253 VINN.n107 4.5005
R68332 VINN.n326 VINN.n107 4.5005
R68333 VINN.n252 VINN.n107 4.5005
R68334 VINN.n328 VINN.n107 4.5005
R68335 VINN.n251 VINN.n107 4.5005
R68336 VINN.n330 VINN.n107 4.5005
R68337 VINN.n250 VINN.n107 4.5005
R68338 VINN.n332 VINN.n107 4.5005
R68339 VINN.n249 VINN.n107 4.5005
R68340 VINN.n334 VINN.n107 4.5005
R68341 VINN.n248 VINN.n107 4.5005
R68342 VINN.n336 VINN.n107 4.5005
R68343 VINN.n247 VINN.n107 4.5005
R68344 VINN.n338 VINN.n107 4.5005
R68345 VINN.n246 VINN.n107 4.5005
R68346 VINN.n340 VINN.n107 4.5005
R68347 VINN.n245 VINN.n107 4.5005
R68348 VINN.n342 VINN.n107 4.5005
R68349 VINN.n244 VINN.n107 4.5005
R68350 VINN.n344 VINN.n107 4.5005
R68351 VINN.n243 VINN.n107 4.5005
R68352 VINN.n346 VINN.n107 4.5005
R68353 VINN.n242 VINN.n107 4.5005
R68354 VINN.n348 VINN.n107 4.5005
R68355 VINN.n241 VINN.n107 4.5005
R68356 VINN.n350 VINN.n107 4.5005
R68357 VINN.n240 VINN.n107 4.5005
R68358 VINN.n352 VINN.n107 4.5005
R68359 VINN.n239 VINN.n107 4.5005
R68360 VINN.n354 VINN.n107 4.5005
R68361 VINN.n238 VINN.n107 4.5005
R68362 VINN.n356 VINN.n107 4.5005
R68363 VINN.n237 VINN.n107 4.5005
R68364 VINN.n358 VINN.n107 4.5005
R68365 VINN.n236 VINN.n107 4.5005
R68366 VINN.n360 VINN.n107 4.5005
R68367 VINN.n235 VINN.n107 4.5005
R68368 VINN.n362 VINN.n107 4.5005
R68369 VINN.n234 VINN.n107 4.5005
R68370 VINN.n364 VINN.n107 4.5005
R68371 VINN.n233 VINN.n107 4.5005
R68372 VINN.n366 VINN.n107 4.5005
R68373 VINN.n232 VINN.n107 4.5005
R68374 VINN.n368 VINN.n107 4.5005
R68375 VINN.n231 VINN.n107 4.5005
R68376 VINN.n370 VINN.n107 4.5005
R68377 VINN.n230 VINN.n107 4.5005
R68378 VINN.n372 VINN.n107 4.5005
R68379 VINN.n229 VINN.n107 4.5005
R68380 VINN.n374 VINN.n107 4.5005
R68381 VINN.n228 VINN.n107 4.5005
R68382 VINN.n376 VINN.n107 4.5005
R68383 VINN.n227 VINN.n107 4.5005
R68384 VINN.n378 VINN.n107 4.5005
R68385 VINN.n226 VINN.n107 4.5005
R68386 VINN.n380 VINN.n107 4.5005
R68387 VINN.n225 VINN.n107 4.5005
R68388 VINN.n382 VINN.n107 4.5005
R68389 VINN.n224 VINN.n107 4.5005
R68390 VINN.n384 VINN.n107 4.5005
R68391 VINN.n223 VINN.n107 4.5005
R68392 VINN.n386 VINN.n107 4.5005
R68393 VINN.n222 VINN.n107 4.5005
R68394 VINN.n388 VINN.n107 4.5005
R68395 VINN.n221 VINN.n107 4.5005
R68396 VINN.n390 VINN.n107 4.5005
R68397 VINN.n220 VINN.n107 4.5005
R68398 VINN.n392 VINN.n107 4.5005
R68399 VINN.n219 VINN.n107 4.5005
R68400 VINN.n394 VINN.n107 4.5005
R68401 VINN.n218 VINN.n107 4.5005
R68402 VINN.n396 VINN.n107 4.5005
R68403 VINN.n217 VINN.n107 4.5005
R68404 VINN.n398 VINN.n107 4.5005
R68405 VINN.n216 VINN.n107 4.5005
R68406 VINN.n400 VINN.n107 4.5005
R68407 VINN.n215 VINN.n107 4.5005
R68408 VINN.n654 VINN.n107 4.5005
R68409 VINN.n656 VINN.n107 4.5005
R68410 VINN.n107 VINN.n0 4.5005
R68411 VINN.n278 VINN.n194 4.5005
R68412 VINN.n276 VINN.n194 4.5005
R68413 VINN.n280 VINN.n194 4.5005
R68414 VINN.n275 VINN.n194 4.5005
R68415 VINN.n282 VINN.n194 4.5005
R68416 VINN.n274 VINN.n194 4.5005
R68417 VINN.n284 VINN.n194 4.5005
R68418 VINN.n273 VINN.n194 4.5005
R68419 VINN.n286 VINN.n194 4.5005
R68420 VINN.n272 VINN.n194 4.5005
R68421 VINN.n288 VINN.n194 4.5005
R68422 VINN.n271 VINN.n194 4.5005
R68423 VINN.n290 VINN.n194 4.5005
R68424 VINN.n270 VINN.n194 4.5005
R68425 VINN.n292 VINN.n194 4.5005
R68426 VINN.n269 VINN.n194 4.5005
R68427 VINN.n294 VINN.n194 4.5005
R68428 VINN.n268 VINN.n194 4.5005
R68429 VINN.n296 VINN.n194 4.5005
R68430 VINN.n267 VINN.n194 4.5005
R68431 VINN.n298 VINN.n194 4.5005
R68432 VINN.n266 VINN.n194 4.5005
R68433 VINN.n300 VINN.n194 4.5005
R68434 VINN.n265 VINN.n194 4.5005
R68435 VINN.n302 VINN.n194 4.5005
R68436 VINN.n264 VINN.n194 4.5005
R68437 VINN.n304 VINN.n194 4.5005
R68438 VINN.n263 VINN.n194 4.5005
R68439 VINN.n306 VINN.n194 4.5005
R68440 VINN.n262 VINN.n194 4.5005
R68441 VINN.n308 VINN.n194 4.5005
R68442 VINN.n261 VINN.n194 4.5005
R68443 VINN.n310 VINN.n194 4.5005
R68444 VINN.n260 VINN.n194 4.5005
R68445 VINN.n312 VINN.n194 4.5005
R68446 VINN.n259 VINN.n194 4.5005
R68447 VINN.n314 VINN.n194 4.5005
R68448 VINN.n258 VINN.n194 4.5005
R68449 VINN.n316 VINN.n194 4.5005
R68450 VINN.n257 VINN.n194 4.5005
R68451 VINN.n318 VINN.n194 4.5005
R68452 VINN.n256 VINN.n194 4.5005
R68453 VINN.n320 VINN.n194 4.5005
R68454 VINN.n255 VINN.n194 4.5005
R68455 VINN.n322 VINN.n194 4.5005
R68456 VINN.n254 VINN.n194 4.5005
R68457 VINN.n324 VINN.n194 4.5005
R68458 VINN.n253 VINN.n194 4.5005
R68459 VINN.n326 VINN.n194 4.5005
R68460 VINN.n252 VINN.n194 4.5005
R68461 VINN.n328 VINN.n194 4.5005
R68462 VINN.n251 VINN.n194 4.5005
R68463 VINN.n330 VINN.n194 4.5005
R68464 VINN.n250 VINN.n194 4.5005
R68465 VINN.n332 VINN.n194 4.5005
R68466 VINN.n249 VINN.n194 4.5005
R68467 VINN.n334 VINN.n194 4.5005
R68468 VINN.n248 VINN.n194 4.5005
R68469 VINN.n336 VINN.n194 4.5005
R68470 VINN.n247 VINN.n194 4.5005
R68471 VINN.n338 VINN.n194 4.5005
R68472 VINN.n246 VINN.n194 4.5005
R68473 VINN.n340 VINN.n194 4.5005
R68474 VINN.n245 VINN.n194 4.5005
R68475 VINN.n342 VINN.n194 4.5005
R68476 VINN.n244 VINN.n194 4.5005
R68477 VINN.n344 VINN.n194 4.5005
R68478 VINN.n243 VINN.n194 4.5005
R68479 VINN.n346 VINN.n194 4.5005
R68480 VINN.n242 VINN.n194 4.5005
R68481 VINN.n348 VINN.n194 4.5005
R68482 VINN.n241 VINN.n194 4.5005
R68483 VINN.n350 VINN.n194 4.5005
R68484 VINN.n240 VINN.n194 4.5005
R68485 VINN.n352 VINN.n194 4.5005
R68486 VINN.n239 VINN.n194 4.5005
R68487 VINN.n354 VINN.n194 4.5005
R68488 VINN.n238 VINN.n194 4.5005
R68489 VINN.n356 VINN.n194 4.5005
R68490 VINN.n237 VINN.n194 4.5005
R68491 VINN.n358 VINN.n194 4.5005
R68492 VINN.n236 VINN.n194 4.5005
R68493 VINN.n360 VINN.n194 4.5005
R68494 VINN.n235 VINN.n194 4.5005
R68495 VINN.n362 VINN.n194 4.5005
R68496 VINN.n234 VINN.n194 4.5005
R68497 VINN.n364 VINN.n194 4.5005
R68498 VINN.n233 VINN.n194 4.5005
R68499 VINN.n366 VINN.n194 4.5005
R68500 VINN.n232 VINN.n194 4.5005
R68501 VINN.n368 VINN.n194 4.5005
R68502 VINN.n231 VINN.n194 4.5005
R68503 VINN.n370 VINN.n194 4.5005
R68504 VINN.n230 VINN.n194 4.5005
R68505 VINN.n372 VINN.n194 4.5005
R68506 VINN.n229 VINN.n194 4.5005
R68507 VINN.n374 VINN.n194 4.5005
R68508 VINN.n228 VINN.n194 4.5005
R68509 VINN.n376 VINN.n194 4.5005
R68510 VINN.n227 VINN.n194 4.5005
R68511 VINN.n378 VINN.n194 4.5005
R68512 VINN.n226 VINN.n194 4.5005
R68513 VINN.n380 VINN.n194 4.5005
R68514 VINN.n225 VINN.n194 4.5005
R68515 VINN.n382 VINN.n194 4.5005
R68516 VINN.n224 VINN.n194 4.5005
R68517 VINN.n384 VINN.n194 4.5005
R68518 VINN.n223 VINN.n194 4.5005
R68519 VINN.n386 VINN.n194 4.5005
R68520 VINN.n222 VINN.n194 4.5005
R68521 VINN.n388 VINN.n194 4.5005
R68522 VINN.n221 VINN.n194 4.5005
R68523 VINN.n390 VINN.n194 4.5005
R68524 VINN.n220 VINN.n194 4.5005
R68525 VINN.n392 VINN.n194 4.5005
R68526 VINN.n219 VINN.n194 4.5005
R68527 VINN.n394 VINN.n194 4.5005
R68528 VINN.n218 VINN.n194 4.5005
R68529 VINN.n396 VINN.n194 4.5005
R68530 VINN.n217 VINN.n194 4.5005
R68531 VINN.n398 VINN.n194 4.5005
R68532 VINN.n216 VINN.n194 4.5005
R68533 VINN.n400 VINN.n194 4.5005
R68534 VINN.n215 VINN.n194 4.5005
R68535 VINN.n654 VINN.n194 4.5005
R68536 VINN.n656 VINN.n194 4.5005
R68537 VINN.n194 VINN.n0 4.5005
R68538 VINN.n278 VINN.n106 4.5005
R68539 VINN.n276 VINN.n106 4.5005
R68540 VINN.n280 VINN.n106 4.5005
R68541 VINN.n275 VINN.n106 4.5005
R68542 VINN.n282 VINN.n106 4.5005
R68543 VINN.n274 VINN.n106 4.5005
R68544 VINN.n284 VINN.n106 4.5005
R68545 VINN.n273 VINN.n106 4.5005
R68546 VINN.n286 VINN.n106 4.5005
R68547 VINN.n272 VINN.n106 4.5005
R68548 VINN.n288 VINN.n106 4.5005
R68549 VINN.n271 VINN.n106 4.5005
R68550 VINN.n290 VINN.n106 4.5005
R68551 VINN.n270 VINN.n106 4.5005
R68552 VINN.n292 VINN.n106 4.5005
R68553 VINN.n269 VINN.n106 4.5005
R68554 VINN.n294 VINN.n106 4.5005
R68555 VINN.n268 VINN.n106 4.5005
R68556 VINN.n296 VINN.n106 4.5005
R68557 VINN.n267 VINN.n106 4.5005
R68558 VINN.n298 VINN.n106 4.5005
R68559 VINN.n266 VINN.n106 4.5005
R68560 VINN.n300 VINN.n106 4.5005
R68561 VINN.n265 VINN.n106 4.5005
R68562 VINN.n302 VINN.n106 4.5005
R68563 VINN.n264 VINN.n106 4.5005
R68564 VINN.n304 VINN.n106 4.5005
R68565 VINN.n263 VINN.n106 4.5005
R68566 VINN.n306 VINN.n106 4.5005
R68567 VINN.n262 VINN.n106 4.5005
R68568 VINN.n308 VINN.n106 4.5005
R68569 VINN.n261 VINN.n106 4.5005
R68570 VINN.n310 VINN.n106 4.5005
R68571 VINN.n260 VINN.n106 4.5005
R68572 VINN.n312 VINN.n106 4.5005
R68573 VINN.n259 VINN.n106 4.5005
R68574 VINN.n314 VINN.n106 4.5005
R68575 VINN.n258 VINN.n106 4.5005
R68576 VINN.n316 VINN.n106 4.5005
R68577 VINN.n257 VINN.n106 4.5005
R68578 VINN.n318 VINN.n106 4.5005
R68579 VINN.n256 VINN.n106 4.5005
R68580 VINN.n320 VINN.n106 4.5005
R68581 VINN.n255 VINN.n106 4.5005
R68582 VINN.n322 VINN.n106 4.5005
R68583 VINN.n254 VINN.n106 4.5005
R68584 VINN.n324 VINN.n106 4.5005
R68585 VINN.n253 VINN.n106 4.5005
R68586 VINN.n326 VINN.n106 4.5005
R68587 VINN.n252 VINN.n106 4.5005
R68588 VINN.n328 VINN.n106 4.5005
R68589 VINN.n251 VINN.n106 4.5005
R68590 VINN.n330 VINN.n106 4.5005
R68591 VINN.n250 VINN.n106 4.5005
R68592 VINN.n332 VINN.n106 4.5005
R68593 VINN.n249 VINN.n106 4.5005
R68594 VINN.n334 VINN.n106 4.5005
R68595 VINN.n248 VINN.n106 4.5005
R68596 VINN.n336 VINN.n106 4.5005
R68597 VINN.n247 VINN.n106 4.5005
R68598 VINN.n338 VINN.n106 4.5005
R68599 VINN.n246 VINN.n106 4.5005
R68600 VINN.n340 VINN.n106 4.5005
R68601 VINN.n245 VINN.n106 4.5005
R68602 VINN.n342 VINN.n106 4.5005
R68603 VINN.n244 VINN.n106 4.5005
R68604 VINN.n344 VINN.n106 4.5005
R68605 VINN.n243 VINN.n106 4.5005
R68606 VINN.n346 VINN.n106 4.5005
R68607 VINN.n242 VINN.n106 4.5005
R68608 VINN.n348 VINN.n106 4.5005
R68609 VINN.n241 VINN.n106 4.5005
R68610 VINN.n350 VINN.n106 4.5005
R68611 VINN.n240 VINN.n106 4.5005
R68612 VINN.n352 VINN.n106 4.5005
R68613 VINN.n239 VINN.n106 4.5005
R68614 VINN.n354 VINN.n106 4.5005
R68615 VINN.n238 VINN.n106 4.5005
R68616 VINN.n356 VINN.n106 4.5005
R68617 VINN.n237 VINN.n106 4.5005
R68618 VINN.n358 VINN.n106 4.5005
R68619 VINN.n236 VINN.n106 4.5005
R68620 VINN.n360 VINN.n106 4.5005
R68621 VINN.n235 VINN.n106 4.5005
R68622 VINN.n362 VINN.n106 4.5005
R68623 VINN.n234 VINN.n106 4.5005
R68624 VINN.n364 VINN.n106 4.5005
R68625 VINN.n233 VINN.n106 4.5005
R68626 VINN.n366 VINN.n106 4.5005
R68627 VINN.n232 VINN.n106 4.5005
R68628 VINN.n368 VINN.n106 4.5005
R68629 VINN.n231 VINN.n106 4.5005
R68630 VINN.n370 VINN.n106 4.5005
R68631 VINN.n230 VINN.n106 4.5005
R68632 VINN.n372 VINN.n106 4.5005
R68633 VINN.n229 VINN.n106 4.5005
R68634 VINN.n374 VINN.n106 4.5005
R68635 VINN.n228 VINN.n106 4.5005
R68636 VINN.n376 VINN.n106 4.5005
R68637 VINN.n227 VINN.n106 4.5005
R68638 VINN.n378 VINN.n106 4.5005
R68639 VINN.n226 VINN.n106 4.5005
R68640 VINN.n380 VINN.n106 4.5005
R68641 VINN.n225 VINN.n106 4.5005
R68642 VINN.n382 VINN.n106 4.5005
R68643 VINN.n224 VINN.n106 4.5005
R68644 VINN.n384 VINN.n106 4.5005
R68645 VINN.n223 VINN.n106 4.5005
R68646 VINN.n386 VINN.n106 4.5005
R68647 VINN.n222 VINN.n106 4.5005
R68648 VINN.n388 VINN.n106 4.5005
R68649 VINN.n221 VINN.n106 4.5005
R68650 VINN.n390 VINN.n106 4.5005
R68651 VINN.n220 VINN.n106 4.5005
R68652 VINN.n392 VINN.n106 4.5005
R68653 VINN.n219 VINN.n106 4.5005
R68654 VINN.n394 VINN.n106 4.5005
R68655 VINN.n218 VINN.n106 4.5005
R68656 VINN.n396 VINN.n106 4.5005
R68657 VINN.n217 VINN.n106 4.5005
R68658 VINN.n398 VINN.n106 4.5005
R68659 VINN.n216 VINN.n106 4.5005
R68660 VINN.n400 VINN.n106 4.5005
R68661 VINN.n215 VINN.n106 4.5005
R68662 VINN.n654 VINN.n106 4.5005
R68663 VINN.n656 VINN.n106 4.5005
R68664 VINN.n106 VINN.n0 4.5005
R68665 VINN.n278 VINN.n195 4.5005
R68666 VINN.n276 VINN.n195 4.5005
R68667 VINN.n280 VINN.n195 4.5005
R68668 VINN.n275 VINN.n195 4.5005
R68669 VINN.n282 VINN.n195 4.5005
R68670 VINN.n274 VINN.n195 4.5005
R68671 VINN.n284 VINN.n195 4.5005
R68672 VINN.n273 VINN.n195 4.5005
R68673 VINN.n286 VINN.n195 4.5005
R68674 VINN.n272 VINN.n195 4.5005
R68675 VINN.n288 VINN.n195 4.5005
R68676 VINN.n271 VINN.n195 4.5005
R68677 VINN.n290 VINN.n195 4.5005
R68678 VINN.n270 VINN.n195 4.5005
R68679 VINN.n292 VINN.n195 4.5005
R68680 VINN.n269 VINN.n195 4.5005
R68681 VINN.n294 VINN.n195 4.5005
R68682 VINN.n268 VINN.n195 4.5005
R68683 VINN.n296 VINN.n195 4.5005
R68684 VINN.n267 VINN.n195 4.5005
R68685 VINN.n298 VINN.n195 4.5005
R68686 VINN.n266 VINN.n195 4.5005
R68687 VINN.n300 VINN.n195 4.5005
R68688 VINN.n265 VINN.n195 4.5005
R68689 VINN.n302 VINN.n195 4.5005
R68690 VINN.n264 VINN.n195 4.5005
R68691 VINN.n304 VINN.n195 4.5005
R68692 VINN.n263 VINN.n195 4.5005
R68693 VINN.n306 VINN.n195 4.5005
R68694 VINN.n262 VINN.n195 4.5005
R68695 VINN.n308 VINN.n195 4.5005
R68696 VINN.n261 VINN.n195 4.5005
R68697 VINN.n310 VINN.n195 4.5005
R68698 VINN.n260 VINN.n195 4.5005
R68699 VINN.n312 VINN.n195 4.5005
R68700 VINN.n259 VINN.n195 4.5005
R68701 VINN.n314 VINN.n195 4.5005
R68702 VINN.n258 VINN.n195 4.5005
R68703 VINN.n316 VINN.n195 4.5005
R68704 VINN.n257 VINN.n195 4.5005
R68705 VINN.n318 VINN.n195 4.5005
R68706 VINN.n256 VINN.n195 4.5005
R68707 VINN.n320 VINN.n195 4.5005
R68708 VINN.n255 VINN.n195 4.5005
R68709 VINN.n322 VINN.n195 4.5005
R68710 VINN.n254 VINN.n195 4.5005
R68711 VINN.n324 VINN.n195 4.5005
R68712 VINN.n253 VINN.n195 4.5005
R68713 VINN.n326 VINN.n195 4.5005
R68714 VINN.n252 VINN.n195 4.5005
R68715 VINN.n328 VINN.n195 4.5005
R68716 VINN.n251 VINN.n195 4.5005
R68717 VINN.n330 VINN.n195 4.5005
R68718 VINN.n250 VINN.n195 4.5005
R68719 VINN.n332 VINN.n195 4.5005
R68720 VINN.n249 VINN.n195 4.5005
R68721 VINN.n334 VINN.n195 4.5005
R68722 VINN.n248 VINN.n195 4.5005
R68723 VINN.n336 VINN.n195 4.5005
R68724 VINN.n247 VINN.n195 4.5005
R68725 VINN.n338 VINN.n195 4.5005
R68726 VINN.n246 VINN.n195 4.5005
R68727 VINN.n340 VINN.n195 4.5005
R68728 VINN.n245 VINN.n195 4.5005
R68729 VINN.n342 VINN.n195 4.5005
R68730 VINN.n244 VINN.n195 4.5005
R68731 VINN.n344 VINN.n195 4.5005
R68732 VINN.n243 VINN.n195 4.5005
R68733 VINN.n346 VINN.n195 4.5005
R68734 VINN.n242 VINN.n195 4.5005
R68735 VINN.n348 VINN.n195 4.5005
R68736 VINN.n241 VINN.n195 4.5005
R68737 VINN.n350 VINN.n195 4.5005
R68738 VINN.n240 VINN.n195 4.5005
R68739 VINN.n352 VINN.n195 4.5005
R68740 VINN.n239 VINN.n195 4.5005
R68741 VINN.n354 VINN.n195 4.5005
R68742 VINN.n238 VINN.n195 4.5005
R68743 VINN.n356 VINN.n195 4.5005
R68744 VINN.n237 VINN.n195 4.5005
R68745 VINN.n358 VINN.n195 4.5005
R68746 VINN.n236 VINN.n195 4.5005
R68747 VINN.n360 VINN.n195 4.5005
R68748 VINN.n235 VINN.n195 4.5005
R68749 VINN.n362 VINN.n195 4.5005
R68750 VINN.n234 VINN.n195 4.5005
R68751 VINN.n364 VINN.n195 4.5005
R68752 VINN.n233 VINN.n195 4.5005
R68753 VINN.n366 VINN.n195 4.5005
R68754 VINN.n232 VINN.n195 4.5005
R68755 VINN.n368 VINN.n195 4.5005
R68756 VINN.n231 VINN.n195 4.5005
R68757 VINN.n370 VINN.n195 4.5005
R68758 VINN.n230 VINN.n195 4.5005
R68759 VINN.n372 VINN.n195 4.5005
R68760 VINN.n229 VINN.n195 4.5005
R68761 VINN.n374 VINN.n195 4.5005
R68762 VINN.n228 VINN.n195 4.5005
R68763 VINN.n376 VINN.n195 4.5005
R68764 VINN.n227 VINN.n195 4.5005
R68765 VINN.n378 VINN.n195 4.5005
R68766 VINN.n226 VINN.n195 4.5005
R68767 VINN.n380 VINN.n195 4.5005
R68768 VINN.n225 VINN.n195 4.5005
R68769 VINN.n382 VINN.n195 4.5005
R68770 VINN.n224 VINN.n195 4.5005
R68771 VINN.n384 VINN.n195 4.5005
R68772 VINN.n223 VINN.n195 4.5005
R68773 VINN.n386 VINN.n195 4.5005
R68774 VINN.n222 VINN.n195 4.5005
R68775 VINN.n388 VINN.n195 4.5005
R68776 VINN.n221 VINN.n195 4.5005
R68777 VINN.n390 VINN.n195 4.5005
R68778 VINN.n220 VINN.n195 4.5005
R68779 VINN.n392 VINN.n195 4.5005
R68780 VINN.n219 VINN.n195 4.5005
R68781 VINN.n394 VINN.n195 4.5005
R68782 VINN.n218 VINN.n195 4.5005
R68783 VINN.n396 VINN.n195 4.5005
R68784 VINN.n217 VINN.n195 4.5005
R68785 VINN.n398 VINN.n195 4.5005
R68786 VINN.n216 VINN.n195 4.5005
R68787 VINN.n400 VINN.n195 4.5005
R68788 VINN.n215 VINN.n195 4.5005
R68789 VINN.n654 VINN.n195 4.5005
R68790 VINN.n656 VINN.n195 4.5005
R68791 VINN.n195 VINN.n0 4.5005
R68792 VINN.n278 VINN.n105 4.5005
R68793 VINN.n276 VINN.n105 4.5005
R68794 VINN.n280 VINN.n105 4.5005
R68795 VINN.n275 VINN.n105 4.5005
R68796 VINN.n282 VINN.n105 4.5005
R68797 VINN.n274 VINN.n105 4.5005
R68798 VINN.n284 VINN.n105 4.5005
R68799 VINN.n273 VINN.n105 4.5005
R68800 VINN.n286 VINN.n105 4.5005
R68801 VINN.n272 VINN.n105 4.5005
R68802 VINN.n288 VINN.n105 4.5005
R68803 VINN.n271 VINN.n105 4.5005
R68804 VINN.n290 VINN.n105 4.5005
R68805 VINN.n270 VINN.n105 4.5005
R68806 VINN.n292 VINN.n105 4.5005
R68807 VINN.n269 VINN.n105 4.5005
R68808 VINN.n294 VINN.n105 4.5005
R68809 VINN.n268 VINN.n105 4.5005
R68810 VINN.n296 VINN.n105 4.5005
R68811 VINN.n267 VINN.n105 4.5005
R68812 VINN.n298 VINN.n105 4.5005
R68813 VINN.n266 VINN.n105 4.5005
R68814 VINN.n300 VINN.n105 4.5005
R68815 VINN.n265 VINN.n105 4.5005
R68816 VINN.n302 VINN.n105 4.5005
R68817 VINN.n264 VINN.n105 4.5005
R68818 VINN.n304 VINN.n105 4.5005
R68819 VINN.n263 VINN.n105 4.5005
R68820 VINN.n306 VINN.n105 4.5005
R68821 VINN.n262 VINN.n105 4.5005
R68822 VINN.n308 VINN.n105 4.5005
R68823 VINN.n261 VINN.n105 4.5005
R68824 VINN.n310 VINN.n105 4.5005
R68825 VINN.n260 VINN.n105 4.5005
R68826 VINN.n312 VINN.n105 4.5005
R68827 VINN.n259 VINN.n105 4.5005
R68828 VINN.n314 VINN.n105 4.5005
R68829 VINN.n258 VINN.n105 4.5005
R68830 VINN.n316 VINN.n105 4.5005
R68831 VINN.n257 VINN.n105 4.5005
R68832 VINN.n318 VINN.n105 4.5005
R68833 VINN.n256 VINN.n105 4.5005
R68834 VINN.n320 VINN.n105 4.5005
R68835 VINN.n255 VINN.n105 4.5005
R68836 VINN.n322 VINN.n105 4.5005
R68837 VINN.n254 VINN.n105 4.5005
R68838 VINN.n324 VINN.n105 4.5005
R68839 VINN.n253 VINN.n105 4.5005
R68840 VINN.n326 VINN.n105 4.5005
R68841 VINN.n252 VINN.n105 4.5005
R68842 VINN.n328 VINN.n105 4.5005
R68843 VINN.n251 VINN.n105 4.5005
R68844 VINN.n330 VINN.n105 4.5005
R68845 VINN.n250 VINN.n105 4.5005
R68846 VINN.n332 VINN.n105 4.5005
R68847 VINN.n249 VINN.n105 4.5005
R68848 VINN.n334 VINN.n105 4.5005
R68849 VINN.n248 VINN.n105 4.5005
R68850 VINN.n336 VINN.n105 4.5005
R68851 VINN.n247 VINN.n105 4.5005
R68852 VINN.n338 VINN.n105 4.5005
R68853 VINN.n246 VINN.n105 4.5005
R68854 VINN.n340 VINN.n105 4.5005
R68855 VINN.n245 VINN.n105 4.5005
R68856 VINN.n342 VINN.n105 4.5005
R68857 VINN.n244 VINN.n105 4.5005
R68858 VINN.n344 VINN.n105 4.5005
R68859 VINN.n243 VINN.n105 4.5005
R68860 VINN.n346 VINN.n105 4.5005
R68861 VINN.n242 VINN.n105 4.5005
R68862 VINN.n348 VINN.n105 4.5005
R68863 VINN.n241 VINN.n105 4.5005
R68864 VINN.n350 VINN.n105 4.5005
R68865 VINN.n240 VINN.n105 4.5005
R68866 VINN.n352 VINN.n105 4.5005
R68867 VINN.n239 VINN.n105 4.5005
R68868 VINN.n354 VINN.n105 4.5005
R68869 VINN.n238 VINN.n105 4.5005
R68870 VINN.n356 VINN.n105 4.5005
R68871 VINN.n237 VINN.n105 4.5005
R68872 VINN.n358 VINN.n105 4.5005
R68873 VINN.n236 VINN.n105 4.5005
R68874 VINN.n360 VINN.n105 4.5005
R68875 VINN.n235 VINN.n105 4.5005
R68876 VINN.n362 VINN.n105 4.5005
R68877 VINN.n234 VINN.n105 4.5005
R68878 VINN.n364 VINN.n105 4.5005
R68879 VINN.n233 VINN.n105 4.5005
R68880 VINN.n366 VINN.n105 4.5005
R68881 VINN.n232 VINN.n105 4.5005
R68882 VINN.n368 VINN.n105 4.5005
R68883 VINN.n231 VINN.n105 4.5005
R68884 VINN.n370 VINN.n105 4.5005
R68885 VINN.n230 VINN.n105 4.5005
R68886 VINN.n372 VINN.n105 4.5005
R68887 VINN.n229 VINN.n105 4.5005
R68888 VINN.n374 VINN.n105 4.5005
R68889 VINN.n228 VINN.n105 4.5005
R68890 VINN.n376 VINN.n105 4.5005
R68891 VINN.n227 VINN.n105 4.5005
R68892 VINN.n378 VINN.n105 4.5005
R68893 VINN.n226 VINN.n105 4.5005
R68894 VINN.n380 VINN.n105 4.5005
R68895 VINN.n225 VINN.n105 4.5005
R68896 VINN.n382 VINN.n105 4.5005
R68897 VINN.n224 VINN.n105 4.5005
R68898 VINN.n384 VINN.n105 4.5005
R68899 VINN.n223 VINN.n105 4.5005
R68900 VINN.n386 VINN.n105 4.5005
R68901 VINN.n222 VINN.n105 4.5005
R68902 VINN.n388 VINN.n105 4.5005
R68903 VINN.n221 VINN.n105 4.5005
R68904 VINN.n390 VINN.n105 4.5005
R68905 VINN.n220 VINN.n105 4.5005
R68906 VINN.n392 VINN.n105 4.5005
R68907 VINN.n219 VINN.n105 4.5005
R68908 VINN.n394 VINN.n105 4.5005
R68909 VINN.n218 VINN.n105 4.5005
R68910 VINN.n396 VINN.n105 4.5005
R68911 VINN.n217 VINN.n105 4.5005
R68912 VINN.n398 VINN.n105 4.5005
R68913 VINN.n216 VINN.n105 4.5005
R68914 VINN.n400 VINN.n105 4.5005
R68915 VINN.n215 VINN.n105 4.5005
R68916 VINN.n654 VINN.n105 4.5005
R68917 VINN.n656 VINN.n105 4.5005
R68918 VINN.n105 VINN.n0 4.5005
R68919 VINN.n278 VINN.n196 4.5005
R68920 VINN.n276 VINN.n196 4.5005
R68921 VINN.n280 VINN.n196 4.5005
R68922 VINN.n275 VINN.n196 4.5005
R68923 VINN.n282 VINN.n196 4.5005
R68924 VINN.n274 VINN.n196 4.5005
R68925 VINN.n284 VINN.n196 4.5005
R68926 VINN.n273 VINN.n196 4.5005
R68927 VINN.n286 VINN.n196 4.5005
R68928 VINN.n272 VINN.n196 4.5005
R68929 VINN.n288 VINN.n196 4.5005
R68930 VINN.n271 VINN.n196 4.5005
R68931 VINN.n290 VINN.n196 4.5005
R68932 VINN.n270 VINN.n196 4.5005
R68933 VINN.n292 VINN.n196 4.5005
R68934 VINN.n269 VINN.n196 4.5005
R68935 VINN.n294 VINN.n196 4.5005
R68936 VINN.n268 VINN.n196 4.5005
R68937 VINN.n296 VINN.n196 4.5005
R68938 VINN.n267 VINN.n196 4.5005
R68939 VINN.n298 VINN.n196 4.5005
R68940 VINN.n266 VINN.n196 4.5005
R68941 VINN.n300 VINN.n196 4.5005
R68942 VINN.n265 VINN.n196 4.5005
R68943 VINN.n302 VINN.n196 4.5005
R68944 VINN.n264 VINN.n196 4.5005
R68945 VINN.n304 VINN.n196 4.5005
R68946 VINN.n263 VINN.n196 4.5005
R68947 VINN.n306 VINN.n196 4.5005
R68948 VINN.n262 VINN.n196 4.5005
R68949 VINN.n308 VINN.n196 4.5005
R68950 VINN.n261 VINN.n196 4.5005
R68951 VINN.n310 VINN.n196 4.5005
R68952 VINN.n260 VINN.n196 4.5005
R68953 VINN.n312 VINN.n196 4.5005
R68954 VINN.n259 VINN.n196 4.5005
R68955 VINN.n314 VINN.n196 4.5005
R68956 VINN.n258 VINN.n196 4.5005
R68957 VINN.n316 VINN.n196 4.5005
R68958 VINN.n257 VINN.n196 4.5005
R68959 VINN.n318 VINN.n196 4.5005
R68960 VINN.n256 VINN.n196 4.5005
R68961 VINN.n320 VINN.n196 4.5005
R68962 VINN.n255 VINN.n196 4.5005
R68963 VINN.n322 VINN.n196 4.5005
R68964 VINN.n254 VINN.n196 4.5005
R68965 VINN.n324 VINN.n196 4.5005
R68966 VINN.n253 VINN.n196 4.5005
R68967 VINN.n326 VINN.n196 4.5005
R68968 VINN.n252 VINN.n196 4.5005
R68969 VINN.n328 VINN.n196 4.5005
R68970 VINN.n251 VINN.n196 4.5005
R68971 VINN.n330 VINN.n196 4.5005
R68972 VINN.n250 VINN.n196 4.5005
R68973 VINN.n332 VINN.n196 4.5005
R68974 VINN.n249 VINN.n196 4.5005
R68975 VINN.n334 VINN.n196 4.5005
R68976 VINN.n248 VINN.n196 4.5005
R68977 VINN.n336 VINN.n196 4.5005
R68978 VINN.n247 VINN.n196 4.5005
R68979 VINN.n338 VINN.n196 4.5005
R68980 VINN.n246 VINN.n196 4.5005
R68981 VINN.n340 VINN.n196 4.5005
R68982 VINN.n245 VINN.n196 4.5005
R68983 VINN.n342 VINN.n196 4.5005
R68984 VINN.n244 VINN.n196 4.5005
R68985 VINN.n344 VINN.n196 4.5005
R68986 VINN.n243 VINN.n196 4.5005
R68987 VINN.n346 VINN.n196 4.5005
R68988 VINN.n242 VINN.n196 4.5005
R68989 VINN.n348 VINN.n196 4.5005
R68990 VINN.n241 VINN.n196 4.5005
R68991 VINN.n350 VINN.n196 4.5005
R68992 VINN.n240 VINN.n196 4.5005
R68993 VINN.n352 VINN.n196 4.5005
R68994 VINN.n239 VINN.n196 4.5005
R68995 VINN.n354 VINN.n196 4.5005
R68996 VINN.n238 VINN.n196 4.5005
R68997 VINN.n356 VINN.n196 4.5005
R68998 VINN.n237 VINN.n196 4.5005
R68999 VINN.n358 VINN.n196 4.5005
R69000 VINN.n236 VINN.n196 4.5005
R69001 VINN.n360 VINN.n196 4.5005
R69002 VINN.n235 VINN.n196 4.5005
R69003 VINN.n362 VINN.n196 4.5005
R69004 VINN.n234 VINN.n196 4.5005
R69005 VINN.n364 VINN.n196 4.5005
R69006 VINN.n233 VINN.n196 4.5005
R69007 VINN.n366 VINN.n196 4.5005
R69008 VINN.n232 VINN.n196 4.5005
R69009 VINN.n368 VINN.n196 4.5005
R69010 VINN.n231 VINN.n196 4.5005
R69011 VINN.n370 VINN.n196 4.5005
R69012 VINN.n230 VINN.n196 4.5005
R69013 VINN.n372 VINN.n196 4.5005
R69014 VINN.n229 VINN.n196 4.5005
R69015 VINN.n374 VINN.n196 4.5005
R69016 VINN.n228 VINN.n196 4.5005
R69017 VINN.n376 VINN.n196 4.5005
R69018 VINN.n227 VINN.n196 4.5005
R69019 VINN.n378 VINN.n196 4.5005
R69020 VINN.n226 VINN.n196 4.5005
R69021 VINN.n380 VINN.n196 4.5005
R69022 VINN.n225 VINN.n196 4.5005
R69023 VINN.n382 VINN.n196 4.5005
R69024 VINN.n224 VINN.n196 4.5005
R69025 VINN.n384 VINN.n196 4.5005
R69026 VINN.n223 VINN.n196 4.5005
R69027 VINN.n386 VINN.n196 4.5005
R69028 VINN.n222 VINN.n196 4.5005
R69029 VINN.n388 VINN.n196 4.5005
R69030 VINN.n221 VINN.n196 4.5005
R69031 VINN.n390 VINN.n196 4.5005
R69032 VINN.n220 VINN.n196 4.5005
R69033 VINN.n392 VINN.n196 4.5005
R69034 VINN.n219 VINN.n196 4.5005
R69035 VINN.n394 VINN.n196 4.5005
R69036 VINN.n218 VINN.n196 4.5005
R69037 VINN.n396 VINN.n196 4.5005
R69038 VINN.n217 VINN.n196 4.5005
R69039 VINN.n398 VINN.n196 4.5005
R69040 VINN.n216 VINN.n196 4.5005
R69041 VINN.n400 VINN.n196 4.5005
R69042 VINN.n215 VINN.n196 4.5005
R69043 VINN.n654 VINN.n196 4.5005
R69044 VINN.n656 VINN.n196 4.5005
R69045 VINN.n196 VINN.n0 4.5005
R69046 VINN.n278 VINN.n104 4.5005
R69047 VINN.n276 VINN.n104 4.5005
R69048 VINN.n280 VINN.n104 4.5005
R69049 VINN.n275 VINN.n104 4.5005
R69050 VINN.n282 VINN.n104 4.5005
R69051 VINN.n274 VINN.n104 4.5005
R69052 VINN.n284 VINN.n104 4.5005
R69053 VINN.n273 VINN.n104 4.5005
R69054 VINN.n286 VINN.n104 4.5005
R69055 VINN.n272 VINN.n104 4.5005
R69056 VINN.n288 VINN.n104 4.5005
R69057 VINN.n271 VINN.n104 4.5005
R69058 VINN.n290 VINN.n104 4.5005
R69059 VINN.n270 VINN.n104 4.5005
R69060 VINN.n292 VINN.n104 4.5005
R69061 VINN.n269 VINN.n104 4.5005
R69062 VINN.n294 VINN.n104 4.5005
R69063 VINN.n268 VINN.n104 4.5005
R69064 VINN.n296 VINN.n104 4.5005
R69065 VINN.n267 VINN.n104 4.5005
R69066 VINN.n298 VINN.n104 4.5005
R69067 VINN.n266 VINN.n104 4.5005
R69068 VINN.n300 VINN.n104 4.5005
R69069 VINN.n265 VINN.n104 4.5005
R69070 VINN.n302 VINN.n104 4.5005
R69071 VINN.n264 VINN.n104 4.5005
R69072 VINN.n304 VINN.n104 4.5005
R69073 VINN.n263 VINN.n104 4.5005
R69074 VINN.n306 VINN.n104 4.5005
R69075 VINN.n262 VINN.n104 4.5005
R69076 VINN.n308 VINN.n104 4.5005
R69077 VINN.n261 VINN.n104 4.5005
R69078 VINN.n310 VINN.n104 4.5005
R69079 VINN.n260 VINN.n104 4.5005
R69080 VINN.n312 VINN.n104 4.5005
R69081 VINN.n259 VINN.n104 4.5005
R69082 VINN.n314 VINN.n104 4.5005
R69083 VINN.n258 VINN.n104 4.5005
R69084 VINN.n316 VINN.n104 4.5005
R69085 VINN.n257 VINN.n104 4.5005
R69086 VINN.n318 VINN.n104 4.5005
R69087 VINN.n256 VINN.n104 4.5005
R69088 VINN.n320 VINN.n104 4.5005
R69089 VINN.n255 VINN.n104 4.5005
R69090 VINN.n322 VINN.n104 4.5005
R69091 VINN.n254 VINN.n104 4.5005
R69092 VINN.n324 VINN.n104 4.5005
R69093 VINN.n253 VINN.n104 4.5005
R69094 VINN.n326 VINN.n104 4.5005
R69095 VINN.n252 VINN.n104 4.5005
R69096 VINN.n328 VINN.n104 4.5005
R69097 VINN.n251 VINN.n104 4.5005
R69098 VINN.n330 VINN.n104 4.5005
R69099 VINN.n250 VINN.n104 4.5005
R69100 VINN.n332 VINN.n104 4.5005
R69101 VINN.n249 VINN.n104 4.5005
R69102 VINN.n334 VINN.n104 4.5005
R69103 VINN.n248 VINN.n104 4.5005
R69104 VINN.n336 VINN.n104 4.5005
R69105 VINN.n247 VINN.n104 4.5005
R69106 VINN.n338 VINN.n104 4.5005
R69107 VINN.n246 VINN.n104 4.5005
R69108 VINN.n340 VINN.n104 4.5005
R69109 VINN.n245 VINN.n104 4.5005
R69110 VINN.n342 VINN.n104 4.5005
R69111 VINN.n244 VINN.n104 4.5005
R69112 VINN.n344 VINN.n104 4.5005
R69113 VINN.n243 VINN.n104 4.5005
R69114 VINN.n346 VINN.n104 4.5005
R69115 VINN.n242 VINN.n104 4.5005
R69116 VINN.n348 VINN.n104 4.5005
R69117 VINN.n241 VINN.n104 4.5005
R69118 VINN.n350 VINN.n104 4.5005
R69119 VINN.n240 VINN.n104 4.5005
R69120 VINN.n352 VINN.n104 4.5005
R69121 VINN.n239 VINN.n104 4.5005
R69122 VINN.n354 VINN.n104 4.5005
R69123 VINN.n238 VINN.n104 4.5005
R69124 VINN.n356 VINN.n104 4.5005
R69125 VINN.n237 VINN.n104 4.5005
R69126 VINN.n358 VINN.n104 4.5005
R69127 VINN.n236 VINN.n104 4.5005
R69128 VINN.n360 VINN.n104 4.5005
R69129 VINN.n235 VINN.n104 4.5005
R69130 VINN.n362 VINN.n104 4.5005
R69131 VINN.n234 VINN.n104 4.5005
R69132 VINN.n364 VINN.n104 4.5005
R69133 VINN.n233 VINN.n104 4.5005
R69134 VINN.n366 VINN.n104 4.5005
R69135 VINN.n232 VINN.n104 4.5005
R69136 VINN.n368 VINN.n104 4.5005
R69137 VINN.n231 VINN.n104 4.5005
R69138 VINN.n370 VINN.n104 4.5005
R69139 VINN.n230 VINN.n104 4.5005
R69140 VINN.n372 VINN.n104 4.5005
R69141 VINN.n229 VINN.n104 4.5005
R69142 VINN.n374 VINN.n104 4.5005
R69143 VINN.n228 VINN.n104 4.5005
R69144 VINN.n376 VINN.n104 4.5005
R69145 VINN.n227 VINN.n104 4.5005
R69146 VINN.n378 VINN.n104 4.5005
R69147 VINN.n226 VINN.n104 4.5005
R69148 VINN.n380 VINN.n104 4.5005
R69149 VINN.n225 VINN.n104 4.5005
R69150 VINN.n382 VINN.n104 4.5005
R69151 VINN.n224 VINN.n104 4.5005
R69152 VINN.n384 VINN.n104 4.5005
R69153 VINN.n223 VINN.n104 4.5005
R69154 VINN.n386 VINN.n104 4.5005
R69155 VINN.n222 VINN.n104 4.5005
R69156 VINN.n388 VINN.n104 4.5005
R69157 VINN.n221 VINN.n104 4.5005
R69158 VINN.n390 VINN.n104 4.5005
R69159 VINN.n220 VINN.n104 4.5005
R69160 VINN.n392 VINN.n104 4.5005
R69161 VINN.n219 VINN.n104 4.5005
R69162 VINN.n394 VINN.n104 4.5005
R69163 VINN.n218 VINN.n104 4.5005
R69164 VINN.n396 VINN.n104 4.5005
R69165 VINN.n217 VINN.n104 4.5005
R69166 VINN.n398 VINN.n104 4.5005
R69167 VINN.n216 VINN.n104 4.5005
R69168 VINN.n400 VINN.n104 4.5005
R69169 VINN.n215 VINN.n104 4.5005
R69170 VINN.n654 VINN.n104 4.5005
R69171 VINN.n656 VINN.n104 4.5005
R69172 VINN.n104 VINN.n0 4.5005
R69173 VINN.n278 VINN.n197 4.5005
R69174 VINN.n276 VINN.n197 4.5005
R69175 VINN.n280 VINN.n197 4.5005
R69176 VINN.n275 VINN.n197 4.5005
R69177 VINN.n282 VINN.n197 4.5005
R69178 VINN.n274 VINN.n197 4.5005
R69179 VINN.n284 VINN.n197 4.5005
R69180 VINN.n273 VINN.n197 4.5005
R69181 VINN.n286 VINN.n197 4.5005
R69182 VINN.n272 VINN.n197 4.5005
R69183 VINN.n288 VINN.n197 4.5005
R69184 VINN.n271 VINN.n197 4.5005
R69185 VINN.n290 VINN.n197 4.5005
R69186 VINN.n270 VINN.n197 4.5005
R69187 VINN.n292 VINN.n197 4.5005
R69188 VINN.n269 VINN.n197 4.5005
R69189 VINN.n294 VINN.n197 4.5005
R69190 VINN.n268 VINN.n197 4.5005
R69191 VINN.n296 VINN.n197 4.5005
R69192 VINN.n267 VINN.n197 4.5005
R69193 VINN.n298 VINN.n197 4.5005
R69194 VINN.n266 VINN.n197 4.5005
R69195 VINN.n300 VINN.n197 4.5005
R69196 VINN.n265 VINN.n197 4.5005
R69197 VINN.n302 VINN.n197 4.5005
R69198 VINN.n264 VINN.n197 4.5005
R69199 VINN.n304 VINN.n197 4.5005
R69200 VINN.n263 VINN.n197 4.5005
R69201 VINN.n306 VINN.n197 4.5005
R69202 VINN.n262 VINN.n197 4.5005
R69203 VINN.n308 VINN.n197 4.5005
R69204 VINN.n261 VINN.n197 4.5005
R69205 VINN.n310 VINN.n197 4.5005
R69206 VINN.n260 VINN.n197 4.5005
R69207 VINN.n312 VINN.n197 4.5005
R69208 VINN.n259 VINN.n197 4.5005
R69209 VINN.n314 VINN.n197 4.5005
R69210 VINN.n258 VINN.n197 4.5005
R69211 VINN.n316 VINN.n197 4.5005
R69212 VINN.n257 VINN.n197 4.5005
R69213 VINN.n318 VINN.n197 4.5005
R69214 VINN.n256 VINN.n197 4.5005
R69215 VINN.n320 VINN.n197 4.5005
R69216 VINN.n255 VINN.n197 4.5005
R69217 VINN.n322 VINN.n197 4.5005
R69218 VINN.n254 VINN.n197 4.5005
R69219 VINN.n324 VINN.n197 4.5005
R69220 VINN.n253 VINN.n197 4.5005
R69221 VINN.n326 VINN.n197 4.5005
R69222 VINN.n252 VINN.n197 4.5005
R69223 VINN.n328 VINN.n197 4.5005
R69224 VINN.n251 VINN.n197 4.5005
R69225 VINN.n330 VINN.n197 4.5005
R69226 VINN.n250 VINN.n197 4.5005
R69227 VINN.n332 VINN.n197 4.5005
R69228 VINN.n249 VINN.n197 4.5005
R69229 VINN.n334 VINN.n197 4.5005
R69230 VINN.n248 VINN.n197 4.5005
R69231 VINN.n336 VINN.n197 4.5005
R69232 VINN.n247 VINN.n197 4.5005
R69233 VINN.n338 VINN.n197 4.5005
R69234 VINN.n246 VINN.n197 4.5005
R69235 VINN.n340 VINN.n197 4.5005
R69236 VINN.n245 VINN.n197 4.5005
R69237 VINN.n342 VINN.n197 4.5005
R69238 VINN.n244 VINN.n197 4.5005
R69239 VINN.n344 VINN.n197 4.5005
R69240 VINN.n243 VINN.n197 4.5005
R69241 VINN.n346 VINN.n197 4.5005
R69242 VINN.n242 VINN.n197 4.5005
R69243 VINN.n348 VINN.n197 4.5005
R69244 VINN.n241 VINN.n197 4.5005
R69245 VINN.n350 VINN.n197 4.5005
R69246 VINN.n240 VINN.n197 4.5005
R69247 VINN.n352 VINN.n197 4.5005
R69248 VINN.n239 VINN.n197 4.5005
R69249 VINN.n354 VINN.n197 4.5005
R69250 VINN.n238 VINN.n197 4.5005
R69251 VINN.n356 VINN.n197 4.5005
R69252 VINN.n237 VINN.n197 4.5005
R69253 VINN.n358 VINN.n197 4.5005
R69254 VINN.n236 VINN.n197 4.5005
R69255 VINN.n360 VINN.n197 4.5005
R69256 VINN.n235 VINN.n197 4.5005
R69257 VINN.n362 VINN.n197 4.5005
R69258 VINN.n234 VINN.n197 4.5005
R69259 VINN.n364 VINN.n197 4.5005
R69260 VINN.n233 VINN.n197 4.5005
R69261 VINN.n366 VINN.n197 4.5005
R69262 VINN.n232 VINN.n197 4.5005
R69263 VINN.n368 VINN.n197 4.5005
R69264 VINN.n231 VINN.n197 4.5005
R69265 VINN.n370 VINN.n197 4.5005
R69266 VINN.n230 VINN.n197 4.5005
R69267 VINN.n372 VINN.n197 4.5005
R69268 VINN.n229 VINN.n197 4.5005
R69269 VINN.n374 VINN.n197 4.5005
R69270 VINN.n228 VINN.n197 4.5005
R69271 VINN.n376 VINN.n197 4.5005
R69272 VINN.n227 VINN.n197 4.5005
R69273 VINN.n378 VINN.n197 4.5005
R69274 VINN.n226 VINN.n197 4.5005
R69275 VINN.n380 VINN.n197 4.5005
R69276 VINN.n225 VINN.n197 4.5005
R69277 VINN.n382 VINN.n197 4.5005
R69278 VINN.n224 VINN.n197 4.5005
R69279 VINN.n384 VINN.n197 4.5005
R69280 VINN.n223 VINN.n197 4.5005
R69281 VINN.n386 VINN.n197 4.5005
R69282 VINN.n222 VINN.n197 4.5005
R69283 VINN.n388 VINN.n197 4.5005
R69284 VINN.n221 VINN.n197 4.5005
R69285 VINN.n390 VINN.n197 4.5005
R69286 VINN.n220 VINN.n197 4.5005
R69287 VINN.n392 VINN.n197 4.5005
R69288 VINN.n219 VINN.n197 4.5005
R69289 VINN.n394 VINN.n197 4.5005
R69290 VINN.n218 VINN.n197 4.5005
R69291 VINN.n396 VINN.n197 4.5005
R69292 VINN.n217 VINN.n197 4.5005
R69293 VINN.n398 VINN.n197 4.5005
R69294 VINN.n216 VINN.n197 4.5005
R69295 VINN.n400 VINN.n197 4.5005
R69296 VINN.n215 VINN.n197 4.5005
R69297 VINN.n654 VINN.n197 4.5005
R69298 VINN.n656 VINN.n197 4.5005
R69299 VINN.n197 VINN.n0 4.5005
R69300 VINN.n278 VINN.n103 4.5005
R69301 VINN.n276 VINN.n103 4.5005
R69302 VINN.n280 VINN.n103 4.5005
R69303 VINN.n275 VINN.n103 4.5005
R69304 VINN.n282 VINN.n103 4.5005
R69305 VINN.n274 VINN.n103 4.5005
R69306 VINN.n284 VINN.n103 4.5005
R69307 VINN.n273 VINN.n103 4.5005
R69308 VINN.n286 VINN.n103 4.5005
R69309 VINN.n272 VINN.n103 4.5005
R69310 VINN.n288 VINN.n103 4.5005
R69311 VINN.n271 VINN.n103 4.5005
R69312 VINN.n290 VINN.n103 4.5005
R69313 VINN.n270 VINN.n103 4.5005
R69314 VINN.n292 VINN.n103 4.5005
R69315 VINN.n269 VINN.n103 4.5005
R69316 VINN.n294 VINN.n103 4.5005
R69317 VINN.n268 VINN.n103 4.5005
R69318 VINN.n296 VINN.n103 4.5005
R69319 VINN.n267 VINN.n103 4.5005
R69320 VINN.n298 VINN.n103 4.5005
R69321 VINN.n266 VINN.n103 4.5005
R69322 VINN.n300 VINN.n103 4.5005
R69323 VINN.n265 VINN.n103 4.5005
R69324 VINN.n302 VINN.n103 4.5005
R69325 VINN.n264 VINN.n103 4.5005
R69326 VINN.n304 VINN.n103 4.5005
R69327 VINN.n263 VINN.n103 4.5005
R69328 VINN.n306 VINN.n103 4.5005
R69329 VINN.n262 VINN.n103 4.5005
R69330 VINN.n308 VINN.n103 4.5005
R69331 VINN.n261 VINN.n103 4.5005
R69332 VINN.n310 VINN.n103 4.5005
R69333 VINN.n260 VINN.n103 4.5005
R69334 VINN.n312 VINN.n103 4.5005
R69335 VINN.n259 VINN.n103 4.5005
R69336 VINN.n314 VINN.n103 4.5005
R69337 VINN.n258 VINN.n103 4.5005
R69338 VINN.n316 VINN.n103 4.5005
R69339 VINN.n257 VINN.n103 4.5005
R69340 VINN.n318 VINN.n103 4.5005
R69341 VINN.n256 VINN.n103 4.5005
R69342 VINN.n320 VINN.n103 4.5005
R69343 VINN.n255 VINN.n103 4.5005
R69344 VINN.n322 VINN.n103 4.5005
R69345 VINN.n254 VINN.n103 4.5005
R69346 VINN.n324 VINN.n103 4.5005
R69347 VINN.n253 VINN.n103 4.5005
R69348 VINN.n326 VINN.n103 4.5005
R69349 VINN.n252 VINN.n103 4.5005
R69350 VINN.n328 VINN.n103 4.5005
R69351 VINN.n251 VINN.n103 4.5005
R69352 VINN.n330 VINN.n103 4.5005
R69353 VINN.n250 VINN.n103 4.5005
R69354 VINN.n332 VINN.n103 4.5005
R69355 VINN.n249 VINN.n103 4.5005
R69356 VINN.n334 VINN.n103 4.5005
R69357 VINN.n248 VINN.n103 4.5005
R69358 VINN.n336 VINN.n103 4.5005
R69359 VINN.n247 VINN.n103 4.5005
R69360 VINN.n338 VINN.n103 4.5005
R69361 VINN.n246 VINN.n103 4.5005
R69362 VINN.n340 VINN.n103 4.5005
R69363 VINN.n245 VINN.n103 4.5005
R69364 VINN.n342 VINN.n103 4.5005
R69365 VINN.n244 VINN.n103 4.5005
R69366 VINN.n344 VINN.n103 4.5005
R69367 VINN.n243 VINN.n103 4.5005
R69368 VINN.n346 VINN.n103 4.5005
R69369 VINN.n242 VINN.n103 4.5005
R69370 VINN.n348 VINN.n103 4.5005
R69371 VINN.n241 VINN.n103 4.5005
R69372 VINN.n350 VINN.n103 4.5005
R69373 VINN.n240 VINN.n103 4.5005
R69374 VINN.n352 VINN.n103 4.5005
R69375 VINN.n239 VINN.n103 4.5005
R69376 VINN.n354 VINN.n103 4.5005
R69377 VINN.n238 VINN.n103 4.5005
R69378 VINN.n356 VINN.n103 4.5005
R69379 VINN.n237 VINN.n103 4.5005
R69380 VINN.n358 VINN.n103 4.5005
R69381 VINN.n236 VINN.n103 4.5005
R69382 VINN.n360 VINN.n103 4.5005
R69383 VINN.n235 VINN.n103 4.5005
R69384 VINN.n362 VINN.n103 4.5005
R69385 VINN.n234 VINN.n103 4.5005
R69386 VINN.n364 VINN.n103 4.5005
R69387 VINN.n233 VINN.n103 4.5005
R69388 VINN.n366 VINN.n103 4.5005
R69389 VINN.n232 VINN.n103 4.5005
R69390 VINN.n368 VINN.n103 4.5005
R69391 VINN.n231 VINN.n103 4.5005
R69392 VINN.n370 VINN.n103 4.5005
R69393 VINN.n230 VINN.n103 4.5005
R69394 VINN.n372 VINN.n103 4.5005
R69395 VINN.n229 VINN.n103 4.5005
R69396 VINN.n374 VINN.n103 4.5005
R69397 VINN.n228 VINN.n103 4.5005
R69398 VINN.n376 VINN.n103 4.5005
R69399 VINN.n227 VINN.n103 4.5005
R69400 VINN.n378 VINN.n103 4.5005
R69401 VINN.n226 VINN.n103 4.5005
R69402 VINN.n380 VINN.n103 4.5005
R69403 VINN.n225 VINN.n103 4.5005
R69404 VINN.n382 VINN.n103 4.5005
R69405 VINN.n224 VINN.n103 4.5005
R69406 VINN.n384 VINN.n103 4.5005
R69407 VINN.n223 VINN.n103 4.5005
R69408 VINN.n386 VINN.n103 4.5005
R69409 VINN.n222 VINN.n103 4.5005
R69410 VINN.n388 VINN.n103 4.5005
R69411 VINN.n221 VINN.n103 4.5005
R69412 VINN.n390 VINN.n103 4.5005
R69413 VINN.n220 VINN.n103 4.5005
R69414 VINN.n392 VINN.n103 4.5005
R69415 VINN.n219 VINN.n103 4.5005
R69416 VINN.n394 VINN.n103 4.5005
R69417 VINN.n218 VINN.n103 4.5005
R69418 VINN.n396 VINN.n103 4.5005
R69419 VINN.n217 VINN.n103 4.5005
R69420 VINN.n398 VINN.n103 4.5005
R69421 VINN.n216 VINN.n103 4.5005
R69422 VINN.n400 VINN.n103 4.5005
R69423 VINN.n215 VINN.n103 4.5005
R69424 VINN.n654 VINN.n103 4.5005
R69425 VINN.n656 VINN.n103 4.5005
R69426 VINN.n103 VINN.n0 4.5005
R69427 VINN.n278 VINN.n198 4.5005
R69428 VINN.n276 VINN.n198 4.5005
R69429 VINN.n280 VINN.n198 4.5005
R69430 VINN.n275 VINN.n198 4.5005
R69431 VINN.n282 VINN.n198 4.5005
R69432 VINN.n274 VINN.n198 4.5005
R69433 VINN.n284 VINN.n198 4.5005
R69434 VINN.n273 VINN.n198 4.5005
R69435 VINN.n286 VINN.n198 4.5005
R69436 VINN.n272 VINN.n198 4.5005
R69437 VINN.n288 VINN.n198 4.5005
R69438 VINN.n271 VINN.n198 4.5005
R69439 VINN.n290 VINN.n198 4.5005
R69440 VINN.n270 VINN.n198 4.5005
R69441 VINN.n292 VINN.n198 4.5005
R69442 VINN.n269 VINN.n198 4.5005
R69443 VINN.n294 VINN.n198 4.5005
R69444 VINN.n268 VINN.n198 4.5005
R69445 VINN.n296 VINN.n198 4.5005
R69446 VINN.n267 VINN.n198 4.5005
R69447 VINN.n298 VINN.n198 4.5005
R69448 VINN.n266 VINN.n198 4.5005
R69449 VINN.n300 VINN.n198 4.5005
R69450 VINN.n265 VINN.n198 4.5005
R69451 VINN.n302 VINN.n198 4.5005
R69452 VINN.n264 VINN.n198 4.5005
R69453 VINN.n304 VINN.n198 4.5005
R69454 VINN.n263 VINN.n198 4.5005
R69455 VINN.n306 VINN.n198 4.5005
R69456 VINN.n262 VINN.n198 4.5005
R69457 VINN.n308 VINN.n198 4.5005
R69458 VINN.n261 VINN.n198 4.5005
R69459 VINN.n310 VINN.n198 4.5005
R69460 VINN.n260 VINN.n198 4.5005
R69461 VINN.n312 VINN.n198 4.5005
R69462 VINN.n259 VINN.n198 4.5005
R69463 VINN.n314 VINN.n198 4.5005
R69464 VINN.n258 VINN.n198 4.5005
R69465 VINN.n316 VINN.n198 4.5005
R69466 VINN.n257 VINN.n198 4.5005
R69467 VINN.n318 VINN.n198 4.5005
R69468 VINN.n256 VINN.n198 4.5005
R69469 VINN.n320 VINN.n198 4.5005
R69470 VINN.n255 VINN.n198 4.5005
R69471 VINN.n322 VINN.n198 4.5005
R69472 VINN.n254 VINN.n198 4.5005
R69473 VINN.n324 VINN.n198 4.5005
R69474 VINN.n253 VINN.n198 4.5005
R69475 VINN.n326 VINN.n198 4.5005
R69476 VINN.n252 VINN.n198 4.5005
R69477 VINN.n328 VINN.n198 4.5005
R69478 VINN.n251 VINN.n198 4.5005
R69479 VINN.n330 VINN.n198 4.5005
R69480 VINN.n250 VINN.n198 4.5005
R69481 VINN.n332 VINN.n198 4.5005
R69482 VINN.n249 VINN.n198 4.5005
R69483 VINN.n334 VINN.n198 4.5005
R69484 VINN.n248 VINN.n198 4.5005
R69485 VINN.n336 VINN.n198 4.5005
R69486 VINN.n247 VINN.n198 4.5005
R69487 VINN.n338 VINN.n198 4.5005
R69488 VINN.n246 VINN.n198 4.5005
R69489 VINN.n340 VINN.n198 4.5005
R69490 VINN.n245 VINN.n198 4.5005
R69491 VINN.n342 VINN.n198 4.5005
R69492 VINN.n244 VINN.n198 4.5005
R69493 VINN.n344 VINN.n198 4.5005
R69494 VINN.n243 VINN.n198 4.5005
R69495 VINN.n346 VINN.n198 4.5005
R69496 VINN.n242 VINN.n198 4.5005
R69497 VINN.n348 VINN.n198 4.5005
R69498 VINN.n241 VINN.n198 4.5005
R69499 VINN.n350 VINN.n198 4.5005
R69500 VINN.n240 VINN.n198 4.5005
R69501 VINN.n352 VINN.n198 4.5005
R69502 VINN.n239 VINN.n198 4.5005
R69503 VINN.n354 VINN.n198 4.5005
R69504 VINN.n238 VINN.n198 4.5005
R69505 VINN.n356 VINN.n198 4.5005
R69506 VINN.n237 VINN.n198 4.5005
R69507 VINN.n358 VINN.n198 4.5005
R69508 VINN.n236 VINN.n198 4.5005
R69509 VINN.n360 VINN.n198 4.5005
R69510 VINN.n235 VINN.n198 4.5005
R69511 VINN.n362 VINN.n198 4.5005
R69512 VINN.n234 VINN.n198 4.5005
R69513 VINN.n364 VINN.n198 4.5005
R69514 VINN.n233 VINN.n198 4.5005
R69515 VINN.n366 VINN.n198 4.5005
R69516 VINN.n232 VINN.n198 4.5005
R69517 VINN.n368 VINN.n198 4.5005
R69518 VINN.n231 VINN.n198 4.5005
R69519 VINN.n370 VINN.n198 4.5005
R69520 VINN.n230 VINN.n198 4.5005
R69521 VINN.n372 VINN.n198 4.5005
R69522 VINN.n229 VINN.n198 4.5005
R69523 VINN.n374 VINN.n198 4.5005
R69524 VINN.n228 VINN.n198 4.5005
R69525 VINN.n376 VINN.n198 4.5005
R69526 VINN.n227 VINN.n198 4.5005
R69527 VINN.n378 VINN.n198 4.5005
R69528 VINN.n226 VINN.n198 4.5005
R69529 VINN.n380 VINN.n198 4.5005
R69530 VINN.n225 VINN.n198 4.5005
R69531 VINN.n382 VINN.n198 4.5005
R69532 VINN.n224 VINN.n198 4.5005
R69533 VINN.n384 VINN.n198 4.5005
R69534 VINN.n223 VINN.n198 4.5005
R69535 VINN.n386 VINN.n198 4.5005
R69536 VINN.n222 VINN.n198 4.5005
R69537 VINN.n388 VINN.n198 4.5005
R69538 VINN.n221 VINN.n198 4.5005
R69539 VINN.n390 VINN.n198 4.5005
R69540 VINN.n220 VINN.n198 4.5005
R69541 VINN.n392 VINN.n198 4.5005
R69542 VINN.n219 VINN.n198 4.5005
R69543 VINN.n394 VINN.n198 4.5005
R69544 VINN.n218 VINN.n198 4.5005
R69545 VINN.n396 VINN.n198 4.5005
R69546 VINN.n217 VINN.n198 4.5005
R69547 VINN.n398 VINN.n198 4.5005
R69548 VINN.n216 VINN.n198 4.5005
R69549 VINN.n400 VINN.n198 4.5005
R69550 VINN.n215 VINN.n198 4.5005
R69551 VINN.n654 VINN.n198 4.5005
R69552 VINN.n656 VINN.n198 4.5005
R69553 VINN.n198 VINN.n0 4.5005
R69554 VINN.n278 VINN.n102 4.5005
R69555 VINN.n276 VINN.n102 4.5005
R69556 VINN.n280 VINN.n102 4.5005
R69557 VINN.n275 VINN.n102 4.5005
R69558 VINN.n282 VINN.n102 4.5005
R69559 VINN.n274 VINN.n102 4.5005
R69560 VINN.n284 VINN.n102 4.5005
R69561 VINN.n273 VINN.n102 4.5005
R69562 VINN.n286 VINN.n102 4.5005
R69563 VINN.n272 VINN.n102 4.5005
R69564 VINN.n288 VINN.n102 4.5005
R69565 VINN.n271 VINN.n102 4.5005
R69566 VINN.n290 VINN.n102 4.5005
R69567 VINN.n270 VINN.n102 4.5005
R69568 VINN.n292 VINN.n102 4.5005
R69569 VINN.n269 VINN.n102 4.5005
R69570 VINN.n294 VINN.n102 4.5005
R69571 VINN.n268 VINN.n102 4.5005
R69572 VINN.n296 VINN.n102 4.5005
R69573 VINN.n267 VINN.n102 4.5005
R69574 VINN.n298 VINN.n102 4.5005
R69575 VINN.n266 VINN.n102 4.5005
R69576 VINN.n300 VINN.n102 4.5005
R69577 VINN.n265 VINN.n102 4.5005
R69578 VINN.n302 VINN.n102 4.5005
R69579 VINN.n264 VINN.n102 4.5005
R69580 VINN.n304 VINN.n102 4.5005
R69581 VINN.n263 VINN.n102 4.5005
R69582 VINN.n306 VINN.n102 4.5005
R69583 VINN.n262 VINN.n102 4.5005
R69584 VINN.n308 VINN.n102 4.5005
R69585 VINN.n261 VINN.n102 4.5005
R69586 VINN.n310 VINN.n102 4.5005
R69587 VINN.n260 VINN.n102 4.5005
R69588 VINN.n312 VINN.n102 4.5005
R69589 VINN.n259 VINN.n102 4.5005
R69590 VINN.n314 VINN.n102 4.5005
R69591 VINN.n258 VINN.n102 4.5005
R69592 VINN.n316 VINN.n102 4.5005
R69593 VINN.n257 VINN.n102 4.5005
R69594 VINN.n318 VINN.n102 4.5005
R69595 VINN.n256 VINN.n102 4.5005
R69596 VINN.n320 VINN.n102 4.5005
R69597 VINN.n255 VINN.n102 4.5005
R69598 VINN.n322 VINN.n102 4.5005
R69599 VINN.n254 VINN.n102 4.5005
R69600 VINN.n324 VINN.n102 4.5005
R69601 VINN.n253 VINN.n102 4.5005
R69602 VINN.n326 VINN.n102 4.5005
R69603 VINN.n252 VINN.n102 4.5005
R69604 VINN.n328 VINN.n102 4.5005
R69605 VINN.n251 VINN.n102 4.5005
R69606 VINN.n330 VINN.n102 4.5005
R69607 VINN.n250 VINN.n102 4.5005
R69608 VINN.n332 VINN.n102 4.5005
R69609 VINN.n249 VINN.n102 4.5005
R69610 VINN.n334 VINN.n102 4.5005
R69611 VINN.n248 VINN.n102 4.5005
R69612 VINN.n336 VINN.n102 4.5005
R69613 VINN.n247 VINN.n102 4.5005
R69614 VINN.n338 VINN.n102 4.5005
R69615 VINN.n246 VINN.n102 4.5005
R69616 VINN.n340 VINN.n102 4.5005
R69617 VINN.n245 VINN.n102 4.5005
R69618 VINN.n342 VINN.n102 4.5005
R69619 VINN.n244 VINN.n102 4.5005
R69620 VINN.n344 VINN.n102 4.5005
R69621 VINN.n243 VINN.n102 4.5005
R69622 VINN.n346 VINN.n102 4.5005
R69623 VINN.n242 VINN.n102 4.5005
R69624 VINN.n348 VINN.n102 4.5005
R69625 VINN.n241 VINN.n102 4.5005
R69626 VINN.n350 VINN.n102 4.5005
R69627 VINN.n240 VINN.n102 4.5005
R69628 VINN.n352 VINN.n102 4.5005
R69629 VINN.n239 VINN.n102 4.5005
R69630 VINN.n354 VINN.n102 4.5005
R69631 VINN.n238 VINN.n102 4.5005
R69632 VINN.n356 VINN.n102 4.5005
R69633 VINN.n237 VINN.n102 4.5005
R69634 VINN.n358 VINN.n102 4.5005
R69635 VINN.n236 VINN.n102 4.5005
R69636 VINN.n360 VINN.n102 4.5005
R69637 VINN.n235 VINN.n102 4.5005
R69638 VINN.n362 VINN.n102 4.5005
R69639 VINN.n234 VINN.n102 4.5005
R69640 VINN.n364 VINN.n102 4.5005
R69641 VINN.n233 VINN.n102 4.5005
R69642 VINN.n366 VINN.n102 4.5005
R69643 VINN.n232 VINN.n102 4.5005
R69644 VINN.n368 VINN.n102 4.5005
R69645 VINN.n231 VINN.n102 4.5005
R69646 VINN.n370 VINN.n102 4.5005
R69647 VINN.n230 VINN.n102 4.5005
R69648 VINN.n372 VINN.n102 4.5005
R69649 VINN.n229 VINN.n102 4.5005
R69650 VINN.n374 VINN.n102 4.5005
R69651 VINN.n228 VINN.n102 4.5005
R69652 VINN.n376 VINN.n102 4.5005
R69653 VINN.n227 VINN.n102 4.5005
R69654 VINN.n378 VINN.n102 4.5005
R69655 VINN.n226 VINN.n102 4.5005
R69656 VINN.n380 VINN.n102 4.5005
R69657 VINN.n225 VINN.n102 4.5005
R69658 VINN.n382 VINN.n102 4.5005
R69659 VINN.n224 VINN.n102 4.5005
R69660 VINN.n384 VINN.n102 4.5005
R69661 VINN.n223 VINN.n102 4.5005
R69662 VINN.n386 VINN.n102 4.5005
R69663 VINN.n222 VINN.n102 4.5005
R69664 VINN.n388 VINN.n102 4.5005
R69665 VINN.n221 VINN.n102 4.5005
R69666 VINN.n390 VINN.n102 4.5005
R69667 VINN.n220 VINN.n102 4.5005
R69668 VINN.n392 VINN.n102 4.5005
R69669 VINN.n219 VINN.n102 4.5005
R69670 VINN.n394 VINN.n102 4.5005
R69671 VINN.n218 VINN.n102 4.5005
R69672 VINN.n396 VINN.n102 4.5005
R69673 VINN.n217 VINN.n102 4.5005
R69674 VINN.n398 VINN.n102 4.5005
R69675 VINN.n216 VINN.n102 4.5005
R69676 VINN.n400 VINN.n102 4.5005
R69677 VINN.n215 VINN.n102 4.5005
R69678 VINN.n654 VINN.n102 4.5005
R69679 VINN.n656 VINN.n102 4.5005
R69680 VINN.n102 VINN.n0 4.5005
R69681 VINN.n278 VINN.n199 4.5005
R69682 VINN.n276 VINN.n199 4.5005
R69683 VINN.n280 VINN.n199 4.5005
R69684 VINN.n275 VINN.n199 4.5005
R69685 VINN.n282 VINN.n199 4.5005
R69686 VINN.n274 VINN.n199 4.5005
R69687 VINN.n284 VINN.n199 4.5005
R69688 VINN.n273 VINN.n199 4.5005
R69689 VINN.n286 VINN.n199 4.5005
R69690 VINN.n272 VINN.n199 4.5005
R69691 VINN.n288 VINN.n199 4.5005
R69692 VINN.n271 VINN.n199 4.5005
R69693 VINN.n290 VINN.n199 4.5005
R69694 VINN.n270 VINN.n199 4.5005
R69695 VINN.n292 VINN.n199 4.5005
R69696 VINN.n269 VINN.n199 4.5005
R69697 VINN.n294 VINN.n199 4.5005
R69698 VINN.n268 VINN.n199 4.5005
R69699 VINN.n296 VINN.n199 4.5005
R69700 VINN.n267 VINN.n199 4.5005
R69701 VINN.n298 VINN.n199 4.5005
R69702 VINN.n266 VINN.n199 4.5005
R69703 VINN.n300 VINN.n199 4.5005
R69704 VINN.n265 VINN.n199 4.5005
R69705 VINN.n302 VINN.n199 4.5005
R69706 VINN.n264 VINN.n199 4.5005
R69707 VINN.n304 VINN.n199 4.5005
R69708 VINN.n263 VINN.n199 4.5005
R69709 VINN.n306 VINN.n199 4.5005
R69710 VINN.n262 VINN.n199 4.5005
R69711 VINN.n308 VINN.n199 4.5005
R69712 VINN.n261 VINN.n199 4.5005
R69713 VINN.n310 VINN.n199 4.5005
R69714 VINN.n260 VINN.n199 4.5005
R69715 VINN.n312 VINN.n199 4.5005
R69716 VINN.n259 VINN.n199 4.5005
R69717 VINN.n314 VINN.n199 4.5005
R69718 VINN.n258 VINN.n199 4.5005
R69719 VINN.n316 VINN.n199 4.5005
R69720 VINN.n257 VINN.n199 4.5005
R69721 VINN.n318 VINN.n199 4.5005
R69722 VINN.n256 VINN.n199 4.5005
R69723 VINN.n320 VINN.n199 4.5005
R69724 VINN.n255 VINN.n199 4.5005
R69725 VINN.n322 VINN.n199 4.5005
R69726 VINN.n254 VINN.n199 4.5005
R69727 VINN.n324 VINN.n199 4.5005
R69728 VINN.n253 VINN.n199 4.5005
R69729 VINN.n326 VINN.n199 4.5005
R69730 VINN.n252 VINN.n199 4.5005
R69731 VINN.n328 VINN.n199 4.5005
R69732 VINN.n251 VINN.n199 4.5005
R69733 VINN.n330 VINN.n199 4.5005
R69734 VINN.n250 VINN.n199 4.5005
R69735 VINN.n332 VINN.n199 4.5005
R69736 VINN.n249 VINN.n199 4.5005
R69737 VINN.n334 VINN.n199 4.5005
R69738 VINN.n248 VINN.n199 4.5005
R69739 VINN.n336 VINN.n199 4.5005
R69740 VINN.n247 VINN.n199 4.5005
R69741 VINN.n338 VINN.n199 4.5005
R69742 VINN.n246 VINN.n199 4.5005
R69743 VINN.n340 VINN.n199 4.5005
R69744 VINN.n245 VINN.n199 4.5005
R69745 VINN.n342 VINN.n199 4.5005
R69746 VINN.n244 VINN.n199 4.5005
R69747 VINN.n344 VINN.n199 4.5005
R69748 VINN.n243 VINN.n199 4.5005
R69749 VINN.n346 VINN.n199 4.5005
R69750 VINN.n242 VINN.n199 4.5005
R69751 VINN.n348 VINN.n199 4.5005
R69752 VINN.n241 VINN.n199 4.5005
R69753 VINN.n350 VINN.n199 4.5005
R69754 VINN.n240 VINN.n199 4.5005
R69755 VINN.n352 VINN.n199 4.5005
R69756 VINN.n239 VINN.n199 4.5005
R69757 VINN.n354 VINN.n199 4.5005
R69758 VINN.n238 VINN.n199 4.5005
R69759 VINN.n356 VINN.n199 4.5005
R69760 VINN.n237 VINN.n199 4.5005
R69761 VINN.n358 VINN.n199 4.5005
R69762 VINN.n236 VINN.n199 4.5005
R69763 VINN.n360 VINN.n199 4.5005
R69764 VINN.n235 VINN.n199 4.5005
R69765 VINN.n362 VINN.n199 4.5005
R69766 VINN.n234 VINN.n199 4.5005
R69767 VINN.n364 VINN.n199 4.5005
R69768 VINN.n233 VINN.n199 4.5005
R69769 VINN.n366 VINN.n199 4.5005
R69770 VINN.n232 VINN.n199 4.5005
R69771 VINN.n368 VINN.n199 4.5005
R69772 VINN.n231 VINN.n199 4.5005
R69773 VINN.n370 VINN.n199 4.5005
R69774 VINN.n230 VINN.n199 4.5005
R69775 VINN.n372 VINN.n199 4.5005
R69776 VINN.n229 VINN.n199 4.5005
R69777 VINN.n374 VINN.n199 4.5005
R69778 VINN.n228 VINN.n199 4.5005
R69779 VINN.n376 VINN.n199 4.5005
R69780 VINN.n227 VINN.n199 4.5005
R69781 VINN.n378 VINN.n199 4.5005
R69782 VINN.n226 VINN.n199 4.5005
R69783 VINN.n380 VINN.n199 4.5005
R69784 VINN.n225 VINN.n199 4.5005
R69785 VINN.n382 VINN.n199 4.5005
R69786 VINN.n224 VINN.n199 4.5005
R69787 VINN.n384 VINN.n199 4.5005
R69788 VINN.n223 VINN.n199 4.5005
R69789 VINN.n386 VINN.n199 4.5005
R69790 VINN.n222 VINN.n199 4.5005
R69791 VINN.n388 VINN.n199 4.5005
R69792 VINN.n221 VINN.n199 4.5005
R69793 VINN.n390 VINN.n199 4.5005
R69794 VINN.n220 VINN.n199 4.5005
R69795 VINN.n392 VINN.n199 4.5005
R69796 VINN.n219 VINN.n199 4.5005
R69797 VINN.n394 VINN.n199 4.5005
R69798 VINN.n218 VINN.n199 4.5005
R69799 VINN.n396 VINN.n199 4.5005
R69800 VINN.n217 VINN.n199 4.5005
R69801 VINN.n398 VINN.n199 4.5005
R69802 VINN.n216 VINN.n199 4.5005
R69803 VINN.n400 VINN.n199 4.5005
R69804 VINN.n215 VINN.n199 4.5005
R69805 VINN.n654 VINN.n199 4.5005
R69806 VINN.n656 VINN.n199 4.5005
R69807 VINN.n199 VINN.n0 4.5005
R69808 VINN.n278 VINN.n101 4.5005
R69809 VINN.n276 VINN.n101 4.5005
R69810 VINN.n280 VINN.n101 4.5005
R69811 VINN.n275 VINN.n101 4.5005
R69812 VINN.n282 VINN.n101 4.5005
R69813 VINN.n274 VINN.n101 4.5005
R69814 VINN.n284 VINN.n101 4.5005
R69815 VINN.n273 VINN.n101 4.5005
R69816 VINN.n286 VINN.n101 4.5005
R69817 VINN.n272 VINN.n101 4.5005
R69818 VINN.n288 VINN.n101 4.5005
R69819 VINN.n271 VINN.n101 4.5005
R69820 VINN.n290 VINN.n101 4.5005
R69821 VINN.n270 VINN.n101 4.5005
R69822 VINN.n292 VINN.n101 4.5005
R69823 VINN.n269 VINN.n101 4.5005
R69824 VINN.n294 VINN.n101 4.5005
R69825 VINN.n268 VINN.n101 4.5005
R69826 VINN.n296 VINN.n101 4.5005
R69827 VINN.n267 VINN.n101 4.5005
R69828 VINN.n298 VINN.n101 4.5005
R69829 VINN.n266 VINN.n101 4.5005
R69830 VINN.n300 VINN.n101 4.5005
R69831 VINN.n265 VINN.n101 4.5005
R69832 VINN.n302 VINN.n101 4.5005
R69833 VINN.n264 VINN.n101 4.5005
R69834 VINN.n304 VINN.n101 4.5005
R69835 VINN.n263 VINN.n101 4.5005
R69836 VINN.n306 VINN.n101 4.5005
R69837 VINN.n262 VINN.n101 4.5005
R69838 VINN.n308 VINN.n101 4.5005
R69839 VINN.n261 VINN.n101 4.5005
R69840 VINN.n310 VINN.n101 4.5005
R69841 VINN.n260 VINN.n101 4.5005
R69842 VINN.n312 VINN.n101 4.5005
R69843 VINN.n259 VINN.n101 4.5005
R69844 VINN.n314 VINN.n101 4.5005
R69845 VINN.n258 VINN.n101 4.5005
R69846 VINN.n316 VINN.n101 4.5005
R69847 VINN.n257 VINN.n101 4.5005
R69848 VINN.n318 VINN.n101 4.5005
R69849 VINN.n256 VINN.n101 4.5005
R69850 VINN.n320 VINN.n101 4.5005
R69851 VINN.n255 VINN.n101 4.5005
R69852 VINN.n322 VINN.n101 4.5005
R69853 VINN.n254 VINN.n101 4.5005
R69854 VINN.n324 VINN.n101 4.5005
R69855 VINN.n253 VINN.n101 4.5005
R69856 VINN.n326 VINN.n101 4.5005
R69857 VINN.n252 VINN.n101 4.5005
R69858 VINN.n328 VINN.n101 4.5005
R69859 VINN.n251 VINN.n101 4.5005
R69860 VINN.n330 VINN.n101 4.5005
R69861 VINN.n250 VINN.n101 4.5005
R69862 VINN.n332 VINN.n101 4.5005
R69863 VINN.n249 VINN.n101 4.5005
R69864 VINN.n334 VINN.n101 4.5005
R69865 VINN.n248 VINN.n101 4.5005
R69866 VINN.n336 VINN.n101 4.5005
R69867 VINN.n247 VINN.n101 4.5005
R69868 VINN.n338 VINN.n101 4.5005
R69869 VINN.n246 VINN.n101 4.5005
R69870 VINN.n340 VINN.n101 4.5005
R69871 VINN.n245 VINN.n101 4.5005
R69872 VINN.n342 VINN.n101 4.5005
R69873 VINN.n244 VINN.n101 4.5005
R69874 VINN.n344 VINN.n101 4.5005
R69875 VINN.n243 VINN.n101 4.5005
R69876 VINN.n346 VINN.n101 4.5005
R69877 VINN.n242 VINN.n101 4.5005
R69878 VINN.n348 VINN.n101 4.5005
R69879 VINN.n241 VINN.n101 4.5005
R69880 VINN.n350 VINN.n101 4.5005
R69881 VINN.n240 VINN.n101 4.5005
R69882 VINN.n352 VINN.n101 4.5005
R69883 VINN.n239 VINN.n101 4.5005
R69884 VINN.n354 VINN.n101 4.5005
R69885 VINN.n238 VINN.n101 4.5005
R69886 VINN.n356 VINN.n101 4.5005
R69887 VINN.n237 VINN.n101 4.5005
R69888 VINN.n358 VINN.n101 4.5005
R69889 VINN.n236 VINN.n101 4.5005
R69890 VINN.n360 VINN.n101 4.5005
R69891 VINN.n235 VINN.n101 4.5005
R69892 VINN.n362 VINN.n101 4.5005
R69893 VINN.n234 VINN.n101 4.5005
R69894 VINN.n364 VINN.n101 4.5005
R69895 VINN.n233 VINN.n101 4.5005
R69896 VINN.n366 VINN.n101 4.5005
R69897 VINN.n232 VINN.n101 4.5005
R69898 VINN.n368 VINN.n101 4.5005
R69899 VINN.n231 VINN.n101 4.5005
R69900 VINN.n370 VINN.n101 4.5005
R69901 VINN.n230 VINN.n101 4.5005
R69902 VINN.n372 VINN.n101 4.5005
R69903 VINN.n229 VINN.n101 4.5005
R69904 VINN.n374 VINN.n101 4.5005
R69905 VINN.n228 VINN.n101 4.5005
R69906 VINN.n376 VINN.n101 4.5005
R69907 VINN.n227 VINN.n101 4.5005
R69908 VINN.n378 VINN.n101 4.5005
R69909 VINN.n226 VINN.n101 4.5005
R69910 VINN.n380 VINN.n101 4.5005
R69911 VINN.n225 VINN.n101 4.5005
R69912 VINN.n382 VINN.n101 4.5005
R69913 VINN.n224 VINN.n101 4.5005
R69914 VINN.n384 VINN.n101 4.5005
R69915 VINN.n223 VINN.n101 4.5005
R69916 VINN.n386 VINN.n101 4.5005
R69917 VINN.n222 VINN.n101 4.5005
R69918 VINN.n388 VINN.n101 4.5005
R69919 VINN.n221 VINN.n101 4.5005
R69920 VINN.n390 VINN.n101 4.5005
R69921 VINN.n220 VINN.n101 4.5005
R69922 VINN.n392 VINN.n101 4.5005
R69923 VINN.n219 VINN.n101 4.5005
R69924 VINN.n394 VINN.n101 4.5005
R69925 VINN.n218 VINN.n101 4.5005
R69926 VINN.n396 VINN.n101 4.5005
R69927 VINN.n217 VINN.n101 4.5005
R69928 VINN.n398 VINN.n101 4.5005
R69929 VINN.n216 VINN.n101 4.5005
R69930 VINN.n400 VINN.n101 4.5005
R69931 VINN.n215 VINN.n101 4.5005
R69932 VINN.n654 VINN.n101 4.5005
R69933 VINN.n656 VINN.n101 4.5005
R69934 VINN.n101 VINN.n0 4.5005
R69935 VINN.n278 VINN.n200 4.5005
R69936 VINN.n276 VINN.n200 4.5005
R69937 VINN.n280 VINN.n200 4.5005
R69938 VINN.n275 VINN.n200 4.5005
R69939 VINN.n282 VINN.n200 4.5005
R69940 VINN.n274 VINN.n200 4.5005
R69941 VINN.n284 VINN.n200 4.5005
R69942 VINN.n273 VINN.n200 4.5005
R69943 VINN.n286 VINN.n200 4.5005
R69944 VINN.n272 VINN.n200 4.5005
R69945 VINN.n288 VINN.n200 4.5005
R69946 VINN.n271 VINN.n200 4.5005
R69947 VINN.n290 VINN.n200 4.5005
R69948 VINN.n270 VINN.n200 4.5005
R69949 VINN.n292 VINN.n200 4.5005
R69950 VINN.n269 VINN.n200 4.5005
R69951 VINN.n294 VINN.n200 4.5005
R69952 VINN.n268 VINN.n200 4.5005
R69953 VINN.n296 VINN.n200 4.5005
R69954 VINN.n267 VINN.n200 4.5005
R69955 VINN.n298 VINN.n200 4.5005
R69956 VINN.n266 VINN.n200 4.5005
R69957 VINN.n300 VINN.n200 4.5005
R69958 VINN.n265 VINN.n200 4.5005
R69959 VINN.n302 VINN.n200 4.5005
R69960 VINN.n264 VINN.n200 4.5005
R69961 VINN.n304 VINN.n200 4.5005
R69962 VINN.n263 VINN.n200 4.5005
R69963 VINN.n306 VINN.n200 4.5005
R69964 VINN.n262 VINN.n200 4.5005
R69965 VINN.n308 VINN.n200 4.5005
R69966 VINN.n261 VINN.n200 4.5005
R69967 VINN.n310 VINN.n200 4.5005
R69968 VINN.n260 VINN.n200 4.5005
R69969 VINN.n312 VINN.n200 4.5005
R69970 VINN.n259 VINN.n200 4.5005
R69971 VINN.n314 VINN.n200 4.5005
R69972 VINN.n258 VINN.n200 4.5005
R69973 VINN.n316 VINN.n200 4.5005
R69974 VINN.n257 VINN.n200 4.5005
R69975 VINN.n318 VINN.n200 4.5005
R69976 VINN.n256 VINN.n200 4.5005
R69977 VINN.n320 VINN.n200 4.5005
R69978 VINN.n255 VINN.n200 4.5005
R69979 VINN.n322 VINN.n200 4.5005
R69980 VINN.n254 VINN.n200 4.5005
R69981 VINN.n324 VINN.n200 4.5005
R69982 VINN.n253 VINN.n200 4.5005
R69983 VINN.n326 VINN.n200 4.5005
R69984 VINN.n252 VINN.n200 4.5005
R69985 VINN.n328 VINN.n200 4.5005
R69986 VINN.n251 VINN.n200 4.5005
R69987 VINN.n330 VINN.n200 4.5005
R69988 VINN.n250 VINN.n200 4.5005
R69989 VINN.n332 VINN.n200 4.5005
R69990 VINN.n249 VINN.n200 4.5005
R69991 VINN.n334 VINN.n200 4.5005
R69992 VINN.n248 VINN.n200 4.5005
R69993 VINN.n336 VINN.n200 4.5005
R69994 VINN.n247 VINN.n200 4.5005
R69995 VINN.n338 VINN.n200 4.5005
R69996 VINN.n246 VINN.n200 4.5005
R69997 VINN.n340 VINN.n200 4.5005
R69998 VINN.n245 VINN.n200 4.5005
R69999 VINN.n342 VINN.n200 4.5005
R70000 VINN.n244 VINN.n200 4.5005
R70001 VINN.n344 VINN.n200 4.5005
R70002 VINN.n243 VINN.n200 4.5005
R70003 VINN.n346 VINN.n200 4.5005
R70004 VINN.n242 VINN.n200 4.5005
R70005 VINN.n348 VINN.n200 4.5005
R70006 VINN.n241 VINN.n200 4.5005
R70007 VINN.n350 VINN.n200 4.5005
R70008 VINN.n240 VINN.n200 4.5005
R70009 VINN.n352 VINN.n200 4.5005
R70010 VINN.n239 VINN.n200 4.5005
R70011 VINN.n354 VINN.n200 4.5005
R70012 VINN.n238 VINN.n200 4.5005
R70013 VINN.n356 VINN.n200 4.5005
R70014 VINN.n237 VINN.n200 4.5005
R70015 VINN.n358 VINN.n200 4.5005
R70016 VINN.n236 VINN.n200 4.5005
R70017 VINN.n360 VINN.n200 4.5005
R70018 VINN.n235 VINN.n200 4.5005
R70019 VINN.n362 VINN.n200 4.5005
R70020 VINN.n234 VINN.n200 4.5005
R70021 VINN.n364 VINN.n200 4.5005
R70022 VINN.n233 VINN.n200 4.5005
R70023 VINN.n366 VINN.n200 4.5005
R70024 VINN.n232 VINN.n200 4.5005
R70025 VINN.n368 VINN.n200 4.5005
R70026 VINN.n231 VINN.n200 4.5005
R70027 VINN.n370 VINN.n200 4.5005
R70028 VINN.n230 VINN.n200 4.5005
R70029 VINN.n372 VINN.n200 4.5005
R70030 VINN.n229 VINN.n200 4.5005
R70031 VINN.n374 VINN.n200 4.5005
R70032 VINN.n228 VINN.n200 4.5005
R70033 VINN.n376 VINN.n200 4.5005
R70034 VINN.n227 VINN.n200 4.5005
R70035 VINN.n378 VINN.n200 4.5005
R70036 VINN.n226 VINN.n200 4.5005
R70037 VINN.n380 VINN.n200 4.5005
R70038 VINN.n225 VINN.n200 4.5005
R70039 VINN.n382 VINN.n200 4.5005
R70040 VINN.n224 VINN.n200 4.5005
R70041 VINN.n384 VINN.n200 4.5005
R70042 VINN.n223 VINN.n200 4.5005
R70043 VINN.n386 VINN.n200 4.5005
R70044 VINN.n222 VINN.n200 4.5005
R70045 VINN.n388 VINN.n200 4.5005
R70046 VINN.n221 VINN.n200 4.5005
R70047 VINN.n390 VINN.n200 4.5005
R70048 VINN.n220 VINN.n200 4.5005
R70049 VINN.n392 VINN.n200 4.5005
R70050 VINN.n219 VINN.n200 4.5005
R70051 VINN.n394 VINN.n200 4.5005
R70052 VINN.n218 VINN.n200 4.5005
R70053 VINN.n396 VINN.n200 4.5005
R70054 VINN.n217 VINN.n200 4.5005
R70055 VINN.n398 VINN.n200 4.5005
R70056 VINN.n216 VINN.n200 4.5005
R70057 VINN.n400 VINN.n200 4.5005
R70058 VINN.n215 VINN.n200 4.5005
R70059 VINN.n654 VINN.n200 4.5005
R70060 VINN.n656 VINN.n200 4.5005
R70061 VINN.n200 VINN.n0 4.5005
R70062 VINN.n278 VINN.n100 4.5005
R70063 VINN.n276 VINN.n100 4.5005
R70064 VINN.n280 VINN.n100 4.5005
R70065 VINN.n275 VINN.n100 4.5005
R70066 VINN.n282 VINN.n100 4.5005
R70067 VINN.n274 VINN.n100 4.5005
R70068 VINN.n284 VINN.n100 4.5005
R70069 VINN.n273 VINN.n100 4.5005
R70070 VINN.n286 VINN.n100 4.5005
R70071 VINN.n272 VINN.n100 4.5005
R70072 VINN.n288 VINN.n100 4.5005
R70073 VINN.n271 VINN.n100 4.5005
R70074 VINN.n290 VINN.n100 4.5005
R70075 VINN.n270 VINN.n100 4.5005
R70076 VINN.n292 VINN.n100 4.5005
R70077 VINN.n269 VINN.n100 4.5005
R70078 VINN.n294 VINN.n100 4.5005
R70079 VINN.n268 VINN.n100 4.5005
R70080 VINN.n296 VINN.n100 4.5005
R70081 VINN.n267 VINN.n100 4.5005
R70082 VINN.n298 VINN.n100 4.5005
R70083 VINN.n266 VINN.n100 4.5005
R70084 VINN.n300 VINN.n100 4.5005
R70085 VINN.n265 VINN.n100 4.5005
R70086 VINN.n302 VINN.n100 4.5005
R70087 VINN.n264 VINN.n100 4.5005
R70088 VINN.n304 VINN.n100 4.5005
R70089 VINN.n263 VINN.n100 4.5005
R70090 VINN.n306 VINN.n100 4.5005
R70091 VINN.n262 VINN.n100 4.5005
R70092 VINN.n308 VINN.n100 4.5005
R70093 VINN.n261 VINN.n100 4.5005
R70094 VINN.n310 VINN.n100 4.5005
R70095 VINN.n260 VINN.n100 4.5005
R70096 VINN.n312 VINN.n100 4.5005
R70097 VINN.n259 VINN.n100 4.5005
R70098 VINN.n314 VINN.n100 4.5005
R70099 VINN.n258 VINN.n100 4.5005
R70100 VINN.n316 VINN.n100 4.5005
R70101 VINN.n257 VINN.n100 4.5005
R70102 VINN.n318 VINN.n100 4.5005
R70103 VINN.n256 VINN.n100 4.5005
R70104 VINN.n320 VINN.n100 4.5005
R70105 VINN.n255 VINN.n100 4.5005
R70106 VINN.n322 VINN.n100 4.5005
R70107 VINN.n254 VINN.n100 4.5005
R70108 VINN.n324 VINN.n100 4.5005
R70109 VINN.n253 VINN.n100 4.5005
R70110 VINN.n326 VINN.n100 4.5005
R70111 VINN.n252 VINN.n100 4.5005
R70112 VINN.n328 VINN.n100 4.5005
R70113 VINN.n251 VINN.n100 4.5005
R70114 VINN.n330 VINN.n100 4.5005
R70115 VINN.n250 VINN.n100 4.5005
R70116 VINN.n332 VINN.n100 4.5005
R70117 VINN.n249 VINN.n100 4.5005
R70118 VINN.n334 VINN.n100 4.5005
R70119 VINN.n248 VINN.n100 4.5005
R70120 VINN.n336 VINN.n100 4.5005
R70121 VINN.n247 VINN.n100 4.5005
R70122 VINN.n338 VINN.n100 4.5005
R70123 VINN.n246 VINN.n100 4.5005
R70124 VINN.n340 VINN.n100 4.5005
R70125 VINN.n245 VINN.n100 4.5005
R70126 VINN.n342 VINN.n100 4.5005
R70127 VINN.n244 VINN.n100 4.5005
R70128 VINN.n344 VINN.n100 4.5005
R70129 VINN.n243 VINN.n100 4.5005
R70130 VINN.n346 VINN.n100 4.5005
R70131 VINN.n242 VINN.n100 4.5005
R70132 VINN.n348 VINN.n100 4.5005
R70133 VINN.n241 VINN.n100 4.5005
R70134 VINN.n350 VINN.n100 4.5005
R70135 VINN.n240 VINN.n100 4.5005
R70136 VINN.n352 VINN.n100 4.5005
R70137 VINN.n239 VINN.n100 4.5005
R70138 VINN.n354 VINN.n100 4.5005
R70139 VINN.n238 VINN.n100 4.5005
R70140 VINN.n356 VINN.n100 4.5005
R70141 VINN.n237 VINN.n100 4.5005
R70142 VINN.n358 VINN.n100 4.5005
R70143 VINN.n236 VINN.n100 4.5005
R70144 VINN.n360 VINN.n100 4.5005
R70145 VINN.n235 VINN.n100 4.5005
R70146 VINN.n362 VINN.n100 4.5005
R70147 VINN.n234 VINN.n100 4.5005
R70148 VINN.n364 VINN.n100 4.5005
R70149 VINN.n233 VINN.n100 4.5005
R70150 VINN.n366 VINN.n100 4.5005
R70151 VINN.n232 VINN.n100 4.5005
R70152 VINN.n368 VINN.n100 4.5005
R70153 VINN.n231 VINN.n100 4.5005
R70154 VINN.n370 VINN.n100 4.5005
R70155 VINN.n230 VINN.n100 4.5005
R70156 VINN.n372 VINN.n100 4.5005
R70157 VINN.n229 VINN.n100 4.5005
R70158 VINN.n374 VINN.n100 4.5005
R70159 VINN.n228 VINN.n100 4.5005
R70160 VINN.n376 VINN.n100 4.5005
R70161 VINN.n227 VINN.n100 4.5005
R70162 VINN.n378 VINN.n100 4.5005
R70163 VINN.n226 VINN.n100 4.5005
R70164 VINN.n380 VINN.n100 4.5005
R70165 VINN.n225 VINN.n100 4.5005
R70166 VINN.n382 VINN.n100 4.5005
R70167 VINN.n224 VINN.n100 4.5005
R70168 VINN.n384 VINN.n100 4.5005
R70169 VINN.n223 VINN.n100 4.5005
R70170 VINN.n386 VINN.n100 4.5005
R70171 VINN.n222 VINN.n100 4.5005
R70172 VINN.n388 VINN.n100 4.5005
R70173 VINN.n221 VINN.n100 4.5005
R70174 VINN.n390 VINN.n100 4.5005
R70175 VINN.n220 VINN.n100 4.5005
R70176 VINN.n392 VINN.n100 4.5005
R70177 VINN.n219 VINN.n100 4.5005
R70178 VINN.n394 VINN.n100 4.5005
R70179 VINN.n218 VINN.n100 4.5005
R70180 VINN.n396 VINN.n100 4.5005
R70181 VINN.n217 VINN.n100 4.5005
R70182 VINN.n398 VINN.n100 4.5005
R70183 VINN.n216 VINN.n100 4.5005
R70184 VINN.n400 VINN.n100 4.5005
R70185 VINN.n215 VINN.n100 4.5005
R70186 VINN.n654 VINN.n100 4.5005
R70187 VINN.n656 VINN.n100 4.5005
R70188 VINN.n100 VINN.n0 4.5005
R70189 VINN.n278 VINN.n201 4.5005
R70190 VINN.n276 VINN.n201 4.5005
R70191 VINN.n280 VINN.n201 4.5005
R70192 VINN.n275 VINN.n201 4.5005
R70193 VINN.n282 VINN.n201 4.5005
R70194 VINN.n274 VINN.n201 4.5005
R70195 VINN.n284 VINN.n201 4.5005
R70196 VINN.n273 VINN.n201 4.5005
R70197 VINN.n286 VINN.n201 4.5005
R70198 VINN.n272 VINN.n201 4.5005
R70199 VINN.n288 VINN.n201 4.5005
R70200 VINN.n271 VINN.n201 4.5005
R70201 VINN.n290 VINN.n201 4.5005
R70202 VINN.n270 VINN.n201 4.5005
R70203 VINN.n292 VINN.n201 4.5005
R70204 VINN.n269 VINN.n201 4.5005
R70205 VINN.n294 VINN.n201 4.5005
R70206 VINN.n268 VINN.n201 4.5005
R70207 VINN.n296 VINN.n201 4.5005
R70208 VINN.n267 VINN.n201 4.5005
R70209 VINN.n298 VINN.n201 4.5005
R70210 VINN.n266 VINN.n201 4.5005
R70211 VINN.n300 VINN.n201 4.5005
R70212 VINN.n265 VINN.n201 4.5005
R70213 VINN.n302 VINN.n201 4.5005
R70214 VINN.n264 VINN.n201 4.5005
R70215 VINN.n304 VINN.n201 4.5005
R70216 VINN.n263 VINN.n201 4.5005
R70217 VINN.n306 VINN.n201 4.5005
R70218 VINN.n262 VINN.n201 4.5005
R70219 VINN.n308 VINN.n201 4.5005
R70220 VINN.n261 VINN.n201 4.5005
R70221 VINN.n310 VINN.n201 4.5005
R70222 VINN.n260 VINN.n201 4.5005
R70223 VINN.n312 VINN.n201 4.5005
R70224 VINN.n259 VINN.n201 4.5005
R70225 VINN.n314 VINN.n201 4.5005
R70226 VINN.n258 VINN.n201 4.5005
R70227 VINN.n316 VINN.n201 4.5005
R70228 VINN.n257 VINN.n201 4.5005
R70229 VINN.n318 VINN.n201 4.5005
R70230 VINN.n256 VINN.n201 4.5005
R70231 VINN.n320 VINN.n201 4.5005
R70232 VINN.n255 VINN.n201 4.5005
R70233 VINN.n322 VINN.n201 4.5005
R70234 VINN.n254 VINN.n201 4.5005
R70235 VINN.n324 VINN.n201 4.5005
R70236 VINN.n253 VINN.n201 4.5005
R70237 VINN.n326 VINN.n201 4.5005
R70238 VINN.n252 VINN.n201 4.5005
R70239 VINN.n328 VINN.n201 4.5005
R70240 VINN.n251 VINN.n201 4.5005
R70241 VINN.n330 VINN.n201 4.5005
R70242 VINN.n250 VINN.n201 4.5005
R70243 VINN.n332 VINN.n201 4.5005
R70244 VINN.n249 VINN.n201 4.5005
R70245 VINN.n334 VINN.n201 4.5005
R70246 VINN.n248 VINN.n201 4.5005
R70247 VINN.n336 VINN.n201 4.5005
R70248 VINN.n247 VINN.n201 4.5005
R70249 VINN.n338 VINN.n201 4.5005
R70250 VINN.n246 VINN.n201 4.5005
R70251 VINN.n340 VINN.n201 4.5005
R70252 VINN.n245 VINN.n201 4.5005
R70253 VINN.n342 VINN.n201 4.5005
R70254 VINN.n244 VINN.n201 4.5005
R70255 VINN.n344 VINN.n201 4.5005
R70256 VINN.n243 VINN.n201 4.5005
R70257 VINN.n346 VINN.n201 4.5005
R70258 VINN.n242 VINN.n201 4.5005
R70259 VINN.n348 VINN.n201 4.5005
R70260 VINN.n241 VINN.n201 4.5005
R70261 VINN.n350 VINN.n201 4.5005
R70262 VINN.n240 VINN.n201 4.5005
R70263 VINN.n352 VINN.n201 4.5005
R70264 VINN.n239 VINN.n201 4.5005
R70265 VINN.n354 VINN.n201 4.5005
R70266 VINN.n238 VINN.n201 4.5005
R70267 VINN.n356 VINN.n201 4.5005
R70268 VINN.n237 VINN.n201 4.5005
R70269 VINN.n358 VINN.n201 4.5005
R70270 VINN.n236 VINN.n201 4.5005
R70271 VINN.n360 VINN.n201 4.5005
R70272 VINN.n235 VINN.n201 4.5005
R70273 VINN.n362 VINN.n201 4.5005
R70274 VINN.n234 VINN.n201 4.5005
R70275 VINN.n364 VINN.n201 4.5005
R70276 VINN.n233 VINN.n201 4.5005
R70277 VINN.n366 VINN.n201 4.5005
R70278 VINN.n232 VINN.n201 4.5005
R70279 VINN.n368 VINN.n201 4.5005
R70280 VINN.n231 VINN.n201 4.5005
R70281 VINN.n370 VINN.n201 4.5005
R70282 VINN.n230 VINN.n201 4.5005
R70283 VINN.n372 VINN.n201 4.5005
R70284 VINN.n229 VINN.n201 4.5005
R70285 VINN.n374 VINN.n201 4.5005
R70286 VINN.n228 VINN.n201 4.5005
R70287 VINN.n376 VINN.n201 4.5005
R70288 VINN.n227 VINN.n201 4.5005
R70289 VINN.n378 VINN.n201 4.5005
R70290 VINN.n226 VINN.n201 4.5005
R70291 VINN.n380 VINN.n201 4.5005
R70292 VINN.n225 VINN.n201 4.5005
R70293 VINN.n382 VINN.n201 4.5005
R70294 VINN.n224 VINN.n201 4.5005
R70295 VINN.n384 VINN.n201 4.5005
R70296 VINN.n223 VINN.n201 4.5005
R70297 VINN.n386 VINN.n201 4.5005
R70298 VINN.n222 VINN.n201 4.5005
R70299 VINN.n388 VINN.n201 4.5005
R70300 VINN.n221 VINN.n201 4.5005
R70301 VINN.n390 VINN.n201 4.5005
R70302 VINN.n220 VINN.n201 4.5005
R70303 VINN.n392 VINN.n201 4.5005
R70304 VINN.n219 VINN.n201 4.5005
R70305 VINN.n394 VINN.n201 4.5005
R70306 VINN.n218 VINN.n201 4.5005
R70307 VINN.n396 VINN.n201 4.5005
R70308 VINN.n217 VINN.n201 4.5005
R70309 VINN.n398 VINN.n201 4.5005
R70310 VINN.n216 VINN.n201 4.5005
R70311 VINN.n400 VINN.n201 4.5005
R70312 VINN.n215 VINN.n201 4.5005
R70313 VINN.n654 VINN.n201 4.5005
R70314 VINN.n656 VINN.n201 4.5005
R70315 VINN.n201 VINN.n0 4.5005
R70316 VINN.n278 VINN.n99 4.5005
R70317 VINN.n276 VINN.n99 4.5005
R70318 VINN.n280 VINN.n99 4.5005
R70319 VINN.n275 VINN.n99 4.5005
R70320 VINN.n282 VINN.n99 4.5005
R70321 VINN.n274 VINN.n99 4.5005
R70322 VINN.n284 VINN.n99 4.5005
R70323 VINN.n273 VINN.n99 4.5005
R70324 VINN.n286 VINN.n99 4.5005
R70325 VINN.n272 VINN.n99 4.5005
R70326 VINN.n288 VINN.n99 4.5005
R70327 VINN.n271 VINN.n99 4.5005
R70328 VINN.n290 VINN.n99 4.5005
R70329 VINN.n270 VINN.n99 4.5005
R70330 VINN.n292 VINN.n99 4.5005
R70331 VINN.n269 VINN.n99 4.5005
R70332 VINN.n294 VINN.n99 4.5005
R70333 VINN.n268 VINN.n99 4.5005
R70334 VINN.n296 VINN.n99 4.5005
R70335 VINN.n267 VINN.n99 4.5005
R70336 VINN.n298 VINN.n99 4.5005
R70337 VINN.n266 VINN.n99 4.5005
R70338 VINN.n300 VINN.n99 4.5005
R70339 VINN.n265 VINN.n99 4.5005
R70340 VINN.n302 VINN.n99 4.5005
R70341 VINN.n264 VINN.n99 4.5005
R70342 VINN.n304 VINN.n99 4.5005
R70343 VINN.n263 VINN.n99 4.5005
R70344 VINN.n306 VINN.n99 4.5005
R70345 VINN.n262 VINN.n99 4.5005
R70346 VINN.n308 VINN.n99 4.5005
R70347 VINN.n261 VINN.n99 4.5005
R70348 VINN.n310 VINN.n99 4.5005
R70349 VINN.n260 VINN.n99 4.5005
R70350 VINN.n312 VINN.n99 4.5005
R70351 VINN.n259 VINN.n99 4.5005
R70352 VINN.n314 VINN.n99 4.5005
R70353 VINN.n258 VINN.n99 4.5005
R70354 VINN.n316 VINN.n99 4.5005
R70355 VINN.n257 VINN.n99 4.5005
R70356 VINN.n318 VINN.n99 4.5005
R70357 VINN.n256 VINN.n99 4.5005
R70358 VINN.n320 VINN.n99 4.5005
R70359 VINN.n255 VINN.n99 4.5005
R70360 VINN.n322 VINN.n99 4.5005
R70361 VINN.n254 VINN.n99 4.5005
R70362 VINN.n324 VINN.n99 4.5005
R70363 VINN.n253 VINN.n99 4.5005
R70364 VINN.n326 VINN.n99 4.5005
R70365 VINN.n252 VINN.n99 4.5005
R70366 VINN.n328 VINN.n99 4.5005
R70367 VINN.n251 VINN.n99 4.5005
R70368 VINN.n330 VINN.n99 4.5005
R70369 VINN.n250 VINN.n99 4.5005
R70370 VINN.n332 VINN.n99 4.5005
R70371 VINN.n249 VINN.n99 4.5005
R70372 VINN.n334 VINN.n99 4.5005
R70373 VINN.n248 VINN.n99 4.5005
R70374 VINN.n336 VINN.n99 4.5005
R70375 VINN.n247 VINN.n99 4.5005
R70376 VINN.n338 VINN.n99 4.5005
R70377 VINN.n246 VINN.n99 4.5005
R70378 VINN.n340 VINN.n99 4.5005
R70379 VINN.n245 VINN.n99 4.5005
R70380 VINN.n342 VINN.n99 4.5005
R70381 VINN.n244 VINN.n99 4.5005
R70382 VINN.n344 VINN.n99 4.5005
R70383 VINN.n243 VINN.n99 4.5005
R70384 VINN.n346 VINN.n99 4.5005
R70385 VINN.n242 VINN.n99 4.5005
R70386 VINN.n348 VINN.n99 4.5005
R70387 VINN.n241 VINN.n99 4.5005
R70388 VINN.n350 VINN.n99 4.5005
R70389 VINN.n240 VINN.n99 4.5005
R70390 VINN.n352 VINN.n99 4.5005
R70391 VINN.n239 VINN.n99 4.5005
R70392 VINN.n354 VINN.n99 4.5005
R70393 VINN.n238 VINN.n99 4.5005
R70394 VINN.n356 VINN.n99 4.5005
R70395 VINN.n237 VINN.n99 4.5005
R70396 VINN.n358 VINN.n99 4.5005
R70397 VINN.n236 VINN.n99 4.5005
R70398 VINN.n360 VINN.n99 4.5005
R70399 VINN.n235 VINN.n99 4.5005
R70400 VINN.n362 VINN.n99 4.5005
R70401 VINN.n234 VINN.n99 4.5005
R70402 VINN.n364 VINN.n99 4.5005
R70403 VINN.n233 VINN.n99 4.5005
R70404 VINN.n366 VINN.n99 4.5005
R70405 VINN.n232 VINN.n99 4.5005
R70406 VINN.n368 VINN.n99 4.5005
R70407 VINN.n231 VINN.n99 4.5005
R70408 VINN.n370 VINN.n99 4.5005
R70409 VINN.n230 VINN.n99 4.5005
R70410 VINN.n372 VINN.n99 4.5005
R70411 VINN.n229 VINN.n99 4.5005
R70412 VINN.n374 VINN.n99 4.5005
R70413 VINN.n228 VINN.n99 4.5005
R70414 VINN.n376 VINN.n99 4.5005
R70415 VINN.n227 VINN.n99 4.5005
R70416 VINN.n378 VINN.n99 4.5005
R70417 VINN.n226 VINN.n99 4.5005
R70418 VINN.n380 VINN.n99 4.5005
R70419 VINN.n225 VINN.n99 4.5005
R70420 VINN.n382 VINN.n99 4.5005
R70421 VINN.n224 VINN.n99 4.5005
R70422 VINN.n384 VINN.n99 4.5005
R70423 VINN.n223 VINN.n99 4.5005
R70424 VINN.n386 VINN.n99 4.5005
R70425 VINN.n222 VINN.n99 4.5005
R70426 VINN.n388 VINN.n99 4.5005
R70427 VINN.n221 VINN.n99 4.5005
R70428 VINN.n390 VINN.n99 4.5005
R70429 VINN.n220 VINN.n99 4.5005
R70430 VINN.n392 VINN.n99 4.5005
R70431 VINN.n219 VINN.n99 4.5005
R70432 VINN.n394 VINN.n99 4.5005
R70433 VINN.n218 VINN.n99 4.5005
R70434 VINN.n396 VINN.n99 4.5005
R70435 VINN.n217 VINN.n99 4.5005
R70436 VINN.n398 VINN.n99 4.5005
R70437 VINN.n216 VINN.n99 4.5005
R70438 VINN.n400 VINN.n99 4.5005
R70439 VINN.n215 VINN.n99 4.5005
R70440 VINN.n654 VINN.n99 4.5005
R70441 VINN.n656 VINN.n99 4.5005
R70442 VINN.n99 VINN.n0 4.5005
R70443 VINN.n278 VINN.n202 4.5005
R70444 VINN.n276 VINN.n202 4.5005
R70445 VINN.n280 VINN.n202 4.5005
R70446 VINN.n275 VINN.n202 4.5005
R70447 VINN.n282 VINN.n202 4.5005
R70448 VINN.n274 VINN.n202 4.5005
R70449 VINN.n284 VINN.n202 4.5005
R70450 VINN.n273 VINN.n202 4.5005
R70451 VINN.n286 VINN.n202 4.5005
R70452 VINN.n272 VINN.n202 4.5005
R70453 VINN.n288 VINN.n202 4.5005
R70454 VINN.n271 VINN.n202 4.5005
R70455 VINN.n290 VINN.n202 4.5005
R70456 VINN.n270 VINN.n202 4.5005
R70457 VINN.n292 VINN.n202 4.5005
R70458 VINN.n269 VINN.n202 4.5005
R70459 VINN.n294 VINN.n202 4.5005
R70460 VINN.n268 VINN.n202 4.5005
R70461 VINN.n296 VINN.n202 4.5005
R70462 VINN.n267 VINN.n202 4.5005
R70463 VINN.n298 VINN.n202 4.5005
R70464 VINN.n266 VINN.n202 4.5005
R70465 VINN.n300 VINN.n202 4.5005
R70466 VINN.n265 VINN.n202 4.5005
R70467 VINN.n302 VINN.n202 4.5005
R70468 VINN.n264 VINN.n202 4.5005
R70469 VINN.n304 VINN.n202 4.5005
R70470 VINN.n263 VINN.n202 4.5005
R70471 VINN.n306 VINN.n202 4.5005
R70472 VINN.n262 VINN.n202 4.5005
R70473 VINN.n308 VINN.n202 4.5005
R70474 VINN.n261 VINN.n202 4.5005
R70475 VINN.n310 VINN.n202 4.5005
R70476 VINN.n260 VINN.n202 4.5005
R70477 VINN.n312 VINN.n202 4.5005
R70478 VINN.n259 VINN.n202 4.5005
R70479 VINN.n314 VINN.n202 4.5005
R70480 VINN.n258 VINN.n202 4.5005
R70481 VINN.n316 VINN.n202 4.5005
R70482 VINN.n257 VINN.n202 4.5005
R70483 VINN.n318 VINN.n202 4.5005
R70484 VINN.n256 VINN.n202 4.5005
R70485 VINN.n320 VINN.n202 4.5005
R70486 VINN.n255 VINN.n202 4.5005
R70487 VINN.n322 VINN.n202 4.5005
R70488 VINN.n254 VINN.n202 4.5005
R70489 VINN.n324 VINN.n202 4.5005
R70490 VINN.n253 VINN.n202 4.5005
R70491 VINN.n326 VINN.n202 4.5005
R70492 VINN.n252 VINN.n202 4.5005
R70493 VINN.n328 VINN.n202 4.5005
R70494 VINN.n251 VINN.n202 4.5005
R70495 VINN.n330 VINN.n202 4.5005
R70496 VINN.n250 VINN.n202 4.5005
R70497 VINN.n332 VINN.n202 4.5005
R70498 VINN.n249 VINN.n202 4.5005
R70499 VINN.n334 VINN.n202 4.5005
R70500 VINN.n248 VINN.n202 4.5005
R70501 VINN.n336 VINN.n202 4.5005
R70502 VINN.n247 VINN.n202 4.5005
R70503 VINN.n338 VINN.n202 4.5005
R70504 VINN.n246 VINN.n202 4.5005
R70505 VINN.n340 VINN.n202 4.5005
R70506 VINN.n245 VINN.n202 4.5005
R70507 VINN.n342 VINN.n202 4.5005
R70508 VINN.n244 VINN.n202 4.5005
R70509 VINN.n344 VINN.n202 4.5005
R70510 VINN.n243 VINN.n202 4.5005
R70511 VINN.n346 VINN.n202 4.5005
R70512 VINN.n242 VINN.n202 4.5005
R70513 VINN.n348 VINN.n202 4.5005
R70514 VINN.n241 VINN.n202 4.5005
R70515 VINN.n350 VINN.n202 4.5005
R70516 VINN.n240 VINN.n202 4.5005
R70517 VINN.n352 VINN.n202 4.5005
R70518 VINN.n239 VINN.n202 4.5005
R70519 VINN.n354 VINN.n202 4.5005
R70520 VINN.n238 VINN.n202 4.5005
R70521 VINN.n356 VINN.n202 4.5005
R70522 VINN.n237 VINN.n202 4.5005
R70523 VINN.n358 VINN.n202 4.5005
R70524 VINN.n236 VINN.n202 4.5005
R70525 VINN.n360 VINN.n202 4.5005
R70526 VINN.n235 VINN.n202 4.5005
R70527 VINN.n362 VINN.n202 4.5005
R70528 VINN.n234 VINN.n202 4.5005
R70529 VINN.n364 VINN.n202 4.5005
R70530 VINN.n233 VINN.n202 4.5005
R70531 VINN.n366 VINN.n202 4.5005
R70532 VINN.n232 VINN.n202 4.5005
R70533 VINN.n368 VINN.n202 4.5005
R70534 VINN.n231 VINN.n202 4.5005
R70535 VINN.n370 VINN.n202 4.5005
R70536 VINN.n230 VINN.n202 4.5005
R70537 VINN.n372 VINN.n202 4.5005
R70538 VINN.n229 VINN.n202 4.5005
R70539 VINN.n374 VINN.n202 4.5005
R70540 VINN.n228 VINN.n202 4.5005
R70541 VINN.n376 VINN.n202 4.5005
R70542 VINN.n227 VINN.n202 4.5005
R70543 VINN.n378 VINN.n202 4.5005
R70544 VINN.n226 VINN.n202 4.5005
R70545 VINN.n380 VINN.n202 4.5005
R70546 VINN.n225 VINN.n202 4.5005
R70547 VINN.n382 VINN.n202 4.5005
R70548 VINN.n224 VINN.n202 4.5005
R70549 VINN.n384 VINN.n202 4.5005
R70550 VINN.n223 VINN.n202 4.5005
R70551 VINN.n386 VINN.n202 4.5005
R70552 VINN.n222 VINN.n202 4.5005
R70553 VINN.n388 VINN.n202 4.5005
R70554 VINN.n221 VINN.n202 4.5005
R70555 VINN.n390 VINN.n202 4.5005
R70556 VINN.n220 VINN.n202 4.5005
R70557 VINN.n392 VINN.n202 4.5005
R70558 VINN.n219 VINN.n202 4.5005
R70559 VINN.n394 VINN.n202 4.5005
R70560 VINN.n218 VINN.n202 4.5005
R70561 VINN.n396 VINN.n202 4.5005
R70562 VINN.n217 VINN.n202 4.5005
R70563 VINN.n398 VINN.n202 4.5005
R70564 VINN.n216 VINN.n202 4.5005
R70565 VINN.n400 VINN.n202 4.5005
R70566 VINN.n215 VINN.n202 4.5005
R70567 VINN.n654 VINN.n202 4.5005
R70568 VINN.n656 VINN.n202 4.5005
R70569 VINN.n202 VINN.n0 4.5005
R70570 VINN.n278 VINN.n98 4.5005
R70571 VINN.n276 VINN.n98 4.5005
R70572 VINN.n280 VINN.n98 4.5005
R70573 VINN.n275 VINN.n98 4.5005
R70574 VINN.n282 VINN.n98 4.5005
R70575 VINN.n274 VINN.n98 4.5005
R70576 VINN.n284 VINN.n98 4.5005
R70577 VINN.n273 VINN.n98 4.5005
R70578 VINN.n286 VINN.n98 4.5005
R70579 VINN.n272 VINN.n98 4.5005
R70580 VINN.n288 VINN.n98 4.5005
R70581 VINN.n271 VINN.n98 4.5005
R70582 VINN.n290 VINN.n98 4.5005
R70583 VINN.n270 VINN.n98 4.5005
R70584 VINN.n292 VINN.n98 4.5005
R70585 VINN.n269 VINN.n98 4.5005
R70586 VINN.n294 VINN.n98 4.5005
R70587 VINN.n268 VINN.n98 4.5005
R70588 VINN.n296 VINN.n98 4.5005
R70589 VINN.n267 VINN.n98 4.5005
R70590 VINN.n298 VINN.n98 4.5005
R70591 VINN.n266 VINN.n98 4.5005
R70592 VINN.n300 VINN.n98 4.5005
R70593 VINN.n265 VINN.n98 4.5005
R70594 VINN.n302 VINN.n98 4.5005
R70595 VINN.n264 VINN.n98 4.5005
R70596 VINN.n304 VINN.n98 4.5005
R70597 VINN.n263 VINN.n98 4.5005
R70598 VINN.n306 VINN.n98 4.5005
R70599 VINN.n262 VINN.n98 4.5005
R70600 VINN.n308 VINN.n98 4.5005
R70601 VINN.n261 VINN.n98 4.5005
R70602 VINN.n310 VINN.n98 4.5005
R70603 VINN.n260 VINN.n98 4.5005
R70604 VINN.n312 VINN.n98 4.5005
R70605 VINN.n259 VINN.n98 4.5005
R70606 VINN.n314 VINN.n98 4.5005
R70607 VINN.n258 VINN.n98 4.5005
R70608 VINN.n316 VINN.n98 4.5005
R70609 VINN.n257 VINN.n98 4.5005
R70610 VINN.n318 VINN.n98 4.5005
R70611 VINN.n256 VINN.n98 4.5005
R70612 VINN.n320 VINN.n98 4.5005
R70613 VINN.n255 VINN.n98 4.5005
R70614 VINN.n322 VINN.n98 4.5005
R70615 VINN.n254 VINN.n98 4.5005
R70616 VINN.n324 VINN.n98 4.5005
R70617 VINN.n253 VINN.n98 4.5005
R70618 VINN.n326 VINN.n98 4.5005
R70619 VINN.n252 VINN.n98 4.5005
R70620 VINN.n328 VINN.n98 4.5005
R70621 VINN.n251 VINN.n98 4.5005
R70622 VINN.n330 VINN.n98 4.5005
R70623 VINN.n250 VINN.n98 4.5005
R70624 VINN.n332 VINN.n98 4.5005
R70625 VINN.n249 VINN.n98 4.5005
R70626 VINN.n334 VINN.n98 4.5005
R70627 VINN.n248 VINN.n98 4.5005
R70628 VINN.n336 VINN.n98 4.5005
R70629 VINN.n247 VINN.n98 4.5005
R70630 VINN.n338 VINN.n98 4.5005
R70631 VINN.n246 VINN.n98 4.5005
R70632 VINN.n340 VINN.n98 4.5005
R70633 VINN.n245 VINN.n98 4.5005
R70634 VINN.n342 VINN.n98 4.5005
R70635 VINN.n244 VINN.n98 4.5005
R70636 VINN.n344 VINN.n98 4.5005
R70637 VINN.n243 VINN.n98 4.5005
R70638 VINN.n346 VINN.n98 4.5005
R70639 VINN.n242 VINN.n98 4.5005
R70640 VINN.n348 VINN.n98 4.5005
R70641 VINN.n241 VINN.n98 4.5005
R70642 VINN.n350 VINN.n98 4.5005
R70643 VINN.n240 VINN.n98 4.5005
R70644 VINN.n352 VINN.n98 4.5005
R70645 VINN.n239 VINN.n98 4.5005
R70646 VINN.n354 VINN.n98 4.5005
R70647 VINN.n238 VINN.n98 4.5005
R70648 VINN.n356 VINN.n98 4.5005
R70649 VINN.n237 VINN.n98 4.5005
R70650 VINN.n358 VINN.n98 4.5005
R70651 VINN.n236 VINN.n98 4.5005
R70652 VINN.n360 VINN.n98 4.5005
R70653 VINN.n235 VINN.n98 4.5005
R70654 VINN.n362 VINN.n98 4.5005
R70655 VINN.n234 VINN.n98 4.5005
R70656 VINN.n364 VINN.n98 4.5005
R70657 VINN.n233 VINN.n98 4.5005
R70658 VINN.n366 VINN.n98 4.5005
R70659 VINN.n232 VINN.n98 4.5005
R70660 VINN.n368 VINN.n98 4.5005
R70661 VINN.n231 VINN.n98 4.5005
R70662 VINN.n370 VINN.n98 4.5005
R70663 VINN.n230 VINN.n98 4.5005
R70664 VINN.n372 VINN.n98 4.5005
R70665 VINN.n229 VINN.n98 4.5005
R70666 VINN.n374 VINN.n98 4.5005
R70667 VINN.n228 VINN.n98 4.5005
R70668 VINN.n376 VINN.n98 4.5005
R70669 VINN.n227 VINN.n98 4.5005
R70670 VINN.n378 VINN.n98 4.5005
R70671 VINN.n226 VINN.n98 4.5005
R70672 VINN.n380 VINN.n98 4.5005
R70673 VINN.n225 VINN.n98 4.5005
R70674 VINN.n382 VINN.n98 4.5005
R70675 VINN.n224 VINN.n98 4.5005
R70676 VINN.n384 VINN.n98 4.5005
R70677 VINN.n223 VINN.n98 4.5005
R70678 VINN.n386 VINN.n98 4.5005
R70679 VINN.n222 VINN.n98 4.5005
R70680 VINN.n388 VINN.n98 4.5005
R70681 VINN.n221 VINN.n98 4.5005
R70682 VINN.n390 VINN.n98 4.5005
R70683 VINN.n220 VINN.n98 4.5005
R70684 VINN.n392 VINN.n98 4.5005
R70685 VINN.n219 VINN.n98 4.5005
R70686 VINN.n394 VINN.n98 4.5005
R70687 VINN.n218 VINN.n98 4.5005
R70688 VINN.n396 VINN.n98 4.5005
R70689 VINN.n217 VINN.n98 4.5005
R70690 VINN.n398 VINN.n98 4.5005
R70691 VINN.n216 VINN.n98 4.5005
R70692 VINN.n400 VINN.n98 4.5005
R70693 VINN.n215 VINN.n98 4.5005
R70694 VINN.n654 VINN.n98 4.5005
R70695 VINN.n656 VINN.n98 4.5005
R70696 VINN.n98 VINN.n0 4.5005
R70697 VINN.n278 VINN.n203 4.5005
R70698 VINN.n276 VINN.n203 4.5005
R70699 VINN.n280 VINN.n203 4.5005
R70700 VINN.n275 VINN.n203 4.5005
R70701 VINN.n282 VINN.n203 4.5005
R70702 VINN.n274 VINN.n203 4.5005
R70703 VINN.n284 VINN.n203 4.5005
R70704 VINN.n273 VINN.n203 4.5005
R70705 VINN.n286 VINN.n203 4.5005
R70706 VINN.n272 VINN.n203 4.5005
R70707 VINN.n288 VINN.n203 4.5005
R70708 VINN.n271 VINN.n203 4.5005
R70709 VINN.n290 VINN.n203 4.5005
R70710 VINN.n270 VINN.n203 4.5005
R70711 VINN.n292 VINN.n203 4.5005
R70712 VINN.n269 VINN.n203 4.5005
R70713 VINN.n294 VINN.n203 4.5005
R70714 VINN.n268 VINN.n203 4.5005
R70715 VINN.n296 VINN.n203 4.5005
R70716 VINN.n267 VINN.n203 4.5005
R70717 VINN.n298 VINN.n203 4.5005
R70718 VINN.n266 VINN.n203 4.5005
R70719 VINN.n300 VINN.n203 4.5005
R70720 VINN.n265 VINN.n203 4.5005
R70721 VINN.n302 VINN.n203 4.5005
R70722 VINN.n264 VINN.n203 4.5005
R70723 VINN.n304 VINN.n203 4.5005
R70724 VINN.n263 VINN.n203 4.5005
R70725 VINN.n306 VINN.n203 4.5005
R70726 VINN.n262 VINN.n203 4.5005
R70727 VINN.n308 VINN.n203 4.5005
R70728 VINN.n261 VINN.n203 4.5005
R70729 VINN.n310 VINN.n203 4.5005
R70730 VINN.n260 VINN.n203 4.5005
R70731 VINN.n312 VINN.n203 4.5005
R70732 VINN.n259 VINN.n203 4.5005
R70733 VINN.n314 VINN.n203 4.5005
R70734 VINN.n258 VINN.n203 4.5005
R70735 VINN.n316 VINN.n203 4.5005
R70736 VINN.n257 VINN.n203 4.5005
R70737 VINN.n318 VINN.n203 4.5005
R70738 VINN.n256 VINN.n203 4.5005
R70739 VINN.n320 VINN.n203 4.5005
R70740 VINN.n255 VINN.n203 4.5005
R70741 VINN.n322 VINN.n203 4.5005
R70742 VINN.n254 VINN.n203 4.5005
R70743 VINN.n324 VINN.n203 4.5005
R70744 VINN.n253 VINN.n203 4.5005
R70745 VINN.n326 VINN.n203 4.5005
R70746 VINN.n252 VINN.n203 4.5005
R70747 VINN.n328 VINN.n203 4.5005
R70748 VINN.n251 VINN.n203 4.5005
R70749 VINN.n330 VINN.n203 4.5005
R70750 VINN.n250 VINN.n203 4.5005
R70751 VINN.n332 VINN.n203 4.5005
R70752 VINN.n249 VINN.n203 4.5005
R70753 VINN.n334 VINN.n203 4.5005
R70754 VINN.n248 VINN.n203 4.5005
R70755 VINN.n336 VINN.n203 4.5005
R70756 VINN.n247 VINN.n203 4.5005
R70757 VINN.n338 VINN.n203 4.5005
R70758 VINN.n246 VINN.n203 4.5005
R70759 VINN.n340 VINN.n203 4.5005
R70760 VINN.n245 VINN.n203 4.5005
R70761 VINN.n342 VINN.n203 4.5005
R70762 VINN.n244 VINN.n203 4.5005
R70763 VINN.n344 VINN.n203 4.5005
R70764 VINN.n243 VINN.n203 4.5005
R70765 VINN.n346 VINN.n203 4.5005
R70766 VINN.n242 VINN.n203 4.5005
R70767 VINN.n348 VINN.n203 4.5005
R70768 VINN.n241 VINN.n203 4.5005
R70769 VINN.n350 VINN.n203 4.5005
R70770 VINN.n240 VINN.n203 4.5005
R70771 VINN.n352 VINN.n203 4.5005
R70772 VINN.n239 VINN.n203 4.5005
R70773 VINN.n354 VINN.n203 4.5005
R70774 VINN.n238 VINN.n203 4.5005
R70775 VINN.n356 VINN.n203 4.5005
R70776 VINN.n237 VINN.n203 4.5005
R70777 VINN.n358 VINN.n203 4.5005
R70778 VINN.n236 VINN.n203 4.5005
R70779 VINN.n360 VINN.n203 4.5005
R70780 VINN.n235 VINN.n203 4.5005
R70781 VINN.n362 VINN.n203 4.5005
R70782 VINN.n234 VINN.n203 4.5005
R70783 VINN.n364 VINN.n203 4.5005
R70784 VINN.n233 VINN.n203 4.5005
R70785 VINN.n366 VINN.n203 4.5005
R70786 VINN.n232 VINN.n203 4.5005
R70787 VINN.n368 VINN.n203 4.5005
R70788 VINN.n231 VINN.n203 4.5005
R70789 VINN.n370 VINN.n203 4.5005
R70790 VINN.n230 VINN.n203 4.5005
R70791 VINN.n372 VINN.n203 4.5005
R70792 VINN.n229 VINN.n203 4.5005
R70793 VINN.n374 VINN.n203 4.5005
R70794 VINN.n228 VINN.n203 4.5005
R70795 VINN.n376 VINN.n203 4.5005
R70796 VINN.n227 VINN.n203 4.5005
R70797 VINN.n378 VINN.n203 4.5005
R70798 VINN.n226 VINN.n203 4.5005
R70799 VINN.n380 VINN.n203 4.5005
R70800 VINN.n225 VINN.n203 4.5005
R70801 VINN.n382 VINN.n203 4.5005
R70802 VINN.n224 VINN.n203 4.5005
R70803 VINN.n384 VINN.n203 4.5005
R70804 VINN.n223 VINN.n203 4.5005
R70805 VINN.n386 VINN.n203 4.5005
R70806 VINN.n222 VINN.n203 4.5005
R70807 VINN.n388 VINN.n203 4.5005
R70808 VINN.n221 VINN.n203 4.5005
R70809 VINN.n390 VINN.n203 4.5005
R70810 VINN.n220 VINN.n203 4.5005
R70811 VINN.n392 VINN.n203 4.5005
R70812 VINN.n219 VINN.n203 4.5005
R70813 VINN.n394 VINN.n203 4.5005
R70814 VINN.n218 VINN.n203 4.5005
R70815 VINN.n396 VINN.n203 4.5005
R70816 VINN.n217 VINN.n203 4.5005
R70817 VINN.n398 VINN.n203 4.5005
R70818 VINN.n216 VINN.n203 4.5005
R70819 VINN.n400 VINN.n203 4.5005
R70820 VINN.n215 VINN.n203 4.5005
R70821 VINN.n654 VINN.n203 4.5005
R70822 VINN.n656 VINN.n203 4.5005
R70823 VINN.n203 VINN.n0 4.5005
R70824 VINN.n278 VINN.n97 4.5005
R70825 VINN.n276 VINN.n97 4.5005
R70826 VINN.n280 VINN.n97 4.5005
R70827 VINN.n275 VINN.n97 4.5005
R70828 VINN.n282 VINN.n97 4.5005
R70829 VINN.n274 VINN.n97 4.5005
R70830 VINN.n284 VINN.n97 4.5005
R70831 VINN.n273 VINN.n97 4.5005
R70832 VINN.n286 VINN.n97 4.5005
R70833 VINN.n272 VINN.n97 4.5005
R70834 VINN.n288 VINN.n97 4.5005
R70835 VINN.n271 VINN.n97 4.5005
R70836 VINN.n290 VINN.n97 4.5005
R70837 VINN.n270 VINN.n97 4.5005
R70838 VINN.n292 VINN.n97 4.5005
R70839 VINN.n269 VINN.n97 4.5005
R70840 VINN.n294 VINN.n97 4.5005
R70841 VINN.n268 VINN.n97 4.5005
R70842 VINN.n296 VINN.n97 4.5005
R70843 VINN.n267 VINN.n97 4.5005
R70844 VINN.n298 VINN.n97 4.5005
R70845 VINN.n266 VINN.n97 4.5005
R70846 VINN.n300 VINN.n97 4.5005
R70847 VINN.n265 VINN.n97 4.5005
R70848 VINN.n302 VINN.n97 4.5005
R70849 VINN.n264 VINN.n97 4.5005
R70850 VINN.n304 VINN.n97 4.5005
R70851 VINN.n263 VINN.n97 4.5005
R70852 VINN.n306 VINN.n97 4.5005
R70853 VINN.n262 VINN.n97 4.5005
R70854 VINN.n308 VINN.n97 4.5005
R70855 VINN.n261 VINN.n97 4.5005
R70856 VINN.n310 VINN.n97 4.5005
R70857 VINN.n260 VINN.n97 4.5005
R70858 VINN.n312 VINN.n97 4.5005
R70859 VINN.n259 VINN.n97 4.5005
R70860 VINN.n314 VINN.n97 4.5005
R70861 VINN.n258 VINN.n97 4.5005
R70862 VINN.n316 VINN.n97 4.5005
R70863 VINN.n257 VINN.n97 4.5005
R70864 VINN.n318 VINN.n97 4.5005
R70865 VINN.n256 VINN.n97 4.5005
R70866 VINN.n320 VINN.n97 4.5005
R70867 VINN.n255 VINN.n97 4.5005
R70868 VINN.n322 VINN.n97 4.5005
R70869 VINN.n254 VINN.n97 4.5005
R70870 VINN.n324 VINN.n97 4.5005
R70871 VINN.n253 VINN.n97 4.5005
R70872 VINN.n326 VINN.n97 4.5005
R70873 VINN.n252 VINN.n97 4.5005
R70874 VINN.n328 VINN.n97 4.5005
R70875 VINN.n251 VINN.n97 4.5005
R70876 VINN.n330 VINN.n97 4.5005
R70877 VINN.n250 VINN.n97 4.5005
R70878 VINN.n332 VINN.n97 4.5005
R70879 VINN.n249 VINN.n97 4.5005
R70880 VINN.n334 VINN.n97 4.5005
R70881 VINN.n248 VINN.n97 4.5005
R70882 VINN.n336 VINN.n97 4.5005
R70883 VINN.n247 VINN.n97 4.5005
R70884 VINN.n338 VINN.n97 4.5005
R70885 VINN.n246 VINN.n97 4.5005
R70886 VINN.n340 VINN.n97 4.5005
R70887 VINN.n245 VINN.n97 4.5005
R70888 VINN.n342 VINN.n97 4.5005
R70889 VINN.n244 VINN.n97 4.5005
R70890 VINN.n344 VINN.n97 4.5005
R70891 VINN.n243 VINN.n97 4.5005
R70892 VINN.n346 VINN.n97 4.5005
R70893 VINN.n242 VINN.n97 4.5005
R70894 VINN.n348 VINN.n97 4.5005
R70895 VINN.n241 VINN.n97 4.5005
R70896 VINN.n350 VINN.n97 4.5005
R70897 VINN.n240 VINN.n97 4.5005
R70898 VINN.n352 VINN.n97 4.5005
R70899 VINN.n239 VINN.n97 4.5005
R70900 VINN.n354 VINN.n97 4.5005
R70901 VINN.n238 VINN.n97 4.5005
R70902 VINN.n356 VINN.n97 4.5005
R70903 VINN.n237 VINN.n97 4.5005
R70904 VINN.n358 VINN.n97 4.5005
R70905 VINN.n236 VINN.n97 4.5005
R70906 VINN.n360 VINN.n97 4.5005
R70907 VINN.n235 VINN.n97 4.5005
R70908 VINN.n362 VINN.n97 4.5005
R70909 VINN.n234 VINN.n97 4.5005
R70910 VINN.n364 VINN.n97 4.5005
R70911 VINN.n233 VINN.n97 4.5005
R70912 VINN.n366 VINN.n97 4.5005
R70913 VINN.n232 VINN.n97 4.5005
R70914 VINN.n368 VINN.n97 4.5005
R70915 VINN.n231 VINN.n97 4.5005
R70916 VINN.n370 VINN.n97 4.5005
R70917 VINN.n230 VINN.n97 4.5005
R70918 VINN.n372 VINN.n97 4.5005
R70919 VINN.n229 VINN.n97 4.5005
R70920 VINN.n374 VINN.n97 4.5005
R70921 VINN.n228 VINN.n97 4.5005
R70922 VINN.n376 VINN.n97 4.5005
R70923 VINN.n227 VINN.n97 4.5005
R70924 VINN.n378 VINN.n97 4.5005
R70925 VINN.n226 VINN.n97 4.5005
R70926 VINN.n380 VINN.n97 4.5005
R70927 VINN.n225 VINN.n97 4.5005
R70928 VINN.n382 VINN.n97 4.5005
R70929 VINN.n224 VINN.n97 4.5005
R70930 VINN.n384 VINN.n97 4.5005
R70931 VINN.n223 VINN.n97 4.5005
R70932 VINN.n386 VINN.n97 4.5005
R70933 VINN.n222 VINN.n97 4.5005
R70934 VINN.n388 VINN.n97 4.5005
R70935 VINN.n221 VINN.n97 4.5005
R70936 VINN.n390 VINN.n97 4.5005
R70937 VINN.n220 VINN.n97 4.5005
R70938 VINN.n392 VINN.n97 4.5005
R70939 VINN.n219 VINN.n97 4.5005
R70940 VINN.n394 VINN.n97 4.5005
R70941 VINN.n218 VINN.n97 4.5005
R70942 VINN.n396 VINN.n97 4.5005
R70943 VINN.n217 VINN.n97 4.5005
R70944 VINN.n398 VINN.n97 4.5005
R70945 VINN.n216 VINN.n97 4.5005
R70946 VINN.n400 VINN.n97 4.5005
R70947 VINN.n215 VINN.n97 4.5005
R70948 VINN.n654 VINN.n97 4.5005
R70949 VINN.n656 VINN.n97 4.5005
R70950 VINN.n97 VINN.n0 4.5005
R70951 VINN.n278 VINN.n204 4.5005
R70952 VINN.n276 VINN.n204 4.5005
R70953 VINN.n280 VINN.n204 4.5005
R70954 VINN.n275 VINN.n204 4.5005
R70955 VINN.n282 VINN.n204 4.5005
R70956 VINN.n274 VINN.n204 4.5005
R70957 VINN.n284 VINN.n204 4.5005
R70958 VINN.n273 VINN.n204 4.5005
R70959 VINN.n286 VINN.n204 4.5005
R70960 VINN.n272 VINN.n204 4.5005
R70961 VINN.n288 VINN.n204 4.5005
R70962 VINN.n271 VINN.n204 4.5005
R70963 VINN.n290 VINN.n204 4.5005
R70964 VINN.n270 VINN.n204 4.5005
R70965 VINN.n292 VINN.n204 4.5005
R70966 VINN.n269 VINN.n204 4.5005
R70967 VINN.n294 VINN.n204 4.5005
R70968 VINN.n268 VINN.n204 4.5005
R70969 VINN.n296 VINN.n204 4.5005
R70970 VINN.n267 VINN.n204 4.5005
R70971 VINN.n298 VINN.n204 4.5005
R70972 VINN.n266 VINN.n204 4.5005
R70973 VINN.n300 VINN.n204 4.5005
R70974 VINN.n265 VINN.n204 4.5005
R70975 VINN.n302 VINN.n204 4.5005
R70976 VINN.n264 VINN.n204 4.5005
R70977 VINN.n304 VINN.n204 4.5005
R70978 VINN.n263 VINN.n204 4.5005
R70979 VINN.n306 VINN.n204 4.5005
R70980 VINN.n262 VINN.n204 4.5005
R70981 VINN.n308 VINN.n204 4.5005
R70982 VINN.n261 VINN.n204 4.5005
R70983 VINN.n310 VINN.n204 4.5005
R70984 VINN.n260 VINN.n204 4.5005
R70985 VINN.n312 VINN.n204 4.5005
R70986 VINN.n259 VINN.n204 4.5005
R70987 VINN.n314 VINN.n204 4.5005
R70988 VINN.n258 VINN.n204 4.5005
R70989 VINN.n316 VINN.n204 4.5005
R70990 VINN.n257 VINN.n204 4.5005
R70991 VINN.n318 VINN.n204 4.5005
R70992 VINN.n256 VINN.n204 4.5005
R70993 VINN.n320 VINN.n204 4.5005
R70994 VINN.n255 VINN.n204 4.5005
R70995 VINN.n322 VINN.n204 4.5005
R70996 VINN.n254 VINN.n204 4.5005
R70997 VINN.n324 VINN.n204 4.5005
R70998 VINN.n253 VINN.n204 4.5005
R70999 VINN.n326 VINN.n204 4.5005
R71000 VINN.n252 VINN.n204 4.5005
R71001 VINN.n328 VINN.n204 4.5005
R71002 VINN.n251 VINN.n204 4.5005
R71003 VINN.n330 VINN.n204 4.5005
R71004 VINN.n250 VINN.n204 4.5005
R71005 VINN.n332 VINN.n204 4.5005
R71006 VINN.n249 VINN.n204 4.5005
R71007 VINN.n334 VINN.n204 4.5005
R71008 VINN.n248 VINN.n204 4.5005
R71009 VINN.n336 VINN.n204 4.5005
R71010 VINN.n247 VINN.n204 4.5005
R71011 VINN.n338 VINN.n204 4.5005
R71012 VINN.n246 VINN.n204 4.5005
R71013 VINN.n340 VINN.n204 4.5005
R71014 VINN.n245 VINN.n204 4.5005
R71015 VINN.n342 VINN.n204 4.5005
R71016 VINN.n244 VINN.n204 4.5005
R71017 VINN.n344 VINN.n204 4.5005
R71018 VINN.n243 VINN.n204 4.5005
R71019 VINN.n346 VINN.n204 4.5005
R71020 VINN.n242 VINN.n204 4.5005
R71021 VINN.n348 VINN.n204 4.5005
R71022 VINN.n241 VINN.n204 4.5005
R71023 VINN.n350 VINN.n204 4.5005
R71024 VINN.n240 VINN.n204 4.5005
R71025 VINN.n352 VINN.n204 4.5005
R71026 VINN.n239 VINN.n204 4.5005
R71027 VINN.n354 VINN.n204 4.5005
R71028 VINN.n238 VINN.n204 4.5005
R71029 VINN.n356 VINN.n204 4.5005
R71030 VINN.n237 VINN.n204 4.5005
R71031 VINN.n358 VINN.n204 4.5005
R71032 VINN.n236 VINN.n204 4.5005
R71033 VINN.n360 VINN.n204 4.5005
R71034 VINN.n235 VINN.n204 4.5005
R71035 VINN.n362 VINN.n204 4.5005
R71036 VINN.n234 VINN.n204 4.5005
R71037 VINN.n364 VINN.n204 4.5005
R71038 VINN.n233 VINN.n204 4.5005
R71039 VINN.n366 VINN.n204 4.5005
R71040 VINN.n232 VINN.n204 4.5005
R71041 VINN.n368 VINN.n204 4.5005
R71042 VINN.n231 VINN.n204 4.5005
R71043 VINN.n370 VINN.n204 4.5005
R71044 VINN.n230 VINN.n204 4.5005
R71045 VINN.n372 VINN.n204 4.5005
R71046 VINN.n229 VINN.n204 4.5005
R71047 VINN.n374 VINN.n204 4.5005
R71048 VINN.n228 VINN.n204 4.5005
R71049 VINN.n376 VINN.n204 4.5005
R71050 VINN.n227 VINN.n204 4.5005
R71051 VINN.n378 VINN.n204 4.5005
R71052 VINN.n226 VINN.n204 4.5005
R71053 VINN.n380 VINN.n204 4.5005
R71054 VINN.n225 VINN.n204 4.5005
R71055 VINN.n382 VINN.n204 4.5005
R71056 VINN.n224 VINN.n204 4.5005
R71057 VINN.n384 VINN.n204 4.5005
R71058 VINN.n223 VINN.n204 4.5005
R71059 VINN.n386 VINN.n204 4.5005
R71060 VINN.n222 VINN.n204 4.5005
R71061 VINN.n388 VINN.n204 4.5005
R71062 VINN.n221 VINN.n204 4.5005
R71063 VINN.n390 VINN.n204 4.5005
R71064 VINN.n220 VINN.n204 4.5005
R71065 VINN.n392 VINN.n204 4.5005
R71066 VINN.n219 VINN.n204 4.5005
R71067 VINN.n394 VINN.n204 4.5005
R71068 VINN.n218 VINN.n204 4.5005
R71069 VINN.n396 VINN.n204 4.5005
R71070 VINN.n217 VINN.n204 4.5005
R71071 VINN.n398 VINN.n204 4.5005
R71072 VINN.n216 VINN.n204 4.5005
R71073 VINN.n400 VINN.n204 4.5005
R71074 VINN.n215 VINN.n204 4.5005
R71075 VINN.n654 VINN.n204 4.5005
R71076 VINN.n656 VINN.n204 4.5005
R71077 VINN.n204 VINN.n0 4.5005
R71078 VINN.n278 VINN.n96 4.5005
R71079 VINN.n276 VINN.n96 4.5005
R71080 VINN.n280 VINN.n96 4.5005
R71081 VINN.n275 VINN.n96 4.5005
R71082 VINN.n282 VINN.n96 4.5005
R71083 VINN.n274 VINN.n96 4.5005
R71084 VINN.n284 VINN.n96 4.5005
R71085 VINN.n273 VINN.n96 4.5005
R71086 VINN.n286 VINN.n96 4.5005
R71087 VINN.n272 VINN.n96 4.5005
R71088 VINN.n288 VINN.n96 4.5005
R71089 VINN.n271 VINN.n96 4.5005
R71090 VINN.n290 VINN.n96 4.5005
R71091 VINN.n270 VINN.n96 4.5005
R71092 VINN.n292 VINN.n96 4.5005
R71093 VINN.n269 VINN.n96 4.5005
R71094 VINN.n294 VINN.n96 4.5005
R71095 VINN.n268 VINN.n96 4.5005
R71096 VINN.n296 VINN.n96 4.5005
R71097 VINN.n267 VINN.n96 4.5005
R71098 VINN.n298 VINN.n96 4.5005
R71099 VINN.n266 VINN.n96 4.5005
R71100 VINN.n300 VINN.n96 4.5005
R71101 VINN.n265 VINN.n96 4.5005
R71102 VINN.n302 VINN.n96 4.5005
R71103 VINN.n264 VINN.n96 4.5005
R71104 VINN.n304 VINN.n96 4.5005
R71105 VINN.n263 VINN.n96 4.5005
R71106 VINN.n306 VINN.n96 4.5005
R71107 VINN.n262 VINN.n96 4.5005
R71108 VINN.n308 VINN.n96 4.5005
R71109 VINN.n261 VINN.n96 4.5005
R71110 VINN.n310 VINN.n96 4.5005
R71111 VINN.n260 VINN.n96 4.5005
R71112 VINN.n312 VINN.n96 4.5005
R71113 VINN.n259 VINN.n96 4.5005
R71114 VINN.n314 VINN.n96 4.5005
R71115 VINN.n258 VINN.n96 4.5005
R71116 VINN.n316 VINN.n96 4.5005
R71117 VINN.n257 VINN.n96 4.5005
R71118 VINN.n318 VINN.n96 4.5005
R71119 VINN.n256 VINN.n96 4.5005
R71120 VINN.n320 VINN.n96 4.5005
R71121 VINN.n255 VINN.n96 4.5005
R71122 VINN.n322 VINN.n96 4.5005
R71123 VINN.n254 VINN.n96 4.5005
R71124 VINN.n324 VINN.n96 4.5005
R71125 VINN.n253 VINN.n96 4.5005
R71126 VINN.n326 VINN.n96 4.5005
R71127 VINN.n252 VINN.n96 4.5005
R71128 VINN.n328 VINN.n96 4.5005
R71129 VINN.n251 VINN.n96 4.5005
R71130 VINN.n330 VINN.n96 4.5005
R71131 VINN.n250 VINN.n96 4.5005
R71132 VINN.n332 VINN.n96 4.5005
R71133 VINN.n249 VINN.n96 4.5005
R71134 VINN.n334 VINN.n96 4.5005
R71135 VINN.n248 VINN.n96 4.5005
R71136 VINN.n336 VINN.n96 4.5005
R71137 VINN.n247 VINN.n96 4.5005
R71138 VINN.n338 VINN.n96 4.5005
R71139 VINN.n246 VINN.n96 4.5005
R71140 VINN.n340 VINN.n96 4.5005
R71141 VINN.n245 VINN.n96 4.5005
R71142 VINN.n342 VINN.n96 4.5005
R71143 VINN.n244 VINN.n96 4.5005
R71144 VINN.n344 VINN.n96 4.5005
R71145 VINN.n243 VINN.n96 4.5005
R71146 VINN.n346 VINN.n96 4.5005
R71147 VINN.n242 VINN.n96 4.5005
R71148 VINN.n348 VINN.n96 4.5005
R71149 VINN.n241 VINN.n96 4.5005
R71150 VINN.n350 VINN.n96 4.5005
R71151 VINN.n240 VINN.n96 4.5005
R71152 VINN.n352 VINN.n96 4.5005
R71153 VINN.n239 VINN.n96 4.5005
R71154 VINN.n354 VINN.n96 4.5005
R71155 VINN.n238 VINN.n96 4.5005
R71156 VINN.n356 VINN.n96 4.5005
R71157 VINN.n237 VINN.n96 4.5005
R71158 VINN.n358 VINN.n96 4.5005
R71159 VINN.n236 VINN.n96 4.5005
R71160 VINN.n360 VINN.n96 4.5005
R71161 VINN.n235 VINN.n96 4.5005
R71162 VINN.n362 VINN.n96 4.5005
R71163 VINN.n234 VINN.n96 4.5005
R71164 VINN.n364 VINN.n96 4.5005
R71165 VINN.n233 VINN.n96 4.5005
R71166 VINN.n366 VINN.n96 4.5005
R71167 VINN.n232 VINN.n96 4.5005
R71168 VINN.n368 VINN.n96 4.5005
R71169 VINN.n231 VINN.n96 4.5005
R71170 VINN.n370 VINN.n96 4.5005
R71171 VINN.n230 VINN.n96 4.5005
R71172 VINN.n372 VINN.n96 4.5005
R71173 VINN.n229 VINN.n96 4.5005
R71174 VINN.n374 VINN.n96 4.5005
R71175 VINN.n228 VINN.n96 4.5005
R71176 VINN.n376 VINN.n96 4.5005
R71177 VINN.n227 VINN.n96 4.5005
R71178 VINN.n378 VINN.n96 4.5005
R71179 VINN.n226 VINN.n96 4.5005
R71180 VINN.n380 VINN.n96 4.5005
R71181 VINN.n225 VINN.n96 4.5005
R71182 VINN.n382 VINN.n96 4.5005
R71183 VINN.n224 VINN.n96 4.5005
R71184 VINN.n384 VINN.n96 4.5005
R71185 VINN.n223 VINN.n96 4.5005
R71186 VINN.n386 VINN.n96 4.5005
R71187 VINN.n222 VINN.n96 4.5005
R71188 VINN.n388 VINN.n96 4.5005
R71189 VINN.n221 VINN.n96 4.5005
R71190 VINN.n390 VINN.n96 4.5005
R71191 VINN.n220 VINN.n96 4.5005
R71192 VINN.n392 VINN.n96 4.5005
R71193 VINN.n219 VINN.n96 4.5005
R71194 VINN.n394 VINN.n96 4.5005
R71195 VINN.n218 VINN.n96 4.5005
R71196 VINN.n396 VINN.n96 4.5005
R71197 VINN.n217 VINN.n96 4.5005
R71198 VINN.n398 VINN.n96 4.5005
R71199 VINN.n216 VINN.n96 4.5005
R71200 VINN.n400 VINN.n96 4.5005
R71201 VINN.n215 VINN.n96 4.5005
R71202 VINN.n654 VINN.n96 4.5005
R71203 VINN.n656 VINN.n96 4.5005
R71204 VINN.n96 VINN.n0 4.5005
R71205 VINN.n278 VINN.n205 4.5005
R71206 VINN.n276 VINN.n205 4.5005
R71207 VINN.n280 VINN.n205 4.5005
R71208 VINN.n275 VINN.n205 4.5005
R71209 VINN.n282 VINN.n205 4.5005
R71210 VINN.n274 VINN.n205 4.5005
R71211 VINN.n284 VINN.n205 4.5005
R71212 VINN.n273 VINN.n205 4.5005
R71213 VINN.n286 VINN.n205 4.5005
R71214 VINN.n272 VINN.n205 4.5005
R71215 VINN.n288 VINN.n205 4.5005
R71216 VINN.n271 VINN.n205 4.5005
R71217 VINN.n290 VINN.n205 4.5005
R71218 VINN.n270 VINN.n205 4.5005
R71219 VINN.n292 VINN.n205 4.5005
R71220 VINN.n269 VINN.n205 4.5005
R71221 VINN.n294 VINN.n205 4.5005
R71222 VINN.n268 VINN.n205 4.5005
R71223 VINN.n296 VINN.n205 4.5005
R71224 VINN.n267 VINN.n205 4.5005
R71225 VINN.n298 VINN.n205 4.5005
R71226 VINN.n266 VINN.n205 4.5005
R71227 VINN.n300 VINN.n205 4.5005
R71228 VINN.n265 VINN.n205 4.5005
R71229 VINN.n302 VINN.n205 4.5005
R71230 VINN.n264 VINN.n205 4.5005
R71231 VINN.n304 VINN.n205 4.5005
R71232 VINN.n263 VINN.n205 4.5005
R71233 VINN.n306 VINN.n205 4.5005
R71234 VINN.n262 VINN.n205 4.5005
R71235 VINN.n308 VINN.n205 4.5005
R71236 VINN.n261 VINN.n205 4.5005
R71237 VINN.n310 VINN.n205 4.5005
R71238 VINN.n260 VINN.n205 4.5005
R71239 VINN.n312 VINN.n205 4.5005
R71240 VINN.n259 VINN.n205 4.5005
R71241 VINN.n314 VINN.n205 4.5005
R71242 VINN.n258 VINN.n205 4.5005
R71243 VINN.n316 VINN.n205 4.5005
R71244 VINN.n257 VINN.n205 4.5005
R71245 VINN.n318 VINN.n205 4.5005
R71246 VINN.n256 VINN.n205 4.5005
R71247 VINN.n320 VINN.n205 4.5005
R71248 VINN.n255 VINN.n205 4.5005
R71249 VINN.n322 VINN.n205 4.5005
R71250 VINN.n254 VINN.n205 4.5005
R71251 VINN.n324 VINN.n205 4.5005
R71252 VINN.n253 VINN.n205 4.5005
R71253 VINN.n326 VINN.n205 4.5005
R71254 VINN.n252 VINN.n205 4.5005
R71255 VINN.n328 VINN.n205 4.5005
R71256 VINN.n251 VINN.n205 4.5005
R71257 VINN.n330 VINN.n205 4.5005
R71258 VINN.n250 VINN.n205 4.5005
R71259 VINN.n332 VINN.n205 4.5005
R71260 VINN.n249 VINN.n205 4.5005
R71261 VINN.n334 VINN.n205 4.5005
R71262 VINN.n248 VINN.n205 4.5005
R71263 VINN.n336 VINN.n205 4.5005
R71264 VINN.n247 VINN.n205 4.5005
R71265 VINN.n338 VINN.n205 4.5005
R71266 VINN.n246 VINN.n205 4.5005
R71267 VINN.n340 VINN.n205 4.5005
R71268 VINN.n245 VINN.n205 4.5005
R71269 VINN.n342 VINN.n205 4.5005
R71270 VINN.n244 VINN.n205 4.5005
R71271 VINN.n344 VINN.n205 4.5005
R71272 VINN.n243 VINN.n205 4.5005
R71273 VINN.n346 VINN.n205 4.5005
R71274 VINN.n242 VINN.n205 4.5005
R71275 VINN.n348 VINN.n205 4.5005
R71276 VINN.n241 VINN.n205 4.5005
R71277 VINN.n350 VINN.n205 4.5005
R71278 VINN.n240 VINN.n205 4.5005
R71279 VINN.n352 VINN.n205 4.5005
R71280 VINN.n239 VINN.n205 4.5005
R71281 VINN.n354 VINN.n205 4.5005
R71282 VINN.n238 VINN.n205 4.5005
R71283 VINN.n356 VINN.n205 4.5005
R71284 VINN.n237 VINN.n205 4.5005
R71285 VINN.n358 VINN.n205 4.5005
R71286 VINN.n236 VINN.n205 4.5005
R71287 VINN.n360 VINN.n205 4.5005
R71288 VINN.n235 VINN.n205 4.5005
R71289 VINN.n362 VINN.n205 4.5005
R71290 VINN.n234 VINN.n205 4.5005
R71291 VINN.n364 VINN.n205 4.5005
R71292 VINN.n233 VINN.n205 4.5005
R71293 VINN.n366 VINN.n205 4.5005
R71294 VINN.n232 VINN.n205 4.5005
R71295 VINN.n368 VINN.n205 4.5005
R71296 VINN.n231 VINN.n205 4.5005
R71297 VINN.n370 VINN.n205 4.5005
R71298 VINN.n230 VINN.n205 4.5005
R71299 VINN.n372 VINN.n205 4.5005
R71300 VINN.n229 VINN.n205 4.5005
R71301 VINN.n374 VINN.n205 4.5005
R71302 VINN.n228 VINN.n205 4.5005
R71303 VINN.n376 VINN.n205 4.5005
R71304 VINN.n227 VINN.n205 4.5005
R71305 VINN.n378 VINN.n205 4.5005
R71306 VINN.n226 VINN.n205 4.5005
R71307 VINN.n380 VINN.n205 4.5005
R71308 VINN.n225 VINN.n205 4.5005
R71309 VINN.n382 VINN.n205 4.5005
R71310 VINN.n224 VINN.n205 4.5005
R71311 VINN.n384 VINN.n205 4.5005
R71312 VINN.n223 VINN.n205 4.5005
R71313 VINN.n386 VINN.n205 4.5005
R71314 VINN.n222 VINN.n205 4.5005
R71315 VINN.n388 VINN.n205 4.5005
R71316 VINN.n221 VINN.n205 4.5005
R71317 VINN.n390 VINN.n205 4.5005
R71318 VINN.n220 VINN.n205 4.5005
R71319 VINN.n392 VINN.n205 4.5005
R71320 VINN.n219 VINN.n205 4.5005
R71321 VINN.n394 VINN.n205 4.5005
R71322 VINN.n218 VINN.n205 4.5005
R71323 VINN.n396 VINN.n205 4.5005
R71324 VINN.n217 VINN.n205 4.5005
R71325 VINN.n398 VINN.n205 4.5005
R71326 VINN.n216 VINN.n205 4.5005
R71327 VINN.n400 VINN.n205 4.5005
R71328 VINN.n215 VINN.n205 4.5005
R71329 VINN.n654 VINN.n205 4.5005
R71330 VINN.n656 VINN.n205 4.5005
R71331 VINN.n205 VINN.n0 4.5005
R71332 VINN.n278 VINN.n95 4.5005
R71333 VINN.n276 VINN.n95 4.5005
R71334 VINN.n280 VINN.n95 4.5005
R71335 VINN.n275 VINN.n95 4.5005
R71336 VINN.n282 VINN.n95 4.5005
R71337 VINN.n274 VINN.n95 4.5005
R71338 VINN.n284 VINN.n95 4.5005
R71339 VINN.n273 VINN.n95 4.5005
R71340 VINN.n286 VINN.n95 4.5005
R71341 VINN.n272 VINN.n95 4.5005
R71342 VINN.n288 VINN.n95 4.5005
R71343 VINN.n271 VINN.n95 4.5005
R71344 VINN.n290 VINN.n95 4.5005
R71345 VINN.n270 VINN.n95 4.5005
R71346 VINN.n292 VINN.n95 4.5005
R71347 VINN.n269 VINN.n95 4.5005
R71348 VINN.n294 VINN.n95 4.5005
R71349 VINN.n268 VINN.n95 4.5005
R71350 VINN.n296 VINN.n95 4.5005
R71351 VINN.n267 VINN.n95 4.5005
R71352 VINN.n298 VINN.n95 4.5005
R71353 VINN.n266 VINN.n95 4.5005
R71354 VINN.n300 VINN.n95 4.5005
R71355 VINN.n265 VINN.n95 4.5005
R71356 VINN.n302 VINN.n95 4.5005
R71357 VINN.n264 VINN.n95 4.5005
R71358 VINN.n304 VINN.n95 4.5005
R71359 VINN.n263 VINN.n95 4.5005
R71360 VINN.n306 VINN.n95 4.5005
R71361 VINN.n262 VINN.n95 4.5005
R71362 VINN.n308 VINN.n95 4.5005
R71363 VINN.n261 VINN.n95 4.5005
R71364 VINN.n310 VINN.n95 4.5005
R71365 VINN.n260 VINN.n95 4.5005
R71366 VINN.n312 VINN.n95 4.5005
R71367 VINN.n259 VINN.n95 4.5005
R71368 VINN.n314 VINN.n95 4.5005
R71369 VINN.n258 VINN.n95 4.5005
R71370 VINN.n316 VINN.n95 4.5005
R71371 VINN.n257 VINN.n95 4.5005
R71372 VINN.n318 VINN.n95 4.5005
R71373 VINN.n256 VINN.n95 4.5005
R71374 VINN.n320 VINN.n95 4.5005
R71375 VINN.n255 VINN.n95 4.5005
R71376 VINN.n322 VINN.n95 4.5005
R71377 VINN.n254 VINN.n95 4.5005
R71378 VINN.n324 VINN.n95 4.5005
R71379 VINN.n253 VINN.n95 4.5005
R71380 VINN.n326 VINN.n95 4.5005
R71381 VINN.n252 VINN.n95 4.5005
R71382 VINN.n328 VINN.n95 4.5005
R71383 VINN.n251 VINN.n95 4.5005
R71384 VINN.n330 VINN.n95 4.5005
R71385 VINN.n250 VINN.n95 4.5005
R71386 VINN.n332 VINN.n95 4.5005
R71387 VINN.n249 VINN.n95 4.5005
R71388 VINN.n334 VINN.n95 4.5005
R71389 VINN.n248 VINN.n95 4.5005
R71390 VINN.n336 VINN.n95 4.5005
R71391 VINN.n247 VINN.n95 4.5005
R71392 VINN.n338 VINN.n95 4.5005
R71393 VINN.n246 VINN.n95 4.5005
R71394 VINN.n340 VINN.n95 4.5005
R71395 VINN.n245 VINN.n95 4.5005
R71396 VINN.n342 VINN.n95 4.5005
R71397 VINN.n244 VINN.n95 4.5005
R71398 VINN.n344 VINN.n95 4.5005
R71399 VINN.n243 VINN.n95 4.5005
R71400 VINN.n346 VINN.n95 4.5005
R71401 VINN.n242 VINN.n95 4.5005
R71402 VINN.n348 VINN.n95 4.5005
R71403 VINN.n241 VINN.n95 4.5005
R71404 VINN.n350 VINN.n95 4.5005
R71405 VINN.n240 VINN.n95 4.5005
R71406 VINN.n352 VINN.n95 4.5005
R71407 VINN.n239 VINN.n95 4.5005
R71408 VINN.n354 VINN.n95 4.5005
R71409 VINN.n238 VINN.n95 4.5005
R71410 VINN.n356 VINN.n95 4.5005
R71411 VINN.n237 VINN.n95 4.5005
R71412 VINN.n358 VINN.n95 4.5005
R71413 VINN.n236 VINN.n95 4.5005
R71414 VINN.n360 VINN.n95 4.5005
R71415 VINN.n235 VINN.n95 4.5005
R71416 VINN.n362 VINN.n95 4.5005
R71417 VINN.n234 VINN.n95 4.5005
R71418 VINN.n364 VINN.n95 4.5005
R71419 VINN.n233 VINN.n95 4.5005
R71420 VINN.n366 VINN.n95 4.5005
R71421 VINN.n232 VINN.n95 4.5005
R71422 VINN.n368 VINN.n95 4.5005
R71423 VINN.n231 VINN.n95 4.5005
R71424 VINN.n370 VINN.n95 4.5005
R71425 VINN.n230 VINN.n95 4.5005
R71426 VINN.n372 VINN.n95 4.5005
R71427 VINN.n229 VINN.n95 4.5005
R71428 VINN.n374 VINN.n95 4.5005
R71429 VINN.n228 VINN.n95 4.5005
R71430 VINN.n376 VINN.n95 4.5005
R71431 VINN.n227 VINN.n95 4.5005
R71432 VINN.n378 VINN.n95 4.5005
R71433 VINN.n226 VINN.n95 4.5005
R71434 VINN.n380 VINN.n95 4.5005
R71435 VINN.n225 VINN.n95 4.5005
R71436 VINN.n382 VINN.n95 4.5005
R71437 VINN.n224 VINN.n95 4.5005
R71438 VINN.n384 VINN.n95 4.5005
R71439 VINN.n223 VINN.n95 4.5005
R71440 VINN.n386 VINN.n95 4.5005
R71441 VINN.n222 VINN.n95 4.5005
R71442 VINN.n388 VINN.n95 4.5005
R71443 VINN.n221 VINN.n95 4.5005
R71444 VINN.n390 VINN.n95 4.5005
R71445 VINN.n220 VINN.n95 4.5005
R71446 VINN.n392 VINN.n95 4.5005
R71447 VINN.n219 VINN.n95 4.5005
R71448 VINN.n394 VINN.n95 4.5005
R71449 VINN.n218 VINN.n95 4.5005
R71450 VINN.n396 VINN.n95 4.5005
R71451 VINN.n217 VINN.n95 4.5005
R71452 VINN.n398 VINN.n95 4.5005
R71453 VINN.n216 VINN.n95 4.5005
R71454 VINN.n400 VINN.n95 4.5005
R71455 VINN.n215 VINN.n95 4.5005
R71456 VINN.n654 VINN.n95 4.5005
R71457 VINN.n656 VINN.n95 4.5005
R71458 VINN.n95 VINN.n0 4.5005
R71459 VINN.n278 VINN.n206 4.5005
R71460 VINN.n276 VINN.n206 4.5005
R71461 VINN.n280 VINN.n206 4.5005
R71462 VINN.n275 VINN.n206 4.5005
R71463 VINN.n282 VINN.n206 4.5005
R71464 VINN.n274 VINN.n206 4.5005
R71465 VINN.n284 VINN.n206 4.5005
R71466 VINN.n273 VINN.n206 4.5005
R71467 VINN.n286 VINN.n206 4.5005
R71468 VINN.n272 VINN.n206 4.5005
R71469 VINN.n288 VINN.n206 4.5005
R71470 VINN.n271 VINN.n206 4.5005
R71471 VINN.n290 VINN.n206 4.5005
R71472 VINN.n270 VINN.n206 4.5005
R71473 VINN.n292 VINN.n206 4.5005
R71474 VINN.n269 VINN.n206 4.5005
R71475 VINN.n294 VINN.n206 4.5005
R71476 VINN.n268 VINN.n206 4.5005
R71477 VINN.n296 VINN.n206 4.5005
R71478 VINN.n267 VINN.n206 4.5005
R71479 VINN.n298 VINN.n206 4.5005
R71480 VINN.n266 VINN.n206 4.5005
R71481 VINN.n300 VINN.n206 4.5005
R71482 VINN.n265 VINN.n206 4.5005
R71483 VINN.n302 VINN.n206 4.5005
R71484 VINN.n264 VINN.n206 4.5005
R71485 VINN.n304 VINN.n206 4.5005
R71486 VINN.n263 VINN.n206 4.5005
R71487 VINN.n306 VINN.n206 4.5005
R71488 VINN.n262 VINN.n206 4.5005
R71489 VINN.n308 VINN.n206 4.5005
R71490 VINN.n261 VINN.n206 4.5005
R71491 VINN.n310 VINN.n206 4.5005
R71492 VINN.n260 VINN.n206 4.5005
R71493 VINN.n312 VINN.n206 4.5005
R71494 VINN.n259 VINN.n206 4.5005
R71495 VINN.n314 VINN.n206 4.5005
R71496 VINN.n258 VINN.n206 4.5005
R71497 VINN.n316 VINN.n206 4.5005
R71498 VINN.n257 VINN.n206 4.5005
R71499 VINN.n318 VINN.n206 4.5005
R71500 VINN.n256 VINN.n206 4.5005
R71501 VINN.n320 VINN.n206 4.5005
R71502 VINN.n255 VINN.n206 4.5005
R71503 VINN.n322 VINN.n206 4.5005
R71504 VINN.n254 VINN.n206 4.5005
R71505 VINN.n324 VINN.n206 4.5005
R71506 VINN.n253 VINN.n206 4.5005
R71507 VINN.n326 VINN.n206 4.5005
R71508 VINN.n252 VINN.n206 4.5005
R71509 VINN.n328 VINN.n206 4.5005
R71510 VINN.n251 VINN.n206 4.5005
R71511 VINN.n330 VINN.n206 4.5005
R71512 VINN.n250 VINN.n206 4.5005
R71513 VINN.n332 VINN.n206 4.5005
R71514 VINN.n249 VINN.n206 4.5005
R71515 VINN.n334 VINN.n206 4.5005
R71516 VINN.n248 VINN.n206 4.5005
R71517 VINN.n336 VINN.n206 4.5005
R71518 VINN.n247 VINN.n206 4.5005
R71519 VINN.n338 VINN.n206 4.5005
R71520 VINN.n246 VINN.n206 4.5005
R71521 VINN.n340 VINN.n206 4.5005
R71522 VINN.n245 VINN.n206 4.5005
R71523 VINN.n342 VINN.n206 4.5005
R71524 VINN.n244 VINN.n206 4.5005
R71525 VINN.n344 VINN.n206 4.5005
R71526 VINN.n243 VINN.n206 4.5005
R71527 VINN.n346 VINN.n206 4.5005
R71528 VINN.n242 VINN.n206 4.5005
R71529 VINN.n348 VINN.n206 4.5005
R71530 VINN.n241 VINN.n206 4.5005
R71531 VINN.n350 VINN.n206 4.5005
R71532 VINN.n240 VINN.n206 4.5005
R71533 VINN.n352 VINN.n206 4.5005
R71534 VINN.n239 VINN.n206 4.5005
R71535 VINN.n354 VINN.n206 4.5005
R71536 VINN.n238 VINN.n206 4.5005
R71537 VINN.n356 VINN.n206 4.5005
R71538 VINN.n237 VINN.n206 4.5005
R71539 VINN.n358 VINN.n206 4.5005
R71540 VINN.n236 VINN.n206 4.5005
R71541 VINN.n360 VINN.n206 4.5005
R71542 VINN.n235 VINN.n206 4.5005
R71543 VINN.n362 VINN.n206 4.5005
R71544 VINN.n234 VINN.n206 4.5005
R71545 VINN.n364 VINN.n206 4.5005
R71546 VINN.n233 VINN.n206 4.5005
R71547 VINN.n366 VINN.n206 4.5005
R71548 VINN.n232 VINN.n206 4.5005
R71549 VINN.n368 VINN.n206 4.5005
R71550 VINN.n231 VINN.n206 4.5005
R71551 VINN.n370 VINN.n206 4.5005
R71552 VINN.n230 VINN.n206 4.5005
R71553 VINN.n372 VINN.n206 4.5005
R71554 VINN.n229 VINN.n206 4.5005
R71555 VINN.n374 VINN.n206 4.5005
R71556 VINN.n228 VINN.n206 4.5005
R71557 VINN.n376 VINN.n206 4.5005
R71558 VINN.n227 VINN.n206 4.5005
R71559 VINN.n378 VINN.n206 4.5005
R71560 VINN.n226 VINN.n206 4.5005
R71561 VINN.n380 VINN.n206 4.5005
R71562 VINN.n225 VINN.n206 4.5005
R71563 VINN.n382 VINN.n206 4.5005
R71564 VINN.n224 VINN.n206 4.5005
R71565 VINN.n384 VINN.n206 4.5005
R71566 VINN.n223 VINN.n206 4.5005
R71567 VINN.n386 VINN.n206 4.5005
R71568 VINN.n222 VINN.n206 4.5005
R71569 VINN.n388 VINN.n206 4.5005
R71570 VINN.n221 VINN.n206 4.5005
R71571 VINN.n390 VINN.n206 4.5005
R71572 VINN.n220 VINN.n206 4.5005
R71573 VINN.n392 VINN.n206 4.5005
R71574 VINN.n219 VINN.n206 4.5005
R71575 VINN.n394 VINN.n206 4.5005
R71576 VINN.n218 VINN.n206 4.5005
R71577 VINN.n396 VINN.n206 4.5005
R71578 VINN.n217 VINN.n206 4.5005
R71579 VINN.n398 VINN.n206 4.5005
R71580 VINN.n216 VINN.n206 4.5005
R71581 VINN.n400 VINN.n206 4.5005
R71582 VINN.n215 VINN.n206 4.5005
R71583 VINN.n654 VINN.n206 4.5005
R71584 VINN.n656 VINN.n206 4.5005
R71585 VINN.n206 VINN.n0 4.5005
R71586 VINN.n278 VINN.n94 4.5005
R71587 VINN.n276 VINN.n94 4.5005
R71588 VINN.n280 VINN.n94 4.5005
R71589 VINN.n275 VINN.n94 4.5005
R71590 VINN.n282 VINN.n94 4.5005
R71591 VINN.n274 VINN.n94 4.5005
R71592 VINN.n284 VINN.n94 4.5005
R71593 VINN.n273 VINN.n94 4.5005
R71594 VINN.n286 VINN.n94 4.5005
R71595 VINN.n272 VINN.n94 4.5005
R71596 VINN.n288 VINN.n94 4.5005
R71597 VINN.n271 VINN.n94 4.5005
R71598 VINN.n290 VINN.n94 4.5005
R71599 VINN.n270 VINN.n94 4.5005
R71600 VINN.n292 VINN.n94 4.5005
R71601 VINN.n269 VINN.n94 4.5005
R71602 VINN.n294 VINN.n94 4.5005
R71603 VINN.n268 VINN.n94 4.5005
R71604 VINN.n296 VINN.n94 4.5005
R71605 VINN.n267 VINN.n94 4.5005
R71606 VINN.n298 VINN.n94 4.5005
R71607 VINN.n266 VINN.n94 4.5005
R71608 VINN.n300 VINN.n94 4.5005
R71609 VINN.n265 VINN.n94 4.5005
R71610 VINN.n302 VINN.n94 4.5005
R71611 VINN.n264 VINN.n94 4.5005
R71612 VINN.n304 VINN.n94 4.5005
R71613 VINN.n263 VINN.n94 4.5005
R71614 VINN.n306 VINN.n94 4.5005
R71615 VINN.n262 VINN.n94 4.5005
R71616 VINN.n308 VINN.n94 4.5005
R71617 VINN.n261 VINN.n94 4.5005
R71618 VINN.n310 VINN.n94 4.5005
R71619 VINN.n260 VINN.n94 4.5005
R71620 VINN.n312 VINN.n94 4.5005
R71621 VINN.n259 VINN.n94 4.5005
R71622 VINN.n314 VINN.n94 4.5005
R71623 VINN.n258 VINN.n94 4.5005
R71624 VINN.n316 VINN.n94 4.5005
R71625 VINN.n257 VINN.n94 4.5005
R71626 VINN.n318 VINN.n94 4.5005
R71627 VINN.n256 VINN.n94 4.5005
R71628 VINN.n320 VINN.n94 4.5005
R71629 VINN.n255 VINN.n94 4.5005
R71630 VINN.n322 VINN.n94 4.5005
R71631 VINN.n254 VINN.n94 4.5005
R71632 VINN.n324 VINN.n94 4.5005
R71633 VINN.n253 VINN.n94 4.5005
R71634 VINN.n326 VINN.n94 4.5005
R71635 VINN.n252 VINN.n94 4.5005
R71636 VINN.n328 VINN.n94 4.5005
R71637 VINN.n251 VINN.n94 4.5005
R71638 VINN.n330 VINN.n94 4.5005
R71639 VINN.n250 VINN.n94 4.5005
R71640 VINN.n332 VINN.n94 4.5005
R71641 VINN.n249 VINN.n94 4.5005
R71642 VINN.n334 VINN.n94 4.5005
R71643 VINN.n248 VINN.n94 4.5005
R71644 VINN.n336 VINN.n94 4.5005
R71645 VINN.n247 VINN.n94 4.5005
R71646 VINN.n338 VINN.n94 4.5005
R71647 VINN.n246 VINN.n94 4.5005
R71648 VINN.n340 VINN.n94 4.5005
R71649 VINN.n245 VINN.n94 4.5005
R71650 VINN.n342 VINN.n94 4.5005
R71651 VINN.n244 VINN.n94 4.5005
R71652 VINN.n344 VINN.n94 4.5005
R71653 VINN.n243 VINN.n94 4.5005
R71654 VINN.n346 VINN.n94 4.5005
R71655 VINN.n242 VINN.n94 4.5005
R71656 VINN.n348 VINN.n94 4.5005
R71657 VINN.n241 VINN.n94 4.5005
R71658 VINN.n350 VINN.n94 4.5005
R71659 VINN.n240 VINN.n94 4.5005
R71660 VINN.n352 VINN.n94 4.5005
R71661 VINN.n239 VINN.n94 4.5005
R71662 VINN.n354 VINN.n94 4.5005
R71663 VINN.n238 VINN.n94 4.5005
R71664 VINN.n356 VINN.n94 4.5005
R71665 VINN.n237 VINN.n94 4.5005
R71666 VINN.n358 VINN.n94 4.5005
R71667 VINN.n236 VINN.n94 4.5005
R71668 VINN.n360 VINN.n94 4.5005
R71669 VINN.n235 VINN.n94 4.5005
R71670 VINN.n362 VINN.n94 4.5005
R71671 VINN.n234 VINN.n94 4.5005
R71672 VINN.n364 VINN.n94 4.5005
R71673 VINN.n233 VINN.n94 4.5005
R71674 VINN.n366 VINN.n94 4.5005
R71675 VINN.n232 VINN.n94 4.5005
R71676 VINN.n368 VINN.n94 4.5005
R71677 VINN.n231 VINN.n94 4.5005
R71678 VINN.n370 VINN.n94 4.5005
R71679 VINN.n230 VINN.n94 4.5005
R71680 VINN.n372 VINN.n94 4.5005
R71681 VINN.n229 VINN.n94 4.5005
R71682 VINN.n374 VINN.n94 4.5005
R71683 VINN.n228 VINN.n94 4.5005
R71684 VINN.n376 VINN.n94 4.5005
R71685 VINN.n227 VINN.n94 4.5005
R71686 VINN.n378 VINN.n94 4.5005
R71687 VINN.n226 VINN.n94 4.5005
R71688 VINN.n380 VINN.n94 4.5005
R71689 VINN.n225 VINN.n94 4.5005
R71690 VINN.n382 VINN.n94 4.5005
R71691 VINN.n224 VINN.n94 4.5005
R71692 VINN.n384 VINN.n94 4.5005
R71693 VINN.n223 VINN.n94 4.5005
R71694 VINN.n386 VINN.n94 4.5005
R71695 VINN.n222 VINN.n94 4.5005
R71696 VINN.n388 VINN.n94 4.5005
R71697 VINN.n221 VINN.n94 4.5005
R71698 VINN.n390 VINN.n94 4.5005
R71699 VINN.n220 VINN.n94 4.5005
R71700 VINN.n392 VINN.n94 4.5005
R71701 VINN.n219 VINN.n94 4.5005
R71702 VINN.n394 VINN.n94 4.5005
R71703 VINN.n218 VINN.n94 4.5005
R71704 VINN.n396 VINN.n94 4.5005
R71705 VINN.n217 VINN.n94 4.5005
R71706 VINN.n398 VINN.n94 4.5005
R71707 VINN.n216 VINN.n94 4.5005
R71708 VINN.n400 VINN.n94 4.5005
R71709 VINN.n215 VINN.n94 4.5005
R71710 VINN.n654 VINN.n94 4.5005
R71711 VINN.n656 VINN.n94 4.5005
R71712 VINN.n94 VINN.n0 4.5005
R71713 VINN.n278 VINN.n207 4.5005
R71714 VINN.n276 VINN.n207 4.5005
R71715 VINN.n280 VINN.n207 4.5005
R71716 VINN.n275 VINN.n207 4.5005
R71717 VINN.n282 VINN.n207 4.5005
R71718 VINN.n274 VINN.n207 4.5005
R71719 VINN.n284 VINN.n207 4.5005
R71720 VINN.n273 VINN.n207 4.5005
R71721 VINN.n286 VINN.n207 4.5005
R71722 VINN.n272 VINN.n207 4.5005
R71723 VINN.n288 VINN.n207 4.5005
R71724 VINN.n271 VINN.n207 4.5005
R71725 VINN.n290 VINN.n207 4.5005
R71726 VINN.n270 VINN.n207 4.5005
R71727 VINN.n292 VINN.n207 4.5005
R71728 VINN.n269 VINN.n207 4.5005
R71729 VINN.n294 VINN.n207 4.5005
R71730 VINN.n268 VINN.n207 4.5005
R71731 VINN.n296 VINN.n207 4.5005
R71732 VINN.n267 VINN.n207 4.5005
R71733 VINN.n298 VINN.n207 4.5005
R71734 VINN.n266 VINN.n207 4.5005
R71735 VINN.n300 VINN.n207 4.5005
R71736 VINN.n265 VINN.n207 4.5005
R71737 VINN.n302 VINN.n207 4.5005
R71738 VINN.n264 VINN.n207 4.5005
R71739 VINN.n304 VINN.n207 4.5005
R71740 VINN.n263 VINN.n207 4.5005
R71741 VINN.n306 VINN.n207 4.5005
R71742 VINN.n262 VINN.n207 4.5005
R71743 VINN.n308 VINN.n207 4.5005
R71744 VINN.n261 VINN.n207 4.5005
R71745 VINN.n310 VINN.n207 4.5005
R71746 VINN.n260 VINN.n207 4.5005
R71747 VINN.n312 VINN.n207 4.5005
R71748 VINN.n259 VINN.n207 4.5005
R71749 VINN.n314 VINN.n207 4.5005
R71750 VINN.n258 VINN.n207 4.5005
R71751 VINN.n316 VINN.n207 4.5005
R71752 VINN.n257 VINN.n207 4.5005
R71753 VINN.n318 VINN.n207 4.5005
R71754 VINN.n256 VINN.n207 4.5005
R71755 VINN.n320 VINN.n207 4.5005
R71756 VINN.n255 VINN.n207 4.5005
R71757 VINN.n322 VINN.n207 4.5005
R71758 VINN.n254 VINN.n207 4.5005
R71759 VINN.n324 VINN.n207 4.5005
R71760 VINN.n253 VINN.n207 4.5005
R71761 VINN.n326 VINN.n207 4.5005
R71762 VINN.n252 VINN.n207 4.5005
R71763 VINN.n328 VINN.n207 4.5005
R71764 VINN.n251 VINN.n207 4.5005
R71765 VINN.n330 VINN.n207 4.5005
R71766 VINN.n250 VINN.n207 4.5005
R71767 VINN.n332 VINN.n207 4.5005
R71768 VINN.n249 VINN.n207 4.5005
R71769 VINN.n334 VINN.n207 4.5005
R71770 VINN.n248 VINN.n207 4.5005
R71771 VINN.n336 VINN.n207 4.5005
R71772 VINN.n247 VINN.n207 4.5005
R71773 VINN.n338 VINN.n207 4.5005
R71774 VINN.n246 VINN.n207 4.5005
R71775 VINN.n340 VINN.n207 4.5005
R71776 VINN.n245 VINN.n207 4.5005
R71777 VINN.n342 VINN.n207 4.5005
R71778 VINN.n244 VINN.n207 4.5005
R71779 VINN.n344 VINN.n207 4.5005
R71780 VINN.n243 VINN.n207 4.5005
R71781 VINN.n346 VINN.n207 4.5005
R71782 VINN.n242 VINN.n207 4.5005
R71783 VINN.n348 VINN.n207 4.5005
R71784 VINN.n241 VINN.n207 4.5005
R71785 VINN.n350 VINN.n207 4.5005
R71786 VINN.n240 VINN.n207 4.5005
R71787 VINN.n352 VINN.n207 4.5005
R71788 VINN.n239 VINN.n207 4.5005
R71789 VINN.n354 VINN.n207 4.5005
R71790 VINN.n238 VINN.n207 4.5005
R71791 VINN.n356 VINN.n207 4.5005
R71792 VINN.n237 VINN.n207 4.5005
R71793 VINN.n358 VINN.n207 4.5005
R71794 VINN.n236 VINN.n207 4.5005
R71795 VINN.n360 VINN.n207 4.5005
R71796 VINN.n235 VINN.n207 4.5005
R71797 VINN.n362 VINN.n207 4.5005
R71798 VINN.n234 VINN.n207 4.5005
R71799 VINN.n364 VINN.n207 4.5005
R71800 VINN.n233 VINN.n207 4.5005
R71801 VINN.n366 VINN.n207 4.5005
R71802 VINN.n232 VINN.n207 4.5005
R71803 VINN.n368 VINN.n207 4.5005
R71804 VINN.n231 VINN.n207 4.5005
R71805 VINN.n370 VINN.n207 4.5005
R71806 VINN.n230 VINN.n207 4.5005
R71807 VINN.n372 VINN.n207 4.5005
R71808 VINN.n229 VINN.n207 4.5005
R71809 VINN.n374 VINN.n207 4.5005
R71810 VINN.n228 VINN.n207 4.5005
R71811 VINN.n376 VINN.n207 4.5005
R71812 VINN.n227 VINN.n207 4.5005
R71813 VINN.n378 VINN.n207 4.5005
R71814 VINN.n226 VINN.n207 4.5005
R71815 VINN.n380 VINN.n207 4.5005
R71816 VINN.n225 VINN.n207 4.5005
R71817 VINN.n382 VINN.n207 4.5005
R71818 VINN.n224 VINN.n207 4.5005
R71819 VINN.n384 VINN.n207 4.5005
R71820 VINN.n223 VINN.n207 4.5005
R71821 VINN.n386 VINN.n207 4.5005
R71822 VINN.n222 VINN.n207 4.5005
R71823 VINN.n388 VINN.n207 4.5005
R71824 VINN.n221 VINN.n207 4.5005
R71825 VINN.n390 VINN.n207 4.5005
R71826 VINN.n220 VINN.n207 4.5005
R71827 VINN.n392 VINN.n207 4.5005
R71828 VINN.n219 VINN.n207 4.5005
R71829 VINN.n394 VINN.n207 4.5005
R71830 VINN.n218 VINN.n207 4.5005
R71831 VINN.n396 VINN.n207 4.5005
R71832 VINN.n217 VINN.n207 4.5005
R71833 VINN.n398 VINN.n207 4.5005
R71834 VINN.n216 VINN.n207 4.5005
R71835 VINN.n400 VINN.n207 4.5005
R71836 VINN.n215 VINN.n207 4.5005
R71837 VINN.n654 VINN.n207 4.5005
R71838 VINN.n656 VINN.n207 4.5005
R71839 VINN.n207 VINN.n0 4.5005
R71840 VINN.n278 VINN.n93 4.5005
R71841 VINN.n276 VINN.n93 4.5005
R71842 VINN.n280 VINN.n93 4.5005
R71843 VINN.n275 VINN.n93 4.5005
R71844 VINN.n282 VINN.n93 4.5005
R71845 VINN.n274 VINN.n93 4.5005
R71846 VINN.n284 VINN.n93 4.5005
R71847 VINN.n273 VINN.n93 4.5005
R71848 VINN.n286 VINN.n93 4.5005
R71849 VINN.n272 VINN.n93 4.5005
R71850 VINN.n288 VINN.n93 4.5005
R71851 VINN.n271 VINN.n93 4.5005
R71852 VINN.n290 VINN.n93 4.5005
R71853 VINN.n270 VINN.n93 4.5005
R71854 VINN.n292 VINN.n93 4.5005
R71855 VINN.n269 VINN.n93 4.5005
R71856 VINN.n294 VINN.n93 4.5005
R71857 VINN.n268 VINN.n93 4.5005
R71858 VINN.n296 VINN.n93 4.5005
R71859 VINN.n267 VINN.n93 4.5005
R71860 VINN.n298 VINN.n93 4.5005
R71861 VINN.n266 VINN.n93 4.5005
R71862 VINN.n300 VINN.n93 4.5005
R71863 VINN.n265 VINN.n93 4.5005
R71864 VINN.n302 VINN.n93 4.5005
R71865 VINN.n264 VINN.n93 4.5005
R71866 VINN.n304 VINN.n93 4.5005
R71867 VINN.n263 VINN.n93 4.5005
R71868 VINN.n306 VINN.n93 4.5005
R71869 VINN.n262 VINN.n93 4.5005
R71870 VINN.n308 VINN.n93 4.5005
R71871 VINN.n261 VINN.n93 4.5005
R71872 VINN.n310 VINN.n93 4.5005
R71873 VINN.n260 VINN.n93 4.5005
R71874 VINN.n312 VINN.n93 4.5005
R71875 VINN.n259 VINN.n93 4.5005
R71876 VINN.n314 VINN.n93 4.5005
R71877 VINN.n258 VINN.n93 4.5005
R71878 VINN.n316 VINN.n93 4.5005
R71879 VINN.n257 VINN.n93 4.5005
R71880 VINN.n318 VINN.n93 4.5005
R71881 VINN.n256 VINN.n93 4.5005
R71882 VINN.n320 VINN.n93 4.5005
R71883 VINN.n255 VINN.n93 4.5005
R71884 VINN.n322 VINN.n93 4.5005
R71885 VINN.n254 VINN.n93 4.5005
R71886 VINN.n324 VINN.n93 4.5005
R71887 VINN.n253 VINN.n93 4.5005
R71888 VINN.n326 VINN.n93 4.5005
R71889 VINN.n252 VINN.n93 4.5005
R71890 VINN.n328 VINN.n93 4.5005
R71891 VINN.n251 VINN.n93 4.5005
R71892 VINN.n330 VINN.n93 4.5005
R71893 VINN.n250 VINN.n93 4.5005
R71894 VINN.n332 VINN.n93 4.5005
R71895 VINN.n249 VINN.n93 4.5005
R71896 VINN.n334 VINN.n93 4.5005
R71897 VINN.n248 VINN.n93 4.5005
R71898 VINN.n336 VINN.n93 4.5005
R71899 VINN.n247 VINN.n93 4.5005
R71900 VINN.n338 VINN.n93 4.5005
R71901 VINN.n246 VINN.n93 4.5005
R71902 VINN.n340 VINN.n93 4.5005
R71903 VINN.n245 VINN.n93 4.5005
R71904 VINN.n342 VINN.n93 4.5005
R71905 VINN.n244 VINN.n93 4.5005
R71906 VINN.n344 VINN.n93 4.5005
R71907 VINN.n243 VINN.n93 4.5005
R71908 VINN.n346 VINN.n93 4.5005
R71909 VINN.n242 VINN.n93 4.5005
R71910 VINN.n348 VINN.n93 4.5005
R71911 VINN.n241 VINN.n93 4.5005
R71912 VINN.n350 VINN.n93 4.5005
R71913 VINN.n240 VINN.n93 4.5005
R71914 VINN.n352 VINN.n93 4.5005
R71915 VINN.n239 VINN.n93 4.5005
R71916 VINN.n354 VINN.n93 4.5005
R71917 VINN.n238 VINN.n93 4.5005
R71918 VINN.n356 VINN.n93 4.5005
R71919 VINN.n237 VINN.n93 4.5005
R71920 VINN.n358 VINN.n93 4.5005
R71921 VINN.n236 VINN.n93 4.5005
R71922 VINN.n360 VINN.n93 4.5005
R71923 VINN.n235 VINN.n93 4.5005
R71924 VINN.n362 VINN.n93 4.5005
R71925 VINN.n234 VINN.n93 4.5005
R71926 VINN.n364 VINN.n93 4.5005
R71927 VINN.n233 VINN.n93 4.5005
R71928 VINN.n366 VINN.n93 4.5005
R71929 VINN.n232 VINN.n93 4.5005
R71930 VINN.n368 VINN.n93 4.5005
R71931 VINN.n231 VINN.n93 4.5005
R71932 VINN.n370 VINN.n93 4.5005
R71933 VINN.n230 VINN.n93 4.5005
R71934 VINN.n372 VINN.n93 4.5005
R71935 VINN.n229 VINN.n93 4.5005
R71936 VINN.n374 VINN.n93 4.5005
R71937 VINN.n228 VINN.n93 4.5005
R71938 VINN.n376 VINN.n93 4.5005
R71939 VINN.n227 VINN.n93 4.5005
R71940 VINN.n378 VINN.n93 4.5005
R71941 VINN.n226 VINN.n93 4.5005
R71942 VINN.n380 VINN.n93 4.5005
R71943 VINN.n225 VINN.n93 4.5005
R71944 VINN.n382 VINN.n93 4.5005
R71945 VINN.n224 VINN.n93 4.5005
R71946 VINN.n384 VINN.n93 4.5005
R71947 VINN.n223 VINN.n93 4.5005
R71948 VINN.n386 VINN.n93 4.5005
R71949 VINN.n222 VINN.n93 4.5005
R71950 VINN.n388 VINN.n93 4.5005
R71951 VINN.n221 VINN.n93 4.5005
R71952 VINN.n390 VINN.n93 4.5005
R71953 VINN.n220 VINN.n93 4.5005
R71954 VINN.n392 VINN.n93 4.5005
R71955 VINN.n219 VINN.n93 4.5005
R71956 VINN.n394 VINN.n93 4.5005
R71957 VINN.n218 VINN.n93 4.5005
R71958 VINN.n396 VINN.n93 4.5005
R71959 VINN.n217 VINN.n93 4.5005
R71960 VINN.n398 VINN.n93 4.5005
R71961 VINN.n216 VINN.n93 4.5005
R71962 VINN.n400 VINN.n93 4.5005
R71963 VINN.n215 VINN.n93 4.5005
R71964 VINN.n654 VINN.n93 4.5005
R71965 VINN.n656 VINN.n93 4.5005
R71966 VINN.n93 VINN.n0 4.5005
R71967 VINN.n278 VINN.n208 4.5005
R71968 VINN.n276 VINN.n208 4.5005
R71969 VINN.n280 VINN.n208 4.5005
R71970 VINN.n275 VINN.n208 4.5005
R71971 VINN.n282 VINN.n208 4.5005
R71972 VINN.n274 VINN.n208 4.5005
R71973 VINN.n284 VINN.n208 4.5005
R71974 VINN.n273 VINN.n208 4.5005
R71975 VINN.n286 VINN.n208 4.5005
R71976 VINN.n272 VINN.n208 4.5005
R71977 VINN.n288 VINN.n208 4.5005
R71978 VINN.n271 VINN.n208 4.5005
R71979 VINN.n290 VINN.n208 4.5005
R71980 VINN.n270 VINN.n208 4.5005
R71981 VINN.n292 VINN.n208 4.5005
R71982 VINN.n269 VINN.n208 4.5005
R71983 VINN.n294 VINN.n208 4.5005
R71984 VINN.n268 VINN.n208 4.5005
R71985 VINN.n296 VINN.n208 4.5005
R71986 VINN.n267 VINN.n208 4.5005
R71987 VINN.n298 VINN.n208 4.5005
R71988 VINN.n266 VINN.n208 4.5005
R71989 VINN.n300 VINN.n208 4.5005
R71990 VINN.n265 VINN.n208 4.5005
R71991 VINN.n302 VINN.n208 4.5005
R71992 VINN.n264 VINN.n208 4.5005
R71993 VINN.n304 VINN.n208 4.5005
R71994 VINN.n263 VINN.n208 4.5005
R71995 VINN.n306 VINN.n208 4.5005
R71996 VINN.n262 VINN.n208 4.5005
R71997 VINN.n308 VINN.n208 4.5005
R71998 VINN.n261 VINN.n208 4.5005
R71999 VINN.n310 VINN.n208 4.5005
R72000 VINN.n260 VINN.n208 4.5005
R72001 VINN.n312 VINN.n208 4.5005
R72002 VINN.n259 VINN.n208 4.5005
R72003 VINN.n314 VINN.n208 4.5005
R72004 VINN.n258 VINN.n208 4.5005
R72005 VINN.n316 VINN.n208 4.5005
R72006 VINN.n257 VINN.n208 4.5005
R72007 VINN.n318 VINN.n208 4.5005
R72008 VINN.n256 VINN.n208 4.5005
R72009 VINN.n320 VINN.n208 4.5005
R72010 VINN.n255 VINN.n208 4.5005
R72011 VINN.n322 VINN.n208 4.5005
R72012 VINN.n254 VINN.n208 4.5005
R72013 VINN.n324 VINN.n208 4.5005
R72014 VINN.n253 VINN.n208 4.5005
R72015 VINN.n326 VINN.n208 4.5005
R72016 VINN.n252 VINN.n208 4.5005
R72017 VINN.n328 VINN.n208 4.5005
R72018 VINN.n251 VINN.n208 4.5005
R72019 VINN.n330 VINN.n208 4.5005
R72020 VINN.n250 VINN.n208 4.5005
R72021 VINN.n332 VINN.n208 4.5005
R72022 VINN.n249 VINN.n208 4.5005
R72023 VINN.n334 VINN.n208 4.5005
R72024 VINN.n248 VINN.n208 4.5005
R72025 VINN.n336 VINN.n208 4.5005
R72026 VINN.n247 VINN.n208 4.5005
R72027 VINN.n338 VINN.n208 4.5005
R72028 VINN.n246 VINN.n208 4.5005
R72029 VINN.n340 VINN.n208 4.5005
R72030 VINN.n245 VINN.n208 4.5005
R72031 VINN.n342 VINN.n208 4.5005
R72032 VINN.n244 VINN.n208 4.5005
R72033 VINN.n344 VINN.n208 4.5005
R72034 VINN.n243 VINN.n208 4.5005
R72035 VINN.n346 VINN.n208 4.5005
R72036 VINN.n242 VINN.n208 4.5005
R72037 VINN.n348 VINN.n208 4.5005
R72038 VINN.n241 VINN.n208 4.5005
R72039 VINN.n350 VINN.n208 4.5005
R72040 VINN.n240 VINN.n208 4.5005
R72041 VINN.n352 VINN.n208 4.5005
R72042 VINN.n239 VINN.n208 4.5005
R72043 VINN.n354 VINN.n208 4.5005
R72044 VINN.n238 VINN.n208 4.5005
R72045 VINN.n356 VINN.n208 4.5005
R72046 VINN.n237 VINN.n208 4.5005
R72047 VINN.n358 VINN.n208 4.5005
R72048 VINN.n236 VINN.n208 4.5005
R72049 VINN.n360 VINN.n208 4.5005
R72050 VINN.n235 VINN.n208 4.5005
R72051 VINN.n362 VINN.n208 4.5005
R72052 VINN.n234 VINN.n208 4.5005
R72053 VINN.n364 VINN.n208 4.5005
R72054 VINN.n233 VINN.n208 4.5005
R72055 VINN.n366 VINN.n208 4.5005
R72056 VINN.n232 VINN.n208 4.5005
R72057 VINN.n368 VINN.n208 4.5005
R72058 VINN.n231 VINN.n208 4.5005
R72059 VINN.n370 VINN.n208 4.5005
R72060 VINN.n230 VINN.n208 4.5005
R72061 VINN.n372 VINN.n208 4.5005
R72062 VINN.n229 VINN.n208 4.5005
R72063 VINN.n374 VINN.n208 4.5005
R72064 VINN.n228 VINN.n208 4.5005
R72065 VINN.n376 VINN.n208 4.5005
R72066 VINN.n227 VINN.n208 4.5005
R72067 VINN.n378 VINN.n208 4.5005
R72068 VINN.n226 VINN.n208 4.5005
R72069 VINN.n380 VINN.n208 4.5005
R72070 VINN.n225 VINN.n208 4.5005
R72071 VINN.n382 VINN.n208 4.5005
R72072 VINN.n224 VINN.n208 4.5005
R72073 VINN.n384 VINN.n208 4.5005
R72074 VINN.n223 VINN.n208 4.5005
R72075 VINN.n386 VINN.n208 4.5005
R72076 VINN.n222 VINN.n208 4.5005
R72077 VINN.n388 VINN.n208 4.5005
R72078 VINN.n221 VINN.n208 4.5005
R72079 VINN.n390 VINN.n208 4.5005
R72080 VINN.n220 VINN.n208 4.5005
R72081 VINN.n392 VINN.n208 4.5005
R72082 VINN.n219 VINN.n208 4.5005
R72083 VINN.n394 VINN.n208 4.5005
R72084 VINN.n218 VINN.n208 4.5005
R72085 VINN.n396 VINN.n208 4.5005
R72086 VINN.n217 VINN.n208 4.5005
R72087 VINN.n398 VINN.n208 4.5005
R72088 VINN.n216 VINN.n208 4.5005
R72089 VINN.n400 VINN.n208 4.5005
R72090 VINN.n215 VINN.n208 4.5005
R72091 VINN.n654 VINN.n208 4.5005
R72092 VINN.n656 VINN.n208 4.5005
R72093 VINN.n208 VINN.n0 4.5005
R72094 VINN.n278 VINN.n92 4.5005
R72095 VINN.n276 VINN.n92 4.5005
R72096 VINN.n280 VINN.n92 4.5005
R72097 VINN.n275 VINN.n92 4.5005
R72098 VINN.n282 VINN.n92 4.5005
R72099 VINN.n274 VINN.n92 4.5005
R72100 VINN.n284 VINN.n92 4.5005
R72101 VINN.n273 VINN.n92 4.5005
R72102 VINN.n286 VINN.n92 4.5005
R72103 VINN.n272 VINN.n92 4.5005
R72104 VINN.n288 VINN.n92 4.5005
R72105 VINN.n271 VINN.n92 4.5005
R72106 VINN.n290 VINN.n92 4.5005
R72107 VINN.n270 VINN.n92 4.5005
R72108 VINN.n292 VINN.n92 4.5005
R72109 VINN.n269 VINN.n92 4.5005
R72110 VINN.n294 VINN.n92 4.5005
R72111 VINN.n268 VINN.n92 4.5005
R72112 VINN.n296 VINN.n92 4.5005
R72113 VINN.n267 VINN.n92 4.5005
R72114 VINN.n298 VINN.n92 4.5005
R72115 VINN.n266 VINN.n92 4.5005
R72116 VINN.n300 VINN.n92 4.5005
R72117 VINN.n265 VINN.n92 4.5005
R72118 VINN.n302 VINN.n92 4.5005
R72119 VINN.n264 VINN.n92 4.5005
R72120 VINN.n304 VINN.n92 4.5005
R72121 VINN.n263 VINN.n92 4.5005
R72122 VINN.n306 VINN.n92 4.5005
R72123 VINN.n262 VINN.n92 4.5005
R72124 VINN.n308 VINN.n92 4.5005
R72125 VINN.n261 VINN.n92 4.5005
R72126 VINN.n310 VINN.n92 4.5005
R72127 VINN.n260 VINN.n92 4.5005
R72128 VINN.n312 VINN.n92 4.5005
R72129 VINN.n259 VINN.n92 4.5005
R72130 VINN.n314 VINN.n92 4.5005
R72131 VINN.n258 VINN.n92 4.5005
R72132 VINN.n316 VINN.n92 4.5005
R72133 VINN.n257 VINN.n92 4.5005
R72134 VINN.n318 VINN.n92 4.5005
R72135 VINN.n256 VINN.n92 4.5005
R72136 VINN.n320 VINN.n92 4.5005
R72137 VINN.n255 VINN.n92 4.5005
R72138 VINN.n322 VINN.n92 4.5005
R72139 VINN.n254 VINN.n92 4.5005
R72140 VINN.n324 VINN.n92 4.5005
R72141 VINN.n253 VINN.n92 4.5005
R72142 VINN.n326 VINN.n92 4.5005
R72143 VINN.n252 VINN.n92 4.5005
R72144 VINN.n328 VINN.n92 4.5005
R72145 VINN.n251 VINN.n92 4.5005
R72146 VINN.n330 VINN.n92 4.5005
R72147 VINN.n250 VINN.n92 4.5005
R72148 VINN.n332 VINN.n92 4.5005
R72149 VINN.n249 VINN.n92 4.5005
R72150 VINN.n334 VINN.n92 4.5005
R72151 VINN.n248 VINN.n92 4.5005
R72152 VINN.n336 VINN.n92 4.5005
R72153 VINN.n247 VINN.n92 4.5005
R72154 VINN.n338 VINN.n92 4.5005
R72155 VINN.n246 VINN.n92 4.5005
R72156 VINN.n340 VINN.n92 4.5005
R72157 VINN.n245 VINN.n92 4.5005
R72158 VINN.n342 VINN.n92 4.5005
R72159 VINN.n244 VINN.n92 4.5005
R72160 VINN.n344 VINN.n92 4.5005
R72161 VINN.n243 VINN.n92 4.5005
R72162 VINN.n346 VINN.n92 4.5005
R72163 VINN.n242 VINN.n92 4.5005
R72164 VINN.n348 VINN.n92 4.5005
R72165 VINN.n241 VINN.n92 4.5005
R72166 VINN.n350 VINN.n92 4.5005
R72167 VINN.n240 VINN.n92 4.5005
R72168 VINN.n352 VINN.n92 4.5005
R72169 VINN.n239 VINN.n92 4.5005
R72170 VINN.n354 VINN.n92 4.5005
R72171 VINN.n238 VINN.n92 4.5005
R72172 VINN.n356 VINN.n92 4.5005
R72173 VINN.n237 VINN.n92 4.5005
R72174 VINN.n358 VINN.n92 4.5005
R72175 VINN.n236 VINN.n92 4.5005
R72176 VINN.n360 VINN.n92 4.5005
R72177 VINN.n235 VINN.n92 4.5005
R72178 VINN.n362 VINN.n92 4.5005
R72179 VINN.n234 VINN.n92 4.5005
R72180 VINN.n364 VINN.n92 4.5005
R72181 VINN.n233 VINN.n92 4.5005
R72182 VINN.n366 VINN.n92 4.5005
R72183 VINN.n232 VINN.n92 4.5005
R72184 VINN.n368 VINN.n92 4.5005
R72185 VINN.n231 VINN.n92 4.5005
R72186 VINN.n370 VINN.n92 4.5005
R72187 VINN.n230 VINN.n92 4.5005
R72188 VINN.n372 VINN.n92 4.5005
R72189 VINN.n229 VINN.n92 4.5005
R72190 VINN.n374 VINN.n92 4.5005
R72191 VINN.n228 VINN.n92 4.5005
R72192 VINN.n376 VINN.n92 4.5005
R72193 VINN.n227 VINN.n92 4.5005
R72194 VINN.n378 VINN.n92 4.5005
R72195 VINN.n226 VINN.n92 4.5005
R72196 VINN.n380 VINN.n92 4.5005
R72197 VINN.n225 VINN.n92 4.5005
R72198 VINN.n382 VINN.n92 4.5005
R72199 VINN.n224 VINN.n92 4.5005
R72200 VINN.n384 VINN.n92 4.5005
R72201 VINN.n223 VINN.n92 4.5005
R72202 VINN.n386 VINN.n92 4.5005
R72203 VINN.n222 VINN.n92 4.5005
R72204 VINN.n388 VINN.n92 4.5005
R72205 VINN.n221 VINN.n92 4.5005
R72206 VINN.n390 VINN.n92 4.5005
R72207 VINN.n220 VINN.n92 4.5005
R72208 VINN.n392 VINN.n92 4.5005
R72209 VINN.n219 VINN.n92 4.5005
R72210 VINN.n394 VINN.n92 4.5005
R72211 VINN.n218 VINN.n92 4.5005
R72212 VINN.n396 VINN.n92 4.5005
R72213 VINN.n217 VINN.n92 4.5005
R72214 VINN.n398 VINN.n92 4.5005
R72215 VINN.n216 VINN.n92 4.5005
R72216 VINN.n400 VINN.n92 4.5005
R72217 VINN.n215 VINN.n92 4.5005
R72218 VINN.n654 VINN.n92 4.5005
R72219 VINN.n656 VINN.n92 4.5005
R72220 VINN.n92 VINN.n0 4.5005
R72221 VINN.n278 VINN.n209 4.5005
R72222 VINN.n276 VINN.n209 4.5005
R72223 VINN.n280 VINN.n209 4.5005
R72224 VINN.n275 VINN.n209 4.5005
R72225 VINN.n282 VINN.n209 4.5005
R72226 VINN.n274 VINN.n209 4.5005
R72227 VINN.n284 VINN.n209 4.5005
R72228 VINN.n273 VINN.n209 4.5005
R72229 VINN.n286 VINN.n209 4.5005
R72230 VINN.n272 VINN.n209 4.5005
R72231 VINN.n288 VINN.n209 4.5005
R72232 VINN.n271 VINN.n209 4.5005
R72233 VINN.n290 VINN.n209 4.5005
R72234 VINN.n270 VINN.n209 4.5005
R72235 VINN.n292 VINN.n209 4.5005
R72236 VINN.n269 VINN.n209 4.5005
R72237 VINN.n294 VINN.n209 4.5005
R72238 VINN.n268 VINN.n209 4.5005
R72239 VINN.n296 VINN.n209 4.5005
R72240 VINN.n267 VINN.n209 4.5005
R72241 VINN.n298 VINN.n209 4.5005
R72242 VINN.n266 VINN.n209 4.5005
R72243 VINN.n300 VINN.n209 4.5005
R72244 VINN.n265 VINN.n209 4.5005
R72245 VINN.n302 VINN.n209 4.5005
R72246 VINN.n264 VINN.n209 4.5005
R72247 VINN.n304 VINN.n209 4.5005
R72248 VINN.n263 VINN.n209 4.5005
R72249 VINN.n306 VINN.n209 4.5005
R72250 VINN.n262 VINN.n209 4.5005
R72251 VINN.n308 VINN.n209 4.5005
R72252 VINN.n261 VINN.n209 4.5005
R72253 VINN.n310 VINN.n209 4.5005
R72254 VINN.n260 VINN.n209 4.5005
R72255 VINN.n312 VINN.n209 4.5005
R72256 VINN.n259 VINN.n209 4.5005
R72257 VINN.n314 VINN.n209 4.5005
R72258 VINN.n258 VINN.n209 4.5005
R72259 VINN.n316 VINN.n209 4.5005
R72260 VINN.n257 VINN.n209 4.5005
R72261 VINN.n318 VINN.n209 4.5005
R72262 VINN.n256 VINN.n209 4.5005
R72263 VINN.n320 VINN.n209 4.5005
R72264 VINN.n255 VINN.n209 4.5005
R72265 VINN.n322 VINN.n209 4.5005
R72266 VINN.n254 VINN.n209 4.5005
R72267 VINN.n324 VINN.n209 4.5005
R72268 VINN.n253 VINN.n209 4.5005
R72269 VINN.n326 VINN.n209 4.5005
R72270 VINN.n252 VINN.n209 4.5005
R72271 VINN.n328 VINN.n209 4.5005
R72272 VINN.n251 VINN.n209 4.5005
R72273 VINN.n330 VINN.n209 4.5005
R72274 VINN.n250 VINN.n209 4.5005
R72275 VINN.n332 VINN.n209 4.5005
R72276 VINN.n249 VINN.n209 4.5005
R72277 VINN.n334 VINN.n209 4.5005
R72278 VINN.n248 VINN.n209 4.5005
R72279 VINN.n336 VINN.n209 4.5005
R72280 VINN.n247 VINN.n209 4.5005
R72281 VINN.n338 VINN.n209 4.5005
R72282 VINN.n246 VINN.n209 4.5005
R72283 VINN.n340 VINN.n209 4.5005
R72284 VINN.n245 VINN.n209 4.5005
R72285 VINN.n342 VINN.n209 4.5005
R72286 VINN.n244 VINN.n209 4.5005
R72287 VINN.n344 VINN.n209 4.5005
R72288 VINN.n243 VINN.n209 4.5005
R72289 VINN.n346 VINN.n209 4.5005
R72290 VINN.n242 VINN.n209 4.5005
R72291 VINN.n348 VINN.n209 4.5005
R72292 VINN.n241 VINN.n209 4.5005
R72293 VINN.n350 VINN.n209 4.5005
R72294 VINN.n240 VINN.n209 4.5005
R72295 VINN.n352 VINN.n209 4.5005
R72296 VINN.n239 VINN.n209 4.5005
R72297 VINN.n354 VINN.n209 4.5005
R72298 VINN.n238 VINN.n209 4.5005
R72299 VINN.n356 VINN.n209 4.5005
R72300 VINN.n237 VINN.n209 4.5005
R72301 VINN.n358 VINN.n209 4.5005
R72302 VINN.n236 VINN.n209 4.5005
R72303 VINN.n360 VINN.n209 4.5005
R72304 VINN.n235 VINN.n209 4.5005
R72305 VINN.n362 VINN.n209 4.5005
R72306 VINN.n234 VINN.n209 4.5005
R72307 VINN.n364 VINN.n209 4.5005
R72308 VINN.n233 VINN.n209 4.5005
R72309 VINN.n366 VINN.n209 4.5005
R72310 VINN.n232 VINN.n209 4.5005
R72311 VINN.n368 VINN.n209 4.5005
R72312 VINN.n231 VINN.n209 4.5005
R72313 VINN.n370 VINN.n209 4.5005
R72314 VINN.n230 VINN.n209 4.5005
R72315 VINN.n372 VINN.n209 4.5005
R72316 VINN.n229 VINN.n209 4.5005
R72317 VINN.n374 VINN.n209 4.5005
R72318 VINN.n228 VINN.n209 4.5005
R72319 VINN.n376 VINN.n209 4.5005
R72320 VINN.n227 VINN.n209 4.5005
R72321 VINN.n378 VINN.n209 4.5005
R72322 VINN.n226 VINN.n209 4.5005
R72323 VINN.n380 VINN.n209 4.5005
R72324 VINN.n225 VINN.n209 4.5005
R72325 VINN.n382 VINN.n209 4.5005
R72326 VINN.n224 VINN.n209 4.5005
R72327 VINN.n384 VINN.n209 4.5005
R72328 VINN.n223 VINN.n209 4.5005
R72329 VINN.n386 VINN.n209 4.5005
R72330 VINN.n222 VINN.n209 4.5005
R72331 VINN.n388 VINN.n209 4.5005
R72332 VINN.n221 VINN.n209 4.5005
R72333 VINN.n390 VINN.n209 4.5005
R72334 VINN.n220 VINN.n209 4.5005
R72335 VINN.n392 VINN.n209 4.5005
R72336 VINN.n219 VINN.n209 4.5005
R72337 VINN.n394 VINN.n209 4.5005
R72338 VINN.n218 VINN.n209 4.5005
R72339 VINN.n396 VINN.n209 4.5005
R72340 VINN.n217 VINN.n209 4.5005
R72341 VINN.n398 VINN.n209 4.5005
R72342 VINN.n216 VINN.n209 4.5005
R72343 VINN.n400 VINN.n209 4.5005
R72344 VINN.n215 VINN.n209 4.5005
R72345 VINN.n654 VINN.n209 4.5005
R72346 VINN.n656 VINN.n209 4.5005
R72347 VINN.n209 VINN.n0 4.5005
R72348 VINN.n278 VINN.n91 4.5005
R72349 VINN.n276 VINN.n91 4.5005
R72350 VINN.n280 VINN.n91 4.5005
R72351 VINN.n275 VINN.n91 4.5005
R72352 VINN.n282 VINN.n91 4.5005
R72353 VINN.n274 VINN.n91 4.5005
R72354 VINN.n284 VINN.n91 4.5005
R72355 VINN.n273 VINN.n91 4.5005
R72356 VINN.n286 VINN.n91 4.5005
R72357 VINN.n272 VINN.n91 4.5005
R72358 VINN.n288 VINN.n91 4.5005
R72359 VINN.n271 VINN.n91 4.5005
R72360 VINN.n290 VINN.n91 4.5005
R72361 VINN.n270 VINN.n91 4.5005
R72362 VINN.n292 VINN.n91 4.5005
R72363 VINN.n269 VINN.n91 4.5005
R72364 VINN.n294 VINN.n91 4.5005
R72365 VINN.n268 VINN.n91 4.5005
R72366 VINN.n296 VINN.n91 4.5005
R72367 VINN.n267 VINN.n91 4.5005
R72368 VINN.n298 VINN.n91 4.5005
R72369 VINN.n266 VINN.n91 4.5005
R72370 VINN.n300 VINN.n91 4.5005
R72371 VINN.n265 VINN.n91 4.5005
R72372 VINN.n302 VINN.n91 4.5005
R72373 VINN.n264 VINN.n91 4.5005
R72374 VINN.n304 VINN.n91 4.5005
R72375 VINN.n263 VINN.n91 4.5005
R72376 VINN.n306 VINN.n91 4.5005
R72377 VINN.n262 VINN.n91 4.5005
R72378 VINN.n308 VINN.n91 4.5005
R72379 VINN.n261 VINN.n91 4.5005
R72380 VINN.n310 VINN.n91 4.5005
R72381 VINN.n260 VINN.n91 4.5005
R72382 VINN.n312 VINN.n91 4.5005
R72383 VINN.n259 VINN.n91 4.5005
R72384 VINN.n314 VINN.n91 4.5005
R72385 VINN.n258 VINN.n91 4.5005
R72386 VINN.n316 VINN.n91 4.5005
R72387 VINN.n257 VINN.n91 4.5005
R72388 VINN.n318 VINN.n91 4.5005
R72389 VINN.n256 VINN.n91 4.5005
R72390 VINN.n320 VINN.n91 4.5005
R72391 VINN.n255 VINN.n91 4.5005
R72392 VINN.n322 VINN.n91 4.5005
R72393 VINN.n254 VINN.n91 4.5005
R72394 VINN.n324 VINN.n91 4.5005
R72395 VINN.n253 VINN.n91 4.5005
R72396 VINN.n326 VINN.n91 4.5005
R72397 VINN.n252 VINN.n91 4.5005
R72398 VINN.n328 VINN.n91 4.5005
R72399 VINN.n251 VINN.n91 4.5005
R72400 VINN.n330 VINN.n91 4.5005
R72401 VINN.n250 VINN.n91 4.5005
R72402 VINN.n332 VINN.n91 4.5005
R72403 VINN.n249 VINN.n91 4.5005
R72404 VINN.n334 VINN.n91 4.5005
R72405 VINN.n248 VINN.n91 4.5005
R72406 VINN.n336 VINN.n91 4.5005
R72407 VINN.n247 VINN.n91 4.5005
R72408 VINN.n338 VINN.n91 4.5005
R72409 VINN.n246 VINN.n91 4.5005
R72410 VINN.n340 VINN.n91 4.5005
R72411 VINN.n245 VINN.n91 4.5005
R72412 VINN.n342 VINN.n91 4.5005
R72413 VINN.n244 VINN.n91 4.5005
R72414 VINN.n344 VINN.n91 4.5005
R72415 VINN.n243 VINN.n91 4.5005
R72416 VINN.n346 VINN.n91 4.5005
R72417 VINN.n242 VINN.n91 4.5005
R72418 VINN.n348 VINN.n91 4.5005
R72419 VINN.n241 VINN.n91 4.5005
R72420 VINN.n350 VINN.n91 4.5005
R72421 VINN.n240 VINN.n91 4.5005
R72422 VINN.n352 VINN.n91 4.5005
R72423 VINN.n239 VINN.n91 4.5005
R72424 VINN.n354 VINN.n91 4.5005
R72425 VINN.n238 VINN.n91 4.5005
R72426 VINN.n356 VINN.n91 4.5005
R72427 VINN.n237 VINN.n91 4.5005
R72428 VINN.n358 VINN.n91 4.5005
R72429 VINN.n236 VINN.n91 4.5005
R72430 VINN.n360 VINN.n91 4.5005
R72431 VINN.n235 VINN.n91 4.5005
R72432 VINN.n362 VINN.n91 4.5005
R72433 VINN.n234 VINN.n91 4.5005
R72434 VINN.n364 VINN.n91 4.5005
R72435 VINN.n233 VINN.n91 4.5005
R72436 VINN.n366 VINN.n91 4.5005
R72437 VINN.n232 VINN.n91 4.5005
R72438 VINN.n368 VINN.n91 4.5005
R72439 VINN.n231 VINN.n91 4.5005
R72440 VINN.n370 VINN.n91 4.5005
R72441 VINN.n230 VINN.n91 4.5005
R72442 VINN.n372 VINN.n91 4.5005
R72443 VINN.n229 VINN.n91 4.5005
R72444 VINN.n374 VINN.n91 4.5005
R72445 VINN.n228 VINN.n91 4.5005
R72446 VINN.n376 VINN.n91 4.5005
R72447 VINN.n227 VINN.n91 4.5005
R72448 VINN.n378 VINN.n91 4.5005
R72449 VINN.n226 VINN.n91 4.5005
R72450 VINN.n380 VINN.n91 4.5005
R72451 VINN.n225 VINN.n91 4.5005
R72452 VINN.n382 VINN.n91 4.5005
R72453 VINN.n224 VINN.n91 4.5005
R72454 VINN.n384 VINN.n91 4.5005
R72455 VINN.n223 VINN.n91 4.5005
R72456 VINN.n386 VINN.n91 4.5005
R72457 VINN.n222 VINN.n91 4.5005
R72458 VINN.n388 VINN.n91 4.5005
R72459 VINN.n221 VINN.n91 4.5005
R72460 VINN.n390 VINN.n91 4.5005
R72461 VINN.n220 VINN.n91 4.5005
R72462 VINN.n392 VINN.n91 4.5005
R72463 VINN.n219 VINN.n91 4.5005
R72464 VINN.n394 VINN.n91 4.5005
R72465 VINN.n218 VINN.n91 4.5005
R72466 VINN.n396 VINN.n91 4.5005
R72467 VINN.n217 VINN.n91 4.5005
R72468 VINN.n398 VINN.n91 4.5005
R72469 VINN.n216 VINN.n91 4.5005
R72470 VINN.n400 VINN.n91 4.5005
R72471 VINN.n215 VINN.n91 4.5005
R72472 VINN.n654 VINN.n91 4.5005
R72473 VINN.n656 VINN.n91 4.5005
R72474 VINN.n91 VINN.n0 4.5005
R72475 VINN.n278 VINN.n210 4.5005
R72476 VINN.n276 VINN.n210 4.5005
R72477 VINN.n280 VINN.n210 4.5005
R72478 VINN.n275 VINN.n210 4.5005
R72479 VINN.n282 VINN.n210 4.5005
R72480 VINN.n274 VINN.n210 4.5005
R72481 VINN.n284 VINN.n210 4.5005
R72482 VINN.n273 VINN.n210 4.5005
R72483 VINN.n286 VINN.n210 4.5005
R72484 VINN.n272 VINN.n210 4.5005
R72485 VINN.n288 VINN.n210 4.5005
R72486 VINN.n271 VINN.n210 4.5005
R72487 VINN.n290 VINN.n210 4.5005
R72488 VINN.n270 VINN.n210 4.5005
R72489 VINN.n292 VINN.n210 4.5005
R72490 VINN.n269 VINN.n210 4.5005
R72491 VINN.n294 VINN.n210 4.5005
R72492 VINN.n268 VINN.n210 4.5005
R72493 VINN.n296 VINN.n210 4.5005
R72494 VINN.n267 VINN.n210 4.5005
R72495 VINN.n298 VINN.n210 4.5005
R72496 VINN.n266 VINN.n210 4.5005
R72497 VINN.n300 VINN.n210 4.5005
R72498 VINN.n265 VINN.n210 4.5005
R72499 VINN.n302 VINN.n210 4.5005
R72500 VINN.n264 VINN.n210 4.5005
R72501 VINN.n304 VINN.n210 4.5005
R72502 VINN.n263 VINN.n210 4.5005
R72503 VINN.n306 VINN.n210 4.5005
R72504 VINN.n262 VINN.n210 4.5005
R72505 VINN.n308 VINN.n210 4.5005
R72506 VINN.n261 VINN.n210 4.5005
R72507 VINN.n310 VINN.n210 4.5005
R72508 VINN.n260 VINN.n210 4.5005
R72509 VINN.n312 VINN.n210 4.5005
R72510 VINN.n259 VINN.n210 4.5005
R72511 VINN.n314 VINN.n210 4.5005
R72512 VINN.n258 VINN.n210 4.5005
R72513 VINN.n316 VINN.n210 4.5005
R72514 VINN.n257 VINN.n210 4.5005
R72515 VINN.n318 VINN.n210 4.5005
R72516 VINN.n256 VINN.n210 4.5005
R72517 VINN.n320 VINN.n210 4.5005
R72518 VINN.n255 VINN.n210 4.5005
R72519 VINN.n322 VINN.n210 4.5005
R72520 VINN.n254 VINN.n210 4.5005
R72521 VINN.n324 VINN.n210 4.5005
R72522 VINN.n253 VINN.n210 4.5005
R72523 VINN.n326 VINN.n210 4.5005
R72524 VINN.n252 VINN.n210 4.5005
R72525 VINN.n328 VINN.n210 4.5005
R72526 VINN.n251 VINN.n210 4.5005
R72527 VINN.n330 VINN.n210 4.5005
R72528 VINN.n250 VINN.n210 4.5005
R72529 VINN.n332 VINN.n210 4.5005
R72530 VINN.n249 VINN.n210 4.5005
R72531 VINN.n334 VINN.n210 4.5005
R72532 VINN.n248 VINN.n210 4.5005
R72533 VINN.n336 VINN.n210 4.5005
R72534 VINN.n247 VINN.n210 4.5005
R72535 VINN.n338 VINN.n210 4.5005
R72536 VINN.n246 VINN.n210 4.5005
R72537 VINN.n340 VINN.n210 4.5005
R72538 VINN.n245 VINN.n210 4.5005
R72539 VINN.n342 VINN.n210 4.5005
R72540 VINN.n244 VINN.n210 4.5005
R72541 VINN.n344 VINN.n210 4.5005
R72542 VINN.n243 VINN.n210 4.5005
R72543 VINN.n346 VINN.n210 4.5005
R72544 VINN.n242 VINN.n210 4.5005
R72545 VINN.n348 VINN.n210 4.5005
R72546 VINN.n241 VINN.n210 4.5005
R72547 VINN.n350 VINN.n210 4.5005
R72548 VINN.n240 VINN.n210 4.5005
R72549 VINN.n352 VINN.n210 4.5005
R72550 VINN.n239 VINN.n210 4.5005
R72551 VINN.n354 VINN.n210 4.5005
R72552 VINN.n238 VINN.n210 4.5005
R72553 VINN.n356 VINN.n210 4.5005
R72554 VINN.n237 VINN.n210 4.5005
R72555 VINN.n358 VINN.n210 4.5005
R72556 VINN.n236 VINN.n210 4.5005
R72557 VINN.n360 VINN.n210 4.5005
R72558 VINN.n235 VINN.n210 4.5005
R72559 VINN.n362 VINN.n210 4.5005
R72560 VINN.n234 VINN.n210 4.5005
R72561 VINN.n364 VINN.n210 4.5005
R72562 VINN.n233 VINN.n210 4.5005
R72563 VINN.n366 VINN.n210 4.5005
R72564 VINN.n232 VINN.n210 4.5005
R72565 VINN.n368 VINN.n210 4.5005
R72566 VINN.n231 VINN.n210 4.5005
R72567 VINN.n370 VINN.n210 4.5005
R72568 VINN.n230 VINN.n210 4.5005
R72569 VINN.n372 VINN.n210 4.5005
R72570 VINN.n229 VINN.n210 4.5005
R72571 VINN.n374 VINN.n210 4.5005
R72572 VINN.n228 VINN.n210 4.5005
R72573 VINN.n376 VINN.n210 4.5005
R72574 VINN.n227 VINN.n210 4.5005
R72575 VINN.n378 VINN.n210 4.5005
R72576 VINN.n226 VINN.n210 4.5005
R72577 VINN.n380 VINN.n210 4.5005
R72578 VINN.n225 VINN.n210 4.5005
R72579 VINN.n382 VINN.n210 4.5005
R72580 VINN.n224 VINN.n210 4.5005
R72581 VINN.n384 VINN.n210 4.5005
R72582 VINN.n223 VINN.n210 4.5005
R72583 VINN.n386 VINN.n210 4.5005
R72584 VINN.n222 VINN.n210 4.5005
R72585 VINN.n388 VINN.n210 4.5005
R72586 VINN.n221 VINN.n210 4.5005
R72587 VINN.n390 VINN.n210 4.5005
R72588 VINN.n220 VINN.n210 4.5005
R72589 VINN.n392 VINN.n210 4.5005
R72590 VINN.n219 VINN.n210 4.5005
R72591 VINN.n394 VINN.n210 4.5005
R72592 VINN.n218 VINN.n210 4.5005
R72593 VINN.n396 VINN.n210 4.5005
R72594 VINN.n217 VINN.n210 4.5005
R72595 VINN.n398 VINN.n210 4.5005
R72596 VINN.n216 VINN.n210 4.5005
R72597 VINN.n400 VINN.n210 4.5005
R72598 VINN.n215 VINN.n210 4.5005
R72599 VINN.n654 VINN.n210 4.5005
R72600 VINN.n656 VINN.n210 4.5005
R72601 VINN.n210 VINN.n0 4.5005
R72602 VINN.n278 VINN.n90 4.5005
R72603 VINN.n276 VINN.n90 4.5005
R72604 VINN.n280 VINN.n90 4.5005
R72605 VINN.n275 VINN.n90 4.5005
R72606 VINN.n282 VINN.n90 4.5005
R72607 VINN.n274 VINN.n90 4.5005
R72608 VINN.n284 VINN.n90 4.5005
R72609 VINN.n273 VINN.n90 4.5005
R72610 VINN.n286 VINN.n90 4.5005
R72611 VINN.n272 VINN.n90 4.5005
R72612 VINN.n288 VINN.n90 4.5005
R72613 VINN.n271 VINN.n90 4.5005
R72614 VINN.n290 VINN.n90 4.5005
R72615 VINN.n270 VINN.n90 4.5005
R72616 VINN.n292 VINN.n90 4.5005
R72617 VINN.n269 VINN.n90 4.5005
R72618 VINN.n294 VINN.n90 4.5005
R72619 VINN.n268 VINN.n90 4.5005
R72620 VINN.n296 VINN.n90 4.5005
R72621 VINN.n267 VINN.n90 4.5005
R72622 VINN.n298 VINN.n90 4.5005
R72623 VINN.n266 VINN.n90 4.5005
R72624 VINN.n300 VINN.n90 4.5005
R72625 VINN.n265 VINN.n90 4.5005
R72626 VINN.n302 VINN.n90 4.5005
R72627 VINN.n264 VINN.n90 4.5005
R72628 VINN.n304 VINN.n90 4.5005
R72629 VINN.n263 VINN.n90 4.5005
R72630 VINN.n306 VINN.n90 4.5005
R72631 VINN.n262 VINN.n90 4.5005
R72632 VINN.n308 VINN.n90 4.5005
R72633 VINN.n261 VINN.n90 4.5005
R72634 VINN.n310 VINN.n90 4.5005
R72635 VINN.n260 VINN.n90 4.5005
R72636 VINN.n312 VINN.n90 4.5005
R72637 VINN.n259 VINN.n90 4.5005
R72638 VINN.n314 VINN.n90 4.5005
R72639 VINN.n258 VINN.n90 4.5005
R72640 VINN.n316 VINN.n90 4.5005
R72641 VINN.n257 VINN.n90 4.5005
R72642 VINN.n318 VINN.n90 4.5005
R72643 VINN.n256 VINN.n90 4.5005
R72644 VINN.n320 VINN.n90 4.5005
R72645 VINN.n255 VINN.n90 4.5005
R72646 VINN.n322 VINN.n90 4.5005
R72647 VINN.n254 VINN.n90 4.5005
R72648 VINN.n324 VINN.n90 4.5005
R72649 VINN.n253 VINN.n90 4.5005
R72650 VINN.n326 VINN.n90 4.5005
R72651 VINN.n252 VINN.n90 4.5005
R72652 VINN.n328 VINN.n90 4.5005
R72653 VINN.n251 VINN.n90 4.5005
R72654 VINN.n330 VINN.n90 4.5005
R72655 VINN.n250 VINN.n90 4.5005
R72656 VINN.n332 VINN.n90 4.5005
R72657 VINN.n249 VINN.n90 4.5005
R72658 VINN.n334 VINN.n90 4.5005
R72659 VINN.n248 VINN.n90 4.5005
R72660 VINN.n336 VINN.n90 4.5005
R72661 VINN.n247 VINN.n90 4.5005
R72662 VINN.n338 VINN.n90 4.5005
R72663 VINN.n246 VINN.n90 4.5005
R72664 VINN.n340 VINN.n90 4.5005
R72665 VINN.n245 VINN.n90 4.5005
R72666 VINN.n342 VINN.n90 4.5005
R72667 VINN.n244 VINN.n90 4.5005
R72668 VINN.n344 VINN.n90 4.5005
R72669 VINN.n243 VINN.n90 4.5005
R72670 VINN.n346 VINN.n90 4.5005
R72671 VINN.n242 VINN.n90 4.5005
R72672 VINN.n348 VINN.n90 4.5005
R72673 VINN.n241 VINN.n90 4.5005
R72674 VINN.n350 VINN.n90 4.5005
R72675 VINN.n240 VINN.n90 4.5005
R72676 VINN.n352 VINN.n90 4.5005
R72677 VINN.n239 VINN.n90 4.5005
R72678 VINN.n354 VINN.n90 4.5005
R72679 VINN.n238 VINN.n90 4.5005
R72680 VINN.n356 VINN.n90 4.5005
R72681 VINN.n237 VINN.n90 4.5005
R72682 VINN.n358 VINN.n90 4.5005
R72683 VINN.n236 VINN.n90 4.5005
R72684 VINN.n360 VINN.n90 4.5005
R72685 VINN.n235 VINN.n90 4.5005
R72686 VINN.n362 VINN.n90 4.5005
R72687 VINN.n234 VINN.n90 4.5005
R72688 VINN.n364 VINN.n90 4.5005
R72689 VINN.n233 VINN.n90 4.5005
R72690 VINN.n366 VINN.n90 4.5005
R72691 VINN.n232 VINN.n90 4.5005
R72692 VINN.n368 VINN.n90 4.5005
R72693 VINN.n231 VINN.n90 4.5005
R72694 VINN.n370 VINN.n90 4.5005
R72695 VINN.n230 VINN.n90 4.5005
R72696 VINN.n372 VINN.n90 4.5005
R72697 VINN.n229 VINN.n90 4.5005
R72698 VINN.n374 VINN.n90 4.5005
R72699 VINN.n228 VINN.n90 4.5005
R72700 VINN.n376 VINN.n90 4.5005
R72701 VINN.n227 VINN.n90 4.5005
R72702 VINN.n378 VINN.n90 4.5005
R72703 VINN.n226 VINN.n90 4.5005
R72704 VINN.n380 VINN.n90 4.5005
R72705 VINN.n225 VINN.n90 4.5005
R72706 VINN.n382 VINN.n90 4.5005
R72707 VINN.n224 VINN.n90 4.5005
R72708 VINN.n384 VINN.n90 4.5005
R72709 VINN.n223 VINN.n90 4.5005
R72710 VINN.n386 VINN.n90 4.5005
R72711 VINN.n222 VINN.n90 4.5005
R72712 VINN.n388 VINN.n90 4.5005
R72713 VINN.n221 VINN.n90 4.5005
R72714 VINN.n390 VINN.n90 4.5005
R72715 VINN.n220 VINN.n90 4.5005
R72716 VINN.n392 VINN.n90 4.5005
R72717 VINN.n219 VINN.n90 4.5005
R72718 VINN.n394 VINN.n90 4.5005
R72719 VINN.n218 VINN.n90 4.5005
R72720 VINN.n396 VINN.n90 4.5005
R72721 VINN.n217 VINN.n90 4.5005
R72722 VINN.n398 VINN.n90 4.5005
R72723 VINN.n216 VINN.n90 4.5005
R72724 VINN.n400 VINN.n90 4.5005
R72725 VINN.n215 VINN.n90 4.5005
R72726 VINN.n654 VINN.n90 4.5005
R72727 VINN.n656 VINN.n90 4.5005
R72728 VINN.n90 VINN.n0 4.5005
R72729 VINN.n278 VINN.n211 4.5005
R72730 VINN.n276 VINN.n211 4.5005
R72731 VINN.n280 VINN.n211 4.5005
R72732 VINN.n275 VINN.n211 4.5005
R72733 VINN.n282 VINN.n211 4.5005
R72734 VINN.n274 VINN.n211 4.5005
R72735 VINN.n284 VINN.n211 4.5005
R72736 VINN.n273 VINN.n211 4.5005
R72737 VINN.n286 VINN.n211 4.5005
R72738 VINN.n272 VINN.n211 4.5005
R72739 VINN.n288 VINN.n211 4.5005
R72740 VINN.n271 VINN.n211 4.5005
R72741 VINN.n290 VINN.n211 4.5005
R72742 VINN.n270 VINN.n211 4.5005
R72743 VINN.n292 VINN.n211 4.5005
R72744 VINN.n269 VINN.n211 4.5005
R72745 VINN.n294 VINN.n211 4.5005
R72746 VINN.n268 VINN.n211 4.5005
R72747 VINN.n296 VINN.n211 4.5005
R72748 VINN.n267 VINN.n211 4.5005
R72749 VINN.n298 VINN.n211 4.5005
R72750 VINN.n266 VINN.n211 4.5005
R72751 VINN.n300 VINN.n211 4.5005
R72752 VINN.n265 VINN.n211 4.5005
R72753 VINN.n302 VINN.n211 4.5005
R72754 VINN.n264 VINN.n211 4.5005
R72755 VINN.n304 VINN.n211 4.5005
R72756 VINN.n263 VINN.n211 4.5005
R72757 VINN.n306 VINN.n211 4.5005
R72758 VINN.n262 VINN.n211 4.5005
R72759 VINN.n308 VINN.n211 4.5005
R72760 VINN.n261 VINN.n211 4.5005
R72761 VINN.n310 VINN.n211 4.5005
R72762 VINN.n260 VINN.n211 4.5005
R72763 VINN.n312 VINN.n211 4.5005
R72764 VINN.n259 VINN.n211 4.5005
R72765 VINN.n314 VINN.n211 4.5005
R72766 VINN.n258 VINN.n211 4.5005
R72767 VINN.n316 VINN.n211 4.5005
R72768 VINN.n257 VINN.n211 4.5005
R72769 VINN.n318 VINN.n211 4.5005
R72770 VINN.n256 VINN.n211 4.5005
R72771 VINN.n320 VINN.n211 4.5005
R72772 VINN.n255 VINN.n211 4.5005
R72773 VINN.n322 VINN.n211 4.5005
R72774 VINN.n254 VINN.n211 4.5005
R72775 VINN.n324 VINN.n211 4.5005
R72776 VINN.n253 VINN.n211 4.5005
R72777 VINN.n326 VINN.n211 4.5005
R72778 VINN.n252 VINN.n211 4.5005
R72779 VINN.n328 VINN.n211 4.5005
R72780 VINN.n251 VINN.n211 4.5005
R72781 VINN.n330 VINN.n211 4.5005
R72782 VINN.n250 VINN.n211 4.5005
R72783 VINN.n332 VINN.n211 4.5005
R72784 VINN.n249 VINN.n211 4.5005
R72785 VINN.n334 VINN.n211 4.5005
R72786 VINN.n248 VINN.n211 4.5005
R72787 VINN.n336 VINN.n211 4.5005
R72788 VINN.n247 VINN.n211 4.5005
R72789 VINN.n338 VINN.n211 4.5005
R72790 VINN.n246 VINN.n211 4.5005
R72791 VINN.n340 VINN.n211 4.5005
R72792 VINN.n245 VINN.n211 4.5005
R72793 VINN.n342 VINN.n211 4.5005
R72794 VINN.n244 VINN.n211 4.5005
R72795 VINN.n344 VINN.n211 4.5005
R72796 VINN.n243 VINN.n211 4.5005
R72797 VINN.n346 VINN.n211 4.5005
R72798 VINN.n242 VINN.n211 4.5005
R72799 VINN.n348 VINN.n211 4.5005
R72800 VINN.n241 VINN.n211 4.5005
R72801 VINN.n350 VINN.n211 4.5005
R72802 VINN.n240 VINN.n211 4.5005
R72803 VINN.n352 VINN.n211 4.5005
R72804 VINN.n239 VINN.n211 4.5005
R72805 VINN.n354 VINN.n211 4.5005
R72806 VINN.n238 VINN.n211 4.5005
R72807 VINN.n356 VINN.n211 4.5005
R72808 VINN.n237 VINN.n211 4.5005
R72809 VINN.n358 VINN.n211 4.5005
R72810 VINN.n236 VINN.n211 4.5005
R72811 VINN.n360 VINN.n211 4.5005
R72812 VINN.n235 VINN.n211 4.5005
R72813 VINN.n362 VINN.n211 4.5005
R72814 VINN.n234 VINN.n211 4.5005
R72815 VINN.n364 VINN.n211 4.5005
R72816 VINN.n233 VINN.n211 4.5005
R72817 VINN.n366 VINN.n211 4.5005
R72818 VINN.n232 VINN.n211 4.5005
R72819 VINN.n368 VINN.n211 4.5005
R72820 VINN.n231 VINN.n211 4.5005
R72821 VINN.n370 VINN.n211 4.5005
R72822 VINN.n230 VINN.n211 4.5005
R72823 VINN.n372 VINN.n211 4.5005
R72824 VINN.n229 VINN.n211 4.5005
R72825 VINN.n374 VINN.n211 4.5005
R72826 VINN.n228 VINN.n211 4.5005
R72827 VINN.n376 VINN.n211 4.5005
R72828 VINN.n227 VINN.n211 4.5005
R72829 VINN.n378 VINN.n211 4.5005
R72830 VINN.n226 VINN.n211 4.5005
R72831 VINN.n380 VINN.n211 4.5005
R72832 VINN.n225 VINN.n211 4.5005
R72833 VINN.n382 VINN.n211 4.5005
R72834 VINN.n224 VINN.n211 4.5005
R72835 VINN.n384 VINN.n211 4.5005
R72836 VINN.n223 VINN.n211 4.5005
R72837 VINN.n386 VINN.n211 4.5005
R72838 VINN.n222 VINN.n211 4.5005
R72839 VINN.n388 VINN.n211 4.5005
R72840 VINN.n221 VINN.n211 4.5005
R72841 VINN.n390 VINN.n211 4.5005
R72842 VINN.n220 VINN.n211 4.5005
R72843 VINN.n392 VINN.n211 4.5005
R72844 VINN.n219 VINN.n211 4.5005
R72845 VINN.n394 VINN.n211 4.5005
R72846 VINN.n218 VINN.n211 4.5005
R72847 VINN.n396 VINN.n211 4.5005
R72848 VINN.n217 VINN.n211 4.5005
R72849 VINN.n398 VINN.n211 4.5005
R72850 VINN.n216 VINN.n211 4.5005
R72851 VINN.n400 VINN.n211 4.5005
R72852 VINN.n215 VINN.n211 4.5005
R72853 VINN.n654 VINN.n211 4.5005
R72854 VINN.n656 VINN.n211 4.5005
R72855 VINN.n211 VINN.n0 4.5005
R72856 VINN.n278 VINN.n89 4.5005
R72857 VINN.n276 VINN.n89 4.5005
R72858 VINN.n280 VINN.n89 4.5005
R72859 VINN.n275 VINN.n89 4.5005
R72860 VINN.n282 VINN.n89 4.5005
R72861 VINN.n274 VINN.n89 4.5005
R72862 VINN.n284 VINN.n89 4.5005
R72863 VINN.n273 VINN.n89 4.5005
R72864 VINN.n286 VINN.n89 4.5005
R72865 VINN.n272 VINN.n89 4.5005
R72866 VINN.n288 VINN.n89 4.5005
R72867 VINN.n271 VINN.n89 4.5005
R72868 VINN.n290 VINN.n89 4.5005
R72869 VINN.n270 VINN.n89 4.5005
R72870 VINN.n292 VINN.n89 4.5005
R72871 VINN.n269 VINN.n89 4.5005
R72872 VINN.n294 VINN.n89 4.5005
R72873 VINN.n268 VINN.n89 4.5005
R72874 VINN.n296 VINN.n89 4.5005
R72875 VINN.n267 VINN.n89 4.5005
R72876 VINN.n298 VINN.n89 4.5005
R72877 VINN.n266 VINN.n89 4.5005
R72878 VINN.n300 VINN.n89 4.5005
R72879 VINN.n265 VINN.n89 4.5005
R72880 VINN.n302 VINN.n89 4.5005
R72881 VINN.n264 VINN.n89 4.5005
R72882 VINN.n304 VINN.n89 4.5005
R72883 VINN.n263 VINN.n89 4.5005
R72884 VINN.n306 VINN.n89 4.5005
R72885 VINN.n262 VINN.n89 4.5005
R72886 VINN.n308 VINN.n89 4.5005
R72887 VINN.n261 VINN.n89 4.5005
R72888 VINN.n310 VINN.n89 4.5005
R72889 VINN.n260 VINN.n89 4.5005
R72890 VINN.n312 VINN.n89 4.5005
R72891 VINN.n259 VINN.n89 4.5005
R72892 VINN.n314 VINN.n89 4.5005
R72893 VINN.n258 VINN.n89 4.5005
R72894 VINN.n316 VINN.n89 4.5005
R72895 VINN.n257 VINN.n89 4.5005
R72896 VINN.n318 VINN.n89 4.5005
R72897 VINN.n256 VINN.n89 4.5005
R72898 VINN.n320 VINN.n89 4.5005
R72899 VINN.n255 VINN.n89 4.5005
R72900 VINN.n322 VINN.n89 4.5005
R72901 VINN.n254 VINN.n89 4.5005
R72902 VINN.n324 VINN.n89 4.5005
R72903 VINN.n253 VINN.n89 4.5005
R72904 VINN.n326 VINN.n89 4.5005
R72905 VINN.n252 VINN.n89 4.5005
R72906 VINN.n328 VINN.n89 4.5005
R72907 VINN.n251 VINN.n89 4.5005
R72908 VINN.n330 VINN.n89 4.5005
R72909 VINN.n250 VINN.n89 4.5005
R72910 VINN.n332 VINN.n89 4.5005
R72911 VINN.n249 VINN.n89 4.5005
R72912 VINN.n334 VINN.n89 4.5005
R72913 VINN.n248 VINN.n89 4.5005
R72914 VINN.n336 VINN.n89 4.5005
R72915 VINN.n247 VINN.n89 4.5005
R72916 VINN.n338 VINN.n89 4.5005
R72917 VINN.n246 VINN.n89 4.5005
R72918 VINN.n340 VINN.n89 4.5005
R72919 VINN.n245 VINN.n89 4.5005
R72920 VINN.n342 VINN.n89 4.5005
R72921 VINN.n244 VINN.n89 4.5005
R72922 VINN.n344 VINN.n89 4.5005
R72923 VINN.n243 VINN.n89 4.5005
R72924 VINN.n346 VINN.n89 4.5005
R72925 VINN.n242 VINN.n89 4.5005
R72926 VINN.n348 VINN.n89 4.5005
R72927 VINN.n241 VINN.n89 4.5005
R72928 VINN.n350 VINN.n89 4.5005
R72929 VINN.n240 VINN.n89 4.5005
R72930 VINN.n352 VINN.n89 4.5005
R72931 VINN.n239 VINN.n89 4.5005
R72932 VINN.n354 VINN.n89 4.5005
R72933 VINN.n238 VINN.n89 4.5005
R72934 VINN.n356 VINN.n89 4.5005
R72935 VINN.n237 VINN.n89 4.5005
R72936 VINN.n358 VINN.n89 4.5005
R72937 VINN.n236 VINN.n89 4.5005
R72938 VINN.n360 VINN.n89 4.5005
R72939 VINN.n235 VINN.n89 4.5005
R72940 VINN.n362 VINN.n89 4.5005
R72941 VINN.n234 VINN.n89 4.5005
R72942 VINN.n364 VINN.n89 4.5005
R72943 VINN.n233 VINN.n89 4.5005
R72944 VINN.n366 VINN.n89 4.5005
R72945 VINN.n232 VINN.n89 4.5005
R72946 VINN.n368 VINN.n89 4.5005
R72947 VINN.n231 VINN.n89 4.5005
R72948 VINN.n370 VINN.n89 4.5005
R72949 VINN.n230 VINN.n89 4.5005
R72950 VINN.n372 VINN.n89 4.5005
R72951 VINN.n229 VINN.n89 4.5005
R72952 VINN.n374 VINN.n89 4.5005
R72953 VINN.n228 VINN.n89 4.5005
R72954 VINN.n376 VINN.n89 4.5005
R72955 VINN.n227 VINN.n89 4.5005
R72956 VINN.n378 VINN.n89 4.5005
R72957 VINN.n226 VINN.n89 4.5005
R72958 VINN.n380 VINN.n89 4.5005
R72959 VINN.n225 VINN.n89 4.5005
R72960 VINN.n382 VINN.n89 4.5005
R72961 VINN.n224 VINN.n89 4.5005
R72962 VINN.n384 VINN.n89 4.5005
R72963 VINN.n223 VINN.n89 4.5005
R72964 VINN.n386 VINN.n89 4.5005
R72965 VINN.n222 VINN.n89 4.5005
R72966 VINN.n388 VINN.n89 4.5005
R72967 VINN.n221 VINN.n89 4.5005
R72968 VINN.n390 VINN.n89 4.5005
R72969 VINN.n220 VINN.n89 4.5005
R72970 VINN.n392 VINN.n89 4.5005
R72971 VINN.n219 VINN.n89 4.5005
R72972 VINN.n394 VINN.n89 4.5005
R72973 VINN.n218 VINN.n89 4.5005
R72974 VINN.n396 VINN.n89 4.5005
R72975 VINN.n217 VINN.n89 4.5005
R72976 VINN.n398 VINN.n89 4.5005
R72977 VINN.n216 VINN.n89 4.5005
R72978 VINN.n400 VINN.n89 4.5005
R72979 VINN.n215 VINN.n89 4.5005
R72980 VINN.n654 VINN.n89 4.5005
R72981 VINN.n656 VINN.n89 4.5005
R72982 VINN.n89 VINN.n0 4.5005
R72983 VINN.n278 VINN.n212 4.5005
R72984 VINN.n276 VINN.n212 4.5005
R72985 VINN.n280 VINN.n212 4.5005
R72986 VINN.n275 VINN.n212 4.5005
R72987 VINN.n282 VINN.n212 4.5005
R72988 VINN.n274 VINN.n212 4.5005
R72989 VINN.n284 VINN.n212 4.5005
R72990 VINN.n273 VINN.n212 4.5005
R72991 VINN.n286 VINN.n212 4.5005
R72992 VINN.n272 VINN.n212 4.5005
R72993 VINN.n288 VINN.n212 4.5005
R72994 VINN.n271 VINN.n212 4.5005
R72995 VINN.n290 VINN.n212 4.5005
R72996 VINN.n270 VINN.n212 4.5005
R72997 VINN.n292 VINN.n212 4.5005
R72998 VINN.n269 VINN.n212 4.5005
R72999 VINN.n294 VINN.n212 4.5005
R73000 VINN.n268 VINN.n212 4.5005
R73001 VINN.n296 VINN.n212 4.5005
R73002 VINN.n267 VINN.n212 4.5005
R73003 VINN.n298 VINN.n212 4.5005
R73004 VINN.n266 VINN.n212 4.5005
R73005 VINN.n300 VINN.n212 4.5005
R73006 VINN.n265 VINN.n212 4.5005
R73007 VINN.n302 VINN.n212 4.5005
R73008 VINN.n264 VINN.n212 4.5005
R73009 VINN.n304 VINN.n212 4.5005
R73010 VINN.n263 VINN.n212 4.5005
R73011 VINN.n306 VINN.n212 4.5005
R73012 VINN.n262 VINN.n212 4.5005
R73013 VINN.n308 VINN.n212 4.5005
R73014 VINN.n261 VINN.n212 4.5005
R73015 VINN.n310 VINN.n212 4.5005
R73016 VINN.n260 VINN.n212 4.5005
R73017 VINN.n312 VINN.n212 4.5005
R73018 VINN.n259 VINN.n212 4.5005
R73019 VINN.n314 VINN.n212 4.5005
R73020 VINN.n258 VINN.n212 4.5005
R73021 VINN.n316 VINN.n212 4.5005
R73022 VINN.n257 VINN.n212 4.5005
R73023 VINN.n318 VINN.n212 4.5005
R73024 VINN.n256 VINN.n212 4.5005
R73025 VINN.n320 VINN.n212 4.5005
R73026 VINN.n255 VINN.n212 4.5005
R73027 VINN.n322 VINN.n212 4.5005
R73028 VINN.n254 VINN.n212 4.5005
R73029 VINN.n324 VINN.n212 4.5005
R73030 VINN.n253 VINN.n212 4.5005
R73031 VINN.n326 VINN.n212 4.5005
R73032 VINN.n252 VINN.n212 4.5005
R73033 VINN.n328 VINN.n212 4.5005
R73034 VINN.n251 VINN.n212 4.5005
R73035 VINN.n330 VINN.n212 4.5005
R73036 VINN.n250 VINN.n212 4.5005
R73037 VINN.n332 VINN.n212 4.5005
R73038 VINN.n249 VINN.n212 4.5005
R73039 VINN.n334 VINN.n212 4.5005
R73040 VINN.n248 VINN.n212 4.5005
R73041 VINN.n336 VINN.n212 4.5005
R73042 VINN.n247 VINN.n212 4.5005
R73043 VINN.n338 VINN.n212 4.5005
R73044 VINN.n246 VINN.n212 4.5005
R73045 VINN.n340 VINN.n212 4.5005
R73046 VINN.n245 VINN.n212 4.5005
R73047 VINN.n342 VINN.n212 4.5005
R73048 VINN.n244 VINN.n212 4.5005
R73049 VINN.n344 VINN.n212 4.5005
R73050 VINN.n243 VINN.n212 4.5005
R73051 VINN.n346 VINN.n212 4.5005
R73052 VINN.n242 VINN.n212 4.5005
R73053 VINN.n348 VINN.n212 4.5005
R73054 VINN.n241 VINN.n212 4.5005
R73055 VINN.n350 VINN.n212 4.5005
R73056 VINN.n240 VINN.n212 4.5005
R73057 VINN.n352 VINN.n212 4.5005
R73058 VINN.n239 VINN.n212 4.5005
R73059 VINN.n354 VINN.n212 4.5005
R73060 VINN.n238 VINN.n212 4.5005
R73061 VINN.n356 VINN.n212 4.5005
R73062 VINN.n237 VINN.n212 4.5005
R73063 VINN.n358 VINN.n212 4.5005
R73064 VINN.n236 VINN.n212 4.5005
R73065 VINN.n360 VINN.n212 4.5005
R73066 VINN.n235 VINN.n212 4.5005
R73067 VINN.n362 VINN.n212 4.5005
R73068 VINN.n234 VINN.n212 4.5005
R73069 VINN.n364 VINN.n212 4.5005
R73070 VINN.n233 VINN.n212 4.5005
R73071 VINN.n366 VINN.n212 4.5005
R73072 VINN.n232 VINN.n212 4.5005
R73073 VINN.n368 VINN.n212 4.5005
R73074 VINN.n231 VINN.n212 4.5005
R73075 VINN.n370 VINN.n212 4.5005
R73076 VINN.n230 VINN.n212 4.5005
R73077 VINN.n372 VINN.n212 4.5005
R73078 VINN.n229 VINN.n212 4.5005
R73079 VINN.n374 VINN.n212 4.5005
R73080 VINN.n228 VINN.n212 4.5005
R73081 VINN.n376 VINN.n212 4.5005
R73082 VINN.n227 VINN.n212 4.5005
R73083 VINN.n378 VINN.n212 4.5005
R73084 VINN.n226 VINN.n212 4.5005
R73085 VINN.n380 VINN.n212 4.5005
R73086 VINN.n225 VINN.n212 4.5005
R73087 VINN.n382 VINN.n212 4.5005
R73088 VINN.n224 VINN.n212 4.5005
R73089 VINN.n384 VINN.n212 4.5005
R73090 VINN.n223 VINN.n212 4.5005
R73091 VINN.n386 VINN.n212 4.5005
R73092 VINN.n222 VINN.n212 4.5005
R73093 VINN.n388 VINN.n212 4.5005
R73094 VINN.n221 VINN.n212 4.5005
R73095 VINN.n390 VINN.n212 4.5005
R73096 VINN.n220 VINN.n212 4.5005
R73097 VINN.n392 VINN.n212 4.5005
R73098 VINN.n219 VINN.n212 4.5005
R73099 VINN.n394 VINN.n212 4.5005
R73100 VINN.n218 VINN.n212 4.5005
R73101 VINN.n396 VINN.n212 4.5005
R73102 VINN.n217 VINN.n212 4.5005
R73103 VINN.n398 VINN.n212 4.5005
R73104 VINN.n216 VINN.n212 4.5005
R73105 VINN.n400 VINN.n212 4.5005
R73106 VINN.n215 VINN.n212 4.5005
R73107 VINN.n654 VINN.n212 4.5005
R73108 VINN.n656 VINN.n212 4.5005
R73109 VINN.n212 VINN.n0 4.5005
R73110 VINN.n278 VINN.n88 4.5005
R73111 VINN.n276 VINN.n88 4.5005
R73112 VINN.n280 VINN.n88 4.5005
R73113 VINN.n275 VINN.n88 4.5005
R73114 VINN.n282 VINN.n88 4.5005
R73115 VINN.n274 VINN.n88 4.5005
R73116 VINN.n284 VINN.n88 4.5005
R73117 VINN.n273 VINN.n88 4.5005
R73118 VINN.n286 VINN.n88 4.5005
R73119 VINN.n272 VINN.n88 4.5005
R73120 VINN.n288 VINN.n88 4.5005
R73121 VINN.n271 VINN.n88 4.5005
R73122 VINN.n290 VINN.n88 4.5005
R73123 VINN.n270 VINN.n88 4.5005
R73124 VINN.n292 VINN.n88 4.5005
R73125 VINN.n269 VINN.n88 4.5005
R73126 VINN.n294 VINN.n88 4.5005
R73127 VINN.n268 VINN.n88 4.5005
R73128 VINN.n296 VINN.n88 4.5005
R73129 VINN.n267 VINN.n88 4.5005
R73130 VINN.n298 VINN.n88 4.5005
R73131 VINN.n266 VINN.n88 4.5005
R73132 VINN.n300 VINN.n88 4.5005
R73133 VINN.n265 VINN.n88 4.5005
R73134 VINN.n302 VINN.n88 4.5005
R73135 VINN.n264 VINN.n88 4.5005
R73136 VINN.n304 VINN.n88 4.5005
R73137 VINN.n263 VINN.n88 4.5005
R73138 VINN.n306 VINN.n88 4.5005
R73139 VINN.n262 VINN.n88 4.5005
R73140 VINN.n308 VINN.n88 4.5005
R73141 VINN.n261 VINN.n88 4.5005
R73142 VINN.n310 VINN.n88 4.5005
R73143 VINN.n260 VINN.n88 4.5005
R73144 VINN.n312 VINN.n88 4.5005
R73145 VINN.n259 VINN.n88 4.5005
R73146 VINN.n314 VINN.n88 4.5005
R73147 VINN.n258 VINN.n88 4.5005
R73148 VINN.n316 VINN.n88 4.5005
R73149 VINN.n257 VINN.n88 4.5005
R73150 VINN.n318 VINN.n88 4.5005
R73151 VINN.n256 VINN.n88 4.5005
R73152 VINN.n320 VINN.n88 4.5005
R73153 VINN.n255 VINN.n88 4.5005
R73154 VINN.n322 VINN.n88 4.5005
R73155 VINN.n254 VINN.n88 4.5005
R73156 VINN.n324 VINN.n88 4.5005
R73157 VINN.n253 VINN.n88 4.5005
R73158 VINN.n326 VINN.n88 4.5005
R73159 VINN.n252 VINN.n88 4.5005
R73160 VINN.n328 VINN.n88 4.5005
R73161 VINN.n251 VINN.n88 4.5005
R73162 VINN.n330 VINN.n88 4.5005
R73163 VINN.n250 VINN.n88 4.5005
R73164 VINN.n332 VINN.n88 4.5005
R73165 VINN.n249 VINN.n88 4.5005
R73166 VINN.n334 VINN.n88 4.5005
R73167 VINN.n248 VINN.n88 4.5005
R73168 VINN.n336 VINN.n88 4.5005
R73169 VINN.n247 VINN.n88 4.5005
R73170 VINN.n338 VINN.n88 4.5005
R73171 VINN.n246 VINN.n88 4.5005
R73172 VINN.n340 VINN.n88 4.5005
R73173 VINN.n245 VINN.n88 4.5005
R73174 VINN.n342 VINN.n88 4.5005
R73175 VINN.n244 VINN.n88 4.5005
R73176 VINN.n344 VINN.n88 4.5005
R73177 VINN.n243 VINN.n88 4.5005
R73178 VINN.n346 VINN.n88 4.5005
R73179 VINN.n242 VINN.n88 4.5005
R73180 VINN.n348 VINN.n88 4.5005
R73181 VINN.n241 VINN.n88 4.5005
R73182 VINN.n350 VINN.n88 4.5005
R73183 VINN.n240 VINN.n88 4.5005
R73184 VINN.n352 VINN.n88 4.5005
R73185 VINN.n239 VINN.n88 4.5005
R73186 VINN.n354 VINN.n88 4.5005
R73187 VINN.n238 VINN.n88 4.5005
R73188 VINN.n356 VINN.n88 4.5005
R73189 VINN.n237 VINN.n88 4.5005
R73190 VINN.n358 VINN.n88 4.5005
R73191 VINN.n236 VINN.n88 4.5005
R73192 VINN.n360 VINN.n88 4.5005
R73193 VINN.n235 VINN.n88 4.5005
R73194 VINN.n362 VINN.n88 4.5005
R73195 VINN.n234 VINN.n88 4.5005
R73196 VINN.n364 VINN.n88 4.5005
R73197 VINN.n233 VINN.n88 4.5005
R73198 VINN.n366 VINN.n88 4.5005
R73199 VINN.n232 VINN.n88 4.5005
R73200 VINN.n368 VINN.n88 4.5005
R73201 VINN.n231 VINN.n88 4.5005
R73202 VINN.n370 VINN.n88 4.5005
R73203 VINN.n230 VINN.n88 4.5005
R73204 VINN.n372 VINN.n88 4.5005
R73205 VINN.n229 VINN.n88 4.5005
R73206 VINN.n374 VINN.n88 4.5005
R73207 VINN.n228 VINN.n88 4.5005
R73208 VINN.n376 VINN.n88 4.5005
R73209 VINN.n227 VINN.n88 4.5005
R73210 VINN.n378 VINN.n88 4.5005
R73211 VINN.n226 VINN.n88 4.5005
R73212 VINN.n380 VINN.n88 4.5005
R73213 VINN.n225 VINN.n88 4.5005
R73214 VINN.n382 VINN.n88 4.5005
R73215 VINN.n224 VINN.n88 4.5005
R73216 VINN.n384 VINN.n88 4.5005
R73217 VINN.n223 VINN.n88 4.5005
R73218 VINN.n386 VINN.n88 4.5005
R73219 VINN.n222 VINN.n88 4.5005
R73220 VINN.n388 VINN.n88 4.5005
R73221 VINN.n221 VINN.n88 4.5005
R73222 VINN.n390 VINN.n88 4.5005
R73223 VINN.n220 VINN.n88 4.5005
R73224 VINN.n392 VINN.n88 4.5005
R73225 VINN.n219 VINN.n88 4.5005
R73226 VINN.n394 VINN.n88 4.5005
R73227 VINN.n218 VINN.n88 4.5005
R73228 VINN.n396 VINN.n88 4.5005
R73229 VINN.n217 VINN.n88 4.5005
R73230 VINN.n398 VINN.n88 4.5005
R73231 VINN.n216 VINN.n88 4.5005
R73232 VINN.n400 VINN.n88 4.5005
R73233 VINN.n215 VINN.n88 4.5005
R73234 VINN.n654 VINN.n88 4.5005
R73235 VINN.n656 VINN.n88 4.5005
R73236 VINN.n88 VINN.n0 4.5005
R73237 VINN.n278 VINN.n213 4.5005
R73238 VINN.n276 VINN.n213 4.5005
R73239 VINN.n280 VINN.n213 4.5005
R73240 VINN.n275 VINN.n213 4.5005
R73241 VINN.n282 VINN.n213 4.5005
R73242 VINN.n274 VINN.n213 4.5005
R73243 VINN.n284 VINN.n213 4.5005
R73244 VINN.n273 VINN.n213 4.5005
R73245 VINN.n286 VINN.n213 4.5005
R73246 VINN.n272 VINN.n213 4.5005
R73247 VINN.n288 VINN.n213 4.5005
R73248 VINN.n271 VINN.n213 4.5005
R73249 VINN.n290 VINN.n213 4.5005
R73250 VINN.n270 VINN.n213 4.5005
R73251 VINN.n292 VINN.n213 4.5005
R73252 VINN.n269 VINN.n213 4.5005
R73253 VINN.n294 VINN.n213 4.5005
R73254 VINN.n268 VINN.n213 4.5005
R73255 VINN.n296 VINN.n213 4.5005
R73256 VINN.n267 VINN.n213 4.5005
R73257 VINN.n298 VINN.n213 4.5005
R73258 VINN.n266 VINN.n213 4.5005
R73259 VINN.n300 VINN.n213 4.5005
R73260 VINN.n265 VINN.n213 4.5005
R73261 VINN.n302 VINN.n213 4.5005
R73262 VINN.n264 VINN.n213 4.5005
R73263 VINN.n304 VINN.n213 4.5005
R73264 VINN.n263 VINN.n213 4.5005
R73265 VINN.n306 VINN.n213 4.5005
R73266 VINN.n262 VINN.n213 4.5005
R73267 VINN.n308 VINN.n213 4.5005
R73268 VINN.n261 VINN.n213 4.5005
R73269 VINN.n310 VINN.n213 4.5005
R73270 VINN.n260 VINN.n213 4.5005
R73271 VINN.n312 VINN.n213 4.5005
R73272 VINN.n259 VINN.n213 4.5005
R73273 VINN.n314 VINN.n213 4.5005
R73274 VINN.n258 VINN.n213 4.5005
R73275 VINN.n316 VINN.n213 4.5005
R73276 VINN.n257 VINN.n213 4.5005
R73277 VINN.n318 VINN.n213 4.5005
R73278 VINN.n256 VINN.n213 4.5005
R73279 VINN.n320 VINN.n213 4.5005
R73280 VINN.n255 VINN.n213 4.5005
R73281 VINN.n322 VINN.n213 4.5005
R73282 VINN.n254 VINN.n213 4.5005
R73283 VINN.n324 VINN.n213 4.5005
R73284 VINN.n253 VINN.n213 4.5005
R73285 VINN.n326 VINN.n213 4.5005
R73286 VINN.n252 VINN.n213 4.5005
R73287 VINN.n328 VINN.n213 4.5005
R73288 VINN.n251 VINN.n213 4.5005
R73289 VINN.n330 VINN.n213 4.5005
R73290 VINN.n250 VINN.n213 4.5005
R73291 VINN.n332 VINN.n213 4.5005
R73292 VINN.n249 VINN.n213 4.5005
R73293 VINN.n334 VINN.n213 4.5005
R73294 VINN.n248 VINN.n213 4.5005
R73295 VINN.n336 VINN.n213 4.5005
R73296 VINN.n247 VINN.n213 4.5005
R73297 VINN.n338 VINN.n213 4.5005
R73298 VINN.n246 VINN.n213 4.5005
R73299 VINN.n340 VINN.n213 4.5005
R73300 VINN.n245 VINN.n213 4.5005
R73301 VINN.n342 VINN.n213 4.5005
R73302 VINN.n244 VINN.n213 4.5005
R73303 VINN.n344 VINN.n213 4.5005
R73304 VINN.n243 VINN.n213 4.5005
R73305 VINN.n346 VINN.n213 4.5005
R73306 VINN.n242 VINN.n213 4.5005
R73307 VINN.n348 VINN.n213 4.5005
R73308 VINN.n241 VINN.n213 4.5005
R73309 VINN.n350 VINN.n213 4.5005
R73310 VINN.n240 VINN.n213 4.5005
R73311 VINN.n352 VINN.n213 4.5005
R73312 VINN.n239 VINN.n213 4.5005
R73313 VINN.n354 VINN.n213 4.5005
R73314 VINN.n238 VINN.n213 4.5005
R73315 VINN.n356 VINN.n213 4.5005
R73316 VINN.n237 VINN.n213 4.5005
R73317 VINN.n358 VINN.n213 4.5005
R73318 VINN.n236 VINN.n213 4.5005
R73319 VINN.n360 VINN.n213 4.5005
R73320 VINN.n235 VINN.n213 4.5005
R73321 VINN.n362 VINN.n213 4.5005
R73322 VINN.n234 VINN.n213 4.5005
R73323 VINN.n364 VINN.n213 4.5005
R73324 VINN.n233 VINN.n213 4.5005
R73325 VINN.n366 VINN.n213 4.5005
R73326 VINN.n232 VINN.n213 4.5005
R73327 VINN.n368 VINN.n213 4.5005
R73328 VINN.n231 VINN.n213 4.5005
R73329 VINN.n370 VINN.n213 4.5005
R73330 VINN.n230 VINN.n213 4.5005
R73331 VINN.n372 VINN.n213 4.5005
R73332 VINN.n229 VINN.n213 4.5005
R73333 VINN.n374 VINN.n213 4.5005
R73334 VINN.n228 VINN.n213 4.5005
R73335 VINN.n376 VINN.n213 4.5005
R73336 VINN.n227 VINN.n213 4.5005
R73337 VINN.n378 VINN.n213 4.5005
R73338 VINN.n226 VINN.n213 4.5005
R73339 VINN.n380 VINN.n213 4.5005
R73340 VINN.n225 VINN.n213 4.5005
R73341 VINN.n382 VINN.n213 4.5005
R73342 VINN.n224 VINN.n213 4.5005
R73343 VINN.n384 VINN.n213 4.5005
R73344 VINN.n223 VINN.n213 4.5005
R73345 VINN.n386 VINN.n213 4.5005
R73346 VINN.n222 VINN.n213 4.5005
R73347 VINN.n388 VINN.n213 4.5005
R73348 VINN.n221 VINN.n213 4.5005
R73349 VINN.n390 VINN.n213 4.5005
R73350 VINN.n220 VINN.n213 4.5005
R73351 VINN.n392 VINN.n213 4.5005
R73352 VINN.n219 VINN.n213 4.5005
R73353 VINN.n394 VINN.n213 4.5005
R73354 VINN.n218 VINN.n213 4.5005
R73355 VINN.n396 VINN.n213 4.5005
R73356 VINN.n217 VINN.n213 4.5005
R73357 VINN.n398 VINN.n213 4.5005
R73358 VINN.n216 VINN.n213 4.5005
R73359 VINN.n400 VINN.n213 4.5005
R73360 VINN.n215 VINN.n213 4.5005
R73361 VINN.n654 VINN.n213 4.5005
R73362 VINN.n656 VINN.n213 4.5005
R73363 VINN.n213 VINN.n0 4.5005
R73364 VINN.n278 VINN.n87 4.5005
R73365 VINN.n276 VINN.n87 4.5005
R73366 VINN.n280 VINN.n87 4.5005
R73367 VINN.n275 VINN.n87 4.5005
R73368 VINN.n282 VINN.n87 4.5005
R73369 VINN.n274 VINN.n87 4.5005
R73370 VINN.n284 VINN.n87 4.5005
R73371 VINN.n273 VINN.n87 4.5005
R73372 VINN.n286 VINN.n87 4.5005
R73373 VINN.n272 VINN.n87 4.5005
R73374 VINN.n288 VINN.n87 4.5005
R73375 VINN.n271 VINN.n87 4.5005
R73376 VINN.n290 VINN.n87 4.5005
R73377 VINN.n270 VINN.n87 4.5005
R73378 VINN.n292 VINN.n87 4.5005
R73379 VINN.n269 VINN.n87 4.5005
R73380 VINN.n294 VINN.n87 4.5005
R73381 VINN.n268 VINN.n87 4.5005
R73382 VINN.n296 VINN.n87 4.5005
R73383 VINN.n267 VINN.n87 4.5005
R73384 VINN.n298 VINN.n87 4.5005
R73385 VINN.n266 VINN.n87 4.5005
R73386 VINN.n300 VINN.n87 4.5005
R73387 VINN.n265 VINN.n87 4.5005
R73388 VINN.n302 VINN.n87 4.5005
R73389 VINN.n264 VINN.n87 4.5005
R73390 VINN.n304 VINN.n87 4.5005
R73391 VINN.n263 VINN.n87 4.5005
R73392 VINN.n306 VINN.n87 4.5005
R73393 VINN.n262 VINN.n87 4.5005
R73394 VINN.n308 VINN.n87 4.5005
R73395 VINN.n261 VINN.n87 4.5005
R73396 VINN.n310 VINN.n87 4.5005
R73397 VINN.n260 VINN.n87 4.5005
R73398 VINN.n312 VINN.n87 4.5005
R73399 VINN.n259 VINN.n87 4.5005
R73400 VINN.n314 VINN.n87 4.5005
R73401 VINN.n258 VINN.n87 4.5005
R73402 VINN.n316 VINN.n87 4.5005
R73403 VINN.n257 VINN.n87 4.5005
R73404 VINN.n318 VINN.n87 4.5005
R73405 VINN.n256 VINN.n87 4.5005
R73406 VINN.n320 VINN.n87 4.5005
R73407 VINN.n255 VINN.n87 4.5005
R73408 VINN.n322 VINN.n87 4.5005
R73409 VINN.n254 VINN.n87 4.5005
R73410 VINN.n324 VINN.n87 4.5005
R73411 VINN.n253 VINN.n87 4.5005
R73412 VINN.n326 VINN.n87 4.5005
R73413 VINN.n252 VINN.n87 4.5005
R73414 VINN.n328 VINN.n87 4.5005
R73415 VINN.n251 VINN.n87 4.5005
R73416 VINN.n330 VINN.n87 4.5005
R73417 VINN.n250 VINN.n87 4.5005
R73418 VINN.n332 VINN.n87 4.5005
R73419 VINN.n249 VINN.n87 4.5005
R73420 VINN.n334 VINN.n87 4.5005
R73421 VINN.n248 VINN.n87 4.5005
R73422 VINN.n336 VINN.n87 4.5005
R73423 VINN.n247 VINN.n87 4.5005
R73424 VINN.n338 VINN.n87 4.5005
R73425 VINN.n246 VINN.n87 4.5005
R73426 VINN.n340 VINN.n87 4.5005
R73427 VINN.n245 VINN.n87 4.5005
R73428 VINN.n342 VINN.n87 4.5005
R73429 VINN.n244 VINN.n87 4.5005
R73430 VINN.n344 VINN.n87 4.5005
R73431 VINN.n243 VINN.n87 4.5005
R73432 VINN.n346 VINN.n87 4.5005
R73433 VINN.n242 VINN.n87 4.5005
R73434 VINN.n348 VINN.n87 4.5005
R73435 VINN.n241 VINN.n87 4.5005
R73436 VINN.n350 VINN.n87 4.5005
R73437 VINN.n240 VINN.n87 4.5005
R73438 VINN.n352 VINN.n87 4.5005
R73439 VINN.n239 VINN.n87 4.5005
R73440 VINN.n354 VINN.n87 4.5005
R73441 VINN.n238 VINN.n87 4.5005
R73442 VINN.n356 VINN.n87 4.5005
R73443 VINN.n237 VINN.n87 4.5005
R73444 VINN.n358 VINN.n87 4.5005
R73445 VINN.n236 VINN.n87 4.5005
R73446 VINN.n360 VINN.n87 4.5005
R73447 VINN.n235 VINN.n87 4.5005
R73448 VINN.n362 VINN.n87 4.5005
R73449 VINN.n234 VINN.n87 4.5005
R73450 VINN.n364 VINN.n87 4.5005
R73451 VINN.n233 VINN.n87 4.5005
R73452 VINN.n366 VINN.n87 4.5005
R73453 VINN.n232 VINN.n87 4.5005
R73454 VINN.n368 VINN.n87 4.5005
R73455 VINN.n231 VINN.n87 4.5005
R73456 VINN.n370 VINN.n87 4.5005
R73457 VINN.n230 VINN.n87 4.5005
R73458 VINN.n372 VINN.n87 4.5005
R73459 VINN.n229 VINN.n87 4.5005
R73460 VINN.n374 VINN.n87 4.5005
R73461 VINN.n228 VINN.n87 4.5005
R73462 VINN.n376 VINN.n87 4.5005
R73463 VINN.n227 VINN.n87 4.5005
R73464 VINN.n378 VINN.n87 4.5005
R73465 VINN.n226 VINN.n87 4.5005
R73466 VINN.n380 VINN.n87 4.5005
R73467 VINN.n225 VINN.n87 4.5005
R73468 VINN.n382 VINN.n87 4.5005
R73469 VINN.n224 VINN.n87 4.5005
R73470 VINN.n384 VINN.n87 4.5005
R73471 VINN.n223 VINN.n87 4.5005
R73472 VINN.n386 VINN.n87 4.5005
R73473 VINN.n222 VINN.n87 4.5005
R73474 VINN.n388 VINN.n87 4.5005
R73475 VINN.n221 VINN.n87 4.5005
R73476 VINN.n390 VINN.n87 4.5005
R73477 VINN.n220 VINN.n87 4.5005
R73478 VINN.n392 VINN.n87 4.5005
R73479 VINN.n219 VINN.n87 4.5005
R73480 VINN.n394 VINN.n87 4.5005
R73481 VINN.n218 VINN.n87 4.5005
R73482 VINN.n396 VINN.n87 4.5005
R73483 VINN.n217 VINN.n87 4.5005
R73484 VINN.n398 VINN.n87 4.5005
R73485 VINN.n216 VINN.n87 4.5005
R73486 VINN.n400 VINN.n87 4.5005
R73487 VINN.n215 VINN.n87 4.5005
R73488 VINN.n654 VINN.n87 4.5005
R73489 VINN.n656 VINN.n87 4.5005
R73490 VINN.n87 VINN.n0 4.5005
R73491 VINN.n655 VINN.n278 4.5005
R73492 VINN.n655 VINN.n276 4.5005
R73493 VINN.n655 VINN.n280 4.5005
R73494 VINN.n655 VINN.n275 4.5005
R73495 VINN.n655 VINN.n282 4.5005
R73496 VINN.n655 VINN.n274 4.5005
R73497 VINN.n655 VINN.n284 4.5005
R73498 VINN.n655 VINN.n273 4.5005
R73499 VINN.n655 VINN.n286 4.5005
R73500 VINN.n655 VINN.n272 4.5005
R73501 VINN.n655 VINN.n288 4.5005
R73502 VINN.n655 VINN.n271 4.5005
R73503 VINN.n655 VINN.n290 4.5005
R73504 VINN.n655 VINN.n270 4.5005
R73505 VINN.n655 VINN.n292 4.5005
R73506 VINN.n655 VINN.n269 4.5005
R73507 VINN.n655 VINN.n294 4.5005
R73508 VINN.n655 VINN.n268 4.5005
R73509 VINN.n655 VINN.n296 4.5005
R73510 VINN.n655 VINN.n267 4.5005
R73511 VINN.n655 VINN.n298 4.5005
R73512 VINN.n655 VINN.n266 4.5005
R73513 VINN.n655 VINN.n300 4.5005
R73514 VINN.n655 VINN.n265 4.5005
R73515 VINN.n655 VINN.n302 4.5005
R73516 VINN.n655 VINN.n264 4.5005
R73517 VINN.n655 VINN.n304 4.5005
R73518 VINN.n655 VINN.n263 4.5005
R73519 VINN.n655 VINN.n306 4.5005
R73520 VINN.n655 VINN.n262 4.5005
R73521 VINN.n655 VINN.n308 4.5005
R73522 VINN.n655 VINN.n261 4.5005
R73523 VINN.n655 VINN.n310 4.5005
R73524 VINN.n655 VINN.n260 4.5005
R73525 VINN.n655 VINN.n312 4.5005
R73526 VINN.n655 VINN.n259 4.5005
R73527 VINN.n655 VINN.n314 4.5005
R73528 VINN.n655 VINN.n258 4.5005
R73529 VINN.n655 VINN.n316 4.5005
R73530 VINN.n655 VINN.n257 4.5005
R73531 VINN.n655 VINN.n318 4.5005
R73532 VINN.n655 VINN.n256 4.5005
R73533 VINN.n655 VINN.n320 4.5005
R73534 VINN.n655 VINN.n255 4.5005
R73535 VINN.n655 VINN.n322 4.5005
R73536 VINN.n655 VINN.n254 4.5005
R73537 VINN.n655 VINN.n324 4.5005
R73538 VINN.n655 VINN.n253 4.5005
R73539 VINN.n655 VINN.n326 4.5005
R73540 VINN.n655 VINN.n252 4.5005
R73541 VINN.n655 VINN.n328 4.5005
R73542 VINN.n655 VINN.n251 4.5005
R73543 VINN.n655 VINN.n330 4.5005
R73544 VINN.n655 VINN.n250 4.5005
R73545 VINN.n655 VINN.n332 4.5005
R73546 VINN.n655 VINN.n249 4.5005
R73547 VINN.n655 VINN.n334 4.5005
R73548 VINN.n655 VINN.n248 4.5005
R73549 VINN.n655 VINN.n336 4.5005
R73550 VINN.n655 VINN.n247 4.5005
R73551 VINN.n655 VINN.n338 4.5005
R73552 VINN.n655 VINN.n246 4.5005
R73553 VINN.n655 VINN.n340 4.5005
R73554 VINN.n655 VINN.n245 4.5005
R73555 VINN.n655 VINN.n342 4.5005
R73556 VINN.n655 VINN.n244 4.5005
R73557 VINN.n655 VINN.n344 4.5005
R73558 VINN.n655 VINN.n243 4.5005
R73559 VINN.n655 VINN.n346 4.5005
R73560 VINN.n655 VINN.n242 4.5005
R73561 VINN.n655 VINN.n348 4.5005
R73562 VINN.n655 VINN.n241 4.5005
R73563 VINN.n655 VINN.n350 4.5005
R73564 VINN.n655 VINN.n240 4.5005
R73565 VINN.n655 VINN.n352 4.5005
R73566 VINN.n655 VINN.n239 4.5005
R73567 VINN.n655 VINN.n354 4.5005
R73568 VINN.n655 VINN.n238 4.5005
R73569 VINN.n655 VINN.n356 4.5005
R73570 VINN.n655 VINN.n237 4.5005
R73571 VINN.n655 VINN.n358 4.5005
R73572 VINN.n655 VINN.n236 4.5005
R73573 VINN.n655 VINN.n360 4.5005
R73574 VINN.n655 VINN.n235 4.5005
R73575 VINN.n655 VINN.n362 4.5005
R73576 VINN.n655 VINN.n234 4.5005
R73577 VINN.n655 VINN.n364 4.5005
R73578 VINN.n655 VINN.n233 4.5005
R73579 VINN.n655 VINN.n366 4.5005
R73580 VINN.n655 VINN.n232 4.5005
R73581 VINN.n655 VINN.n368 4.5005
R73582 VINN.n655 VINN.n231 4.5005
R73583 VINN.n655 VINN.n370 4.5005
R73584 VINN.n655 VINN.n230 4.5005
R73585 VINN.n655 VINN.n372 4.5005
R73586 VINN.n655 VINN.n229 4.5005
R73587 VINN.n655 VINN.n374 4.5005
R73588 VINN.n655 VINN.n228 4.5005
R73589 VINN.n655 VINN.n376 4.5005
R73590 VINN.n655 VINN.n227 4.5005
R73591 VINN.n655 VINN.n378 4.5005
R73592 VINN.n655 VINN.n226 4.5005
R73593 VINN.n655 VINN.n380 4.5005
R73594 VINN.n655 VINN.n225 4.5005
R73595 VINN.n655 VINN.n382 4.5005
R73596 VINN.n655 VINN.n224 4.5005
R73597 VINN.n655 VINN.n384 4.5005
R73598 VINN.n655 VINN.n223 4.5005
R73599 VINN.n655 VINN.n386 4.5005
R73600 VINN.n655 VINN.n222 4.5005
R73601 VINN.n655 VINN.n388 4.5005
R73602 VINN.n655 VINN.n221 4.5005
R73603 VINN.n655 VINN.n390 4.5005
R73604 VINN.n655 VINN.n220 4.5005
R73605 VINN.n655 VINN.n392 4.5005
R73606 VINN.n655 VINN.n219 4.5005
R73607 VINN.n655 VINN.n394 4.5005
R73608 VINN.n655 VINN.n218 4.5005
R73609 VINN.n655 VINN.n396 4.5005
R73610 VINN.n655 VINN.n217 4.5005
R73611 VINN.n655 VINN.n398 4.5005
R73612 VINN.n655 VINN.n216 4.5005
R73613 VINN.n655 VINN.n400 4.5005
R73614 VINN.n655 VINN.n215 4.5005
R73615 VINN.n655 VINN.n654 4.5005
R73616 VINN.n656 VINN.n655 4.5005
R73617 VINN.n655 VINN.n0 4.5005
R73618 VINN.n278 VINN.n86 4.5005
R73619 VINN.n276 VINN.n86 4.5005
R73620 VINN.n280 VINN.n86 4.5005
R73621 VINN.n275 VINN.n86 4.5005
R73622 VINN.n282 VINN.n86 4.5005
R73623 VINN.n274 VINN.n86 4.5005
R73624 VINN.n284 VINN.n86 4.5005
R73625 VINN.n273 VINN.n86 4.5005
R73626 VINN.n286 VINN.n86 4.5005
R73627 VINN.n272 VINN.n86 4.5005
R73628 VINN.n288 VINN.n86 4.5005
R73629 VINN.n271 VINN.n86 4.5005
R73630 VINN.n290 VINN.n86 4.5005
R73631 VINN.n270 VINN.n86 4.5005
R73632 VINN.n292 VINN.n86 4.5005
R73633 VINN.n269 VINN.n86 4.5005
R73634 VINN.n294 VINN.n86 4.5005
R73635 VINN.n268 VINN.n86 4.5005
R73636 VINN.n296 VINN.n86 4.5005
R73637 VINN.n267 VINN.n86 4.5005
R73638 VINN.n298 VINN.n86 4.5005
R73639 VINN.n266 VINN.n86 4.5005
R73640 VINN.n300 VINN.n86 4.5005
R73641 VINN.n265 VINN.n86 4.5005
R73642 VINN.n302 VINN.n86 4.5005
R73643 VINN.n264 VINN.n86 4.5005
R73644 VINN.n304 VINN.n86 4.5005
R73645 VINN.n263 VINN.n86 4.5005
R73646 VINN.n306 VINN.n86 4.5005
R73647 VINN.n262 VINN.n86 4.5005
R73648 VINN.n308 VINN.n86 4.5005
R73649 VINN.n261 VINN.n86 4.5005
R73650 VINN.n310 VINN.n86 4.5005
R73651 VINN.n260 VINN.n86 4.5005
R73652 VINN.n312 VINN.n86 4.5005
R73653 VINN.n259 VINN.n86 4.5005
R73654 VINN.n314 VINN.n86 4.5005
R73655 VINN.n258 VINN.n86 4.5005
R73656 VINN.n316 VINN.n86 4.5005
R73657 VINN.n257 VINN.n86 4.5005
R73658 VINN.n318 VINN.n86 4.5005
R73659 VINN.n256 VINN.n86 4.5005
R73660 VINN.n320 VINN.n86 4.5005
R73661 VINN.n255 VINN.n86 4.5005
R73662 VINN.n322 VINN.n86 4.5005
R73663 VINN.n254 VINN.n86 4.5005
R73664 VINN.n324 VINN.n86 4.5005
R73665 VINN.n253 VINN.n86 4.5005
R73666 VINN.n326 VINN.n86 4.5005
R73667 VINN.n252 VINN.n86 4.5005
R73668 VINN.n328 VINN.n86 4.5005
R73669 VINN.n251 VINN.n86 4.5005
R73670 VINN.n330 VINN.n86 4.5005
R73671 VINN.n250 VINN.n86 4.5005
R73672 VINN.n332 VINN.n86 4.5005
R73673 VINN.n249 VINN.n86 4.5005
R73674 VINN.n334 VINN.n86 4.5005
R73675 VINN.n248 VINN.n86 4.5005
R73676 VINN.n336 VINN.n86 4.5005
R73677 VINN.n247 VINN.n86 4.5005
R73678 VINN.n338 VINN.n86 4.5005
R73679 VINN.n246 VINN.n86 4.5005
R73680 VINN.n340 VINN.n86 4.5005
R73681 VINN.n245 VINN.n86 4.5005
R73682 VINN.n342 VINN.n86 4.5005
R73683 VINN.n244 VINN.n86 4.5005
R73684 VINN.n344 VINN.n86 4.5005
R73685 VINN.n243 VINN.n86 4.5005
R73686 VINN.n346 VINN.n86 4.5005
R73687 VINN.n242 VINN.n86 4.5005
R73688 VINN.n348 VINN.n86 4.5005
R73689 VINN.n241 VINN.n86 4.5005
R73690 VINN.n350 VINN.n86 4.5005
R73691 VINN.n240 VINN.n86 4.5005
R73692 VINN.n352 VINN.n86 4.5005
R73693 VINN.n239 VINN.n86 4.5005
R73694 VINN.n354 VINN.n86 4.5005
R73695 VINN.n238 VINN.n86 4.5005
R73696 VINN.n356 VINN.n86 4.5005
R73697 VINN.n237 VINN.n86 4.5005
R73698 VINN.n358 VINN.n86 4.5005
R73699 VINN.n236 VINN.n86 4.5005
R73700 VINN.n360 VINN.n86 4.5005
R73701 VINN.n235 VINN.n86 4.5005
R73702 VINN.n362 VINN.n86 4.5005
R73703 VINN.n234 VINN.n86 4.5005
R73704 VINN.n364 VINN.n86 4.5005
R73705 VINN.n233 VINN.n86 4.5005
R73706 VINN.n366 VINN.n86 4.5005
R73707 VINN.n232 VINN.n86 4.5005
R73708 VINN.n368 VINN.n86 4.5005
R73709 VINN.n231 VINN.n86 4.5005
R73710 VINN.n370 VINN.n86 4.5005
R73711 VINN.n230 VINN.n86 4.5005
R73712 VINN.n372 VINN.n86 4.5005
R73713 VINN.n229 VINN.n86 4.5005
R73714 VINN.n374 VINN.n86 4.5005
R73715 VINN.n228 VINN.n86 4.5005
R73716 VINN.n376 VINN.n86 4.5005
R73717 VINN.n227 VINN.n86 4.5005
R73718 VINN.n378 VINN.n86 4.5005
R73719 VINN.n226 VINN.n86 4.5005
R73720 VINN.n380 VINN.n86 4.5005
R73721 VINN.n225 VINN.n86 4.5005
R73722 VINN.n382 VINN.n86 4.5005
R73723 VINN.n224 VINN.n86 4.5005
R73724 VINN.n384 VINN.n86 4.5005
R73725 VINN.n223 VINN.n86 4.5005
R73726 VINN.n386 VINN.n86 4.5005
R73727 VINN.n222 VINN.n86 4.5005
R73728 VINN.n388 VINN.n86 4.5005
R73729 VINN.n221 VINN.n86 4.5005
R73730 VINN.n390 VINN.n86 4.5005
R73731 VINN.n220 VINN.n86 4.5005
R73732 VINN.n392 VINN.n86 4.5005
R73733 VINN.n219 VINN.n86 4.5005
R73734 VINN.n394 VINN.n86 4.5005
R73735 VINN.n218 VINN.n86 4.5005
R73736 VINN.n396 VINN.n86 4.5005
R73737 VINN.n217 VINN.n86 4.5005
R73738 VINN.n398 VINN.n86 4.5005
R73739 VINN.n216 VINN.n86 4.5005
R73740 VINN.n400 VINN.n86 4.5005
R73741 VINN.n215 VINN.n86 4.5005
R73742 VINN.n654 VINN.n86 4.5005
R73743 VINN.n528 VINN.n86 4.5005
R73744 VINN.n656 VINN.n86 4.5005
R73745 VINN.n86 VINN.n0 4.5005
R73746 VINN.n462 VINN.n278 2.25083
R73747 VINN.n463 VINN.n461 2.25083
R73748 VINN.n463 VINN.n460 2.25083
R73749 VINN.n463 VINN.n459 2.25083
R73750 VINN.n463 VINN.n458 2.25083
R73751 VINN.n463 VINN.n457 2.25083
R73752 VINN.n463 VINN.n456 2.25083
R73753 VINN.n463 VINN.n455 2.25083
R73754 VINN.n463 VINN.n454 2.25083
R73755 VINN.n463 VINN.n453 2.25083
R73756 VINN.n463 VINN.n452 2.25083
R73757 VINN.n463 VINN.n451 2.25083
R73758 VINN.n463 VINN.n450 2.25083
R73759 VINN.n463 VINN.n449 2.25083
R73760 VINN.n463 VINN.n448 2.25083
R73761 VINN.n463 VINN.n447 2.25083
R73762 VINN.n463 VINN.n446 2.25083
R73763 VINN.n463 VINN.n445 2.25083
R73764 VINN.n463 VINN.n444 2.25083
R73765 VINN.n463 VINN.n443 2.25083
R73766 VINN.n463 VINN.n442 2.25083
R73767 VINN.n463 VINN.n441 2.25083
R73768 VINN.n463 VINN.n440 2.25083
R73769 VINN.n463 VINN.n439 2.25083
R73770 VINN.n463 VINN.n438 2.25083
R73771 VINN.n463 VINN.n437 2.25083
R73772 VINN.n463 VINN.n436 2.25083
R73773 VINN.n463 VINN.n435 2.25083
R73774 VINN.n463 VINN.n434 2.25083
R73775 VINN.n463 VINN.n433 2.25083
R73776 VINN.n463 VINN.n432 2.25083
R73777 VINN.n463 VINN.n431 2.25083
R73778 VINN.n463 VINN.n430 2.25083
R73779 VINN.n463 VINN.n429 2.25083
R73780 VINN.n463 VINN.n428 2.25083
R73781 VINN.n463 VINN.n427 2.25083
R73782 VINN.n463 VINN.n426 2.25083
R73783 VINN.n463 VINN.n425 2.25083
R73784 VINN.n463 VINN.n424 2.25083
R73785 VINN.n463 VINN.n423 2.25083
R73786 VINN.n463 VINN.n422 2.25083
R73787 VINN.n463 VINN.n421 2.25083
R73788 VINN.n463 VINN.n420 2.25083
R73789 VINN.n463 VINN.n419 2.25083
R73790 VINN.n463 VINN.n418 2.25083
R73791 VINN.n463 VINN.n417 2.25083
R73792 VINN.n463 VINN.n416 2.25083
R73793 VINN.n463 VINN.n415 2.25083
R73794 VINN.n463 VINN.n414 2.25083
R73795 VINN.n463 VINN.n413 2.25083
R73796 VINN.n463 VINN.n412 2.25083
R73797 VINN.n463 VINN.n411 2.25083
R73798 VINN.n463 VINN.n410 2.25083
R73799 VINN.n463 VINN.n409 2.25083
R73800 VINN.n463 VINN.n408 2.25083
R73801 VINN.n463 VINN.n407 2.25083
R73802 VINN.n463 VINN.n406 2.25083
R73803 VINN.n463 VINN.n405 2.25083
R73804 VINN.n463 VINN.n404 2.25083
R73805 VINN.n463 VINN.n403 2.25083
R73806 VINN.n463 VINN.n402 2.25083
R73807 VINN.n463 VINN.n401 2.25083
R73808 VINN.n464 VINN.n463 2.25083
R73809 VINN.n463 VINN.n150 2.25083
R73810 VINN.n463 VINN.n66 2.25083
R73811 VINN.n279 VINN.n151 2.25083
R73812 VINN.n281 VINN.n151 2.25083
R73813 VINN.n283 VINN.n151 2.25083
R73814 VINN.n285 VINN.n151 2.25083
R73815 VINN.n287 VINN.n151 2.25083
R73816 VINN.n289 VINN.n151 2.25083
R73817 VINN.n291 VINN.n151 2.25083
R73818 VINN.n293 VINN.n151 2.25083
R73819 VINN.n295 VINN.n151 2.25083
R73820 VINN.n297 VINN.n151 2.25083
R73821 VINN.n299 VINN.n151 2.25083
R73822 VINN.n301 VINN.n151 2.25083
R73823 VINN.n303 VINN.n151 2.25083
R73824 VINN.n305 VINN.n151 2.25083
R73825 VINN.n307 VINN.n151 2.25083
R73826 VINN.n309 VINN.n151 2.25083
R73827 VINN.n311 VINN.n151 2.25083
R73828 VINN.n313 VINN.n151 2.25083
R73829 VINN.n315 VINN.n151 2.25083
R73830 VINN.n317 VINN.n151 2.25083
R73831 VINN.n319 VINN.n151 2.25083
R73832 VINN.n321 VINN.n151 2.25083
R73833 VINN.n323 VINN.n151 2.25083
R73834 VINN.n325 VINN.n151 2.25083
R73835 VINN.n327 VINN.n151 2.25083
R73836 VINN.n329 VINN.n151 2.25083
R73837 VINN.n331 VINN.n151 2.25083
R73838 VINN.n333 VINN.n151 2.25083
R73839 VINN.n335 VINN.n151 2.25083
R73840 VINN.n337 VINN.n151 2.25083
R73841 VINN.n339 VINN.n151 2.25083
R73842 VINN.n341 VINN.n151 2.25083
R73843 VINN.n343 VINN.n151 2.25083
R73844 VINN.n345 VINN.n151 2.25083
R73845 VINN.n347 VINN.n151 2.25083
R73846 VINN.n349 VINN.n151 2.25083
R73847 VINN.n351 VINN.n151 2.25083
R73848 VINN.n353 VINN.n151 2.25083
R73849 VINN.n355 VINN.n151 2.25083
R73850 VINN.n357 VINN.n151 2.25083
R73851 VINN.n359 VINN.n151 2.25083
R73852 VINN.n361 VINN.n151 2.25083
R73853 VINN.n363 VINN.n151 2.25083
R73854 VINN.n365 VINN.n151 2.25083
R73855 VINN.n367 VINN.n151 2.25083
R73856 VINN.n369 VINN.n151 2.25083
R73857 VINN.n371 VINN.n151 2.25083
R73858 VINN.n373 VINN.n151 2.25083
R73859 VINN.n375 VINN.n151 2.25083
R73860 VINN.n377 VINN.n151 2.25083
R73861 VINN.n379 VINN.n151 2.25083
R73862 VINN.n381 VINN.n151 2.25083
R73863 VINN.n383 VINN.n151 2.25083
R73864 VINN.n385 VINN.n151 2.25083
R73865 VINN.n387 VINN.n151 2.25083
R73866 VINN.n389 VINN.n151 2.25083
R73867 VINN.n391 VINN.n151 2.25083
R73868 VINN.n393 VINN.n151 2.25083
R73869 VINN.n395 VINN.n151 2.25083
R73870 VINN.n397 VINN.n151 2.25083
R73871 VINN.n399 VINN.n151 2.25083
R73872 VINN.n465 VINN.n151 2.25083
R73873 VINN.n277 VINN.n149 2.25083
R73874 VINN.n657 VINN.n65 2.25083
R73875 VINN.n528 VINN.n466 2.25083
R73876 VINN.n657 VINN.n64 2.25083
R73877 VINN.n528 VINN.n467 2.25083
R73878 VINN.n657 VINN.n63 2.25083
R73879 VINN.n528 VINN.n468 2.25083
R73880 VINN.n657 VINN.n62 2.25083
R73881 VINN.n528 VINN.n469 2.25083
R73882 VINN.n657 VINN.n61 2.25083
R73883 VINN.n528 VINN.n470 2.25083
R73884 VINN.n657 VINN.n60 2.25083
R73885 VINN.n528 VINN.n471 2.25083
R73886 VINN.n657 VINN.n59 2.25083
R73887 VINN.n528 VINN.n472 2.25083
R73888 VINN.n657 VINN.n58 2.25083
R73889 VINN.n528 VINN.n473 2.25083
R73890 VINN.n657 VINN.n57 2.25083
R73891 VINN.n528 VINN.n474 2.25083
R73892 VINN.n657 VINN.n56 2.25083
R73893 VINN.n528 VINN.n475 2.25083
R73894 VINN.n657 VINN.n55 2.25083
R73895 VINN.n528 VINN.n476 2.25083
R73896 VINN.n657 VINN.n54 2.25083
R73897 VINN.n528 VINN.n477 2.25083
R73898 VINN.n657 VINN.n53 2.25083
R73899 VINN.n528 VINN.n478 2.25083
R73900 VINN.n657 VINN.n52 2.25083
R73901 VINN.n528 VINN.n479 2.25083
R73902 VINN.n657 VINN.n51 2.25083
R73903 VINN.n528 VINN.n480 2.25083
R73904 VINN.n657 VINN.n50 2.25083
R73905 VINN.n528 VINN.n481 2.25083
R73906 VINN.n657 VINN.n49 2.25083
R73907 VINN.n528 VINN.n482 2.25083
R73908 VINN.n657 VINN.n48 2.25083
R73909 VINN.n528 VINN.n483 2.25083
R73910 VINN.n657 VINN.n47 2.25083
R73911 VINN.n528 VINN.n484 2.25083
R73912 VINN.n657 VINN.n46 2.25083
R73913 VINN.n528 VINN.n485 2.25083
R73914 VINN.n657 VINN.n45 2.25083
R73915 VINN.n528 VINN.n486 2.25083
R73916 VINN.n657 VINN.n44 2.25083
R73917 VINN.n528 VINN.n487 2.25083
R73918 VINN.n657 VINN.n43 2.25083
R73919 VINN.n528 VINN.n488 2.25083
R73920 VINN.n657 VINN.n42 2.25083
R73921 VINN.n528 VINN.n489 2.25083
R73922 VINN.n657 VINN.n41 2.25083
R73923 VINN.n528 VINN.n490 2.25083
R73924 VINN.n657 VINN.n40 2.25083
R73925 VINN.n528 VINN.n491 2.25083
R73926 VINN.n657 VINN.n39 2.25083
R73927 VINN.n528 VINN.n492 2.25083
R73928 VINN.n657 VINN.n38 2.25083
R73929 VINN.n528 VINN.n493 2.25083
R73930 VINN.n657 VINN.n37 2.25083
R73931 VINN.n528 VINN.n494 2.25083
R73932 VINN.n657 VINN.n36 2.25083
R73933 VINN.n528 VINN.n495 2.25083
R73934 VINN.n657 VINN.n35 2.25083
R73935 VINN.n528 VINN.n496 2.25083
R73936 VINN.n657 VINN.n34 2.25083
R73937 VINN.n528 VINN.n497 2.25083
R73938 VINN.n657 VINN.n33 2.25083
R73939 VINN.n528 VINN.n498 2.25083
R73940 VINN.n657 VINN.n32 2.25083
R73941 VINN.n528 VINN.n499 2.25083
R73942 VINN.n657 VINN.n31 2.25083
R73943 VINN.n528 VINN.n500 2.25083
R73944 VINN.n657 VINN.n30 2.25083
R73945 VINN.n528 VINN.n501 2.25083
R73946 VINN.n657 VINN.n29 2.25083
R73947 VINN.n528 VINN.n502 2.25083
R73948 VINN.n657 VINN.n28 2.25083
R73949 VINN.n528 VINN.n503 2.25083
R73950 VINN.n657 VINN.n27 2.25083
R73951 VINN.n528 VINN.n504 2.25083
R73952 VINN.n657 VINN.n26 2.25083
R73953 VINN.n528 VINN.n505 2.25083
R73954 VINN.n657 VINN.n25 2.25083
R73955 VINN.n528 VINN.n506 2.25083
R73956 VINN.n657 VINN.n24 2.25083
R73957 VINN.n528 VINN.n507 2.25083
R73958 VINN.n657 VINN.n23 2.25083
R73959 VINN.n528 VINN.n508 2.25083
R73960 VINN.n657 VINN.n22 2.25083
R73961 VINN.n528 VINN.n509 2.25083
R73962 VINN.n657 VINN.n21 2.25083
R73963 VINN.n528 VINN.n510 2.25083
R73964 VINN.n657 VINN.n20 2.25083
R73965 VINN.n528 VINN.n511 2.25083
R73966 VINN.n657 VINN.n19 2.25083
R73967 VINN.n528 VINN.n512 2.25083
R73968 VINN.n657 VINN.n18 2.25083
R73969 VINN.n528 VINN.n513 2.25083
R73970 VINN.n657 VINN.n17 2.25083
R73971 VINN.n528 VINN.n514 2.25083
R73972 VINN.n657 VINN.n16 2.25083
R73973 VINN.n528 VINN.n515 2.25083
R73974 VINN.n657 VINN.n15 2.25083
R73975 VINN.n528 VINN.n516 2.25083
R73976 VINN.n657 VINN.n14 2.25083
R73977 VINN.n528 VINN.n517 2.25083
R73978 VINN.n657 VINN.n13 2.25083
R73979 VINN.n528 VINN.n518 2.25083
R73980 VINN.n657 VINN.n12 2.25083
R73981 VINN.n528 VINN.n519 2.25083
R73982 VINN.n657 VINN.n11 2.25083
R73983 VINN.n528 VINN.n520 2.25083
R73984 VINN.n657 VINN.n10 2.25083
R73985 VINN.n528 VINN.n521 2.25083
R73986 VINN.n657 VINN.n9 2.25083
R73987 VINN.n528 VINN.n522 2.25083
R73988 VINN.n657 VINN.n8 2.25083
R73989 VINN.n528 VINN.n523 2.25083
R73990 VINN.n657 VINN.n7 2.25083
R73991 VINN.n528 VINN.n524 2.25083
R73992 VINN.n657 VINN.n6 2.25083
R73993 VINN.n528 VINN.n525 2.25083
R73994 VINN.n657 VINN.n5 2.25083
R73995 VINN.n528 VINN.n526 2.25083
R73996 VINN.n657 VINN.n4 2.25083
R73997 VINN.n528 VINN.n527 2.25083
R73998 VINN.n657 VINN.n3 2.25083
R73999 VINN.n528 VINN.n214 2.25083
R74000 VINN.n657 VINN.n2 2.25083
R74001 VINN.n68 VINN.n67 0.0986818
R74002 VINN.n69 VINN.n68 0.0986818
R74003 VINN.n70 VINN.n69 0.0986818
R74004 VINN.n71 VINN.n70 0.0986818
R74005 VINN.n72 VINN.n71 0.0986818
R74006 VINN.n73 VINN.n72 0.0986818
R74007 VINN.n74 VINN.n73 0.0986818
R74008 VINN.n75 VINN.n74 0.0986818
R74009 VINN.n76 VINN.n75 0.0986818
R74010 VINN.n77 VINN.n76 0.0986818
R74011 VINN.n78 VINN.n77 0.0986818
R74012 VINN.n79 VINN.n78 0.0986818
R74013 VINN.n80 VINN.n79 0.0986818
R74014 VINN.n81 VINN.n80 0.0986818
R74015 VINN.n82 VINN.n81 0.0986818
R74016 VINN.n83 VINN.n82 0.0986818
R74017 VINN.n84 VINN.n83 0.0986818
R74018 VINN.n85 VINN.n84 0.0985091
R74019 VINN.n658 VINN.n0 0.0358487
R74020 VINN.n530 VINN.n278 0.0358487
R74021 VINN.n658 VINN.n657 0.0353837
R74022 VINN.n656 VINN.n1 0.0353837
R74023 VINN.n529 VINN.n528 0.0353837
R74024 VINN.n654 VINN.n653 0.0353837
R74025 VINN.n652 VINN.n215 0.0353837
R74026 VINN.n651 VINN.n400 0.0353837
R74027 VINN.n650 VINN.n216 0.0353837
R74028 VINN.n649 VINN.n398 0.0353837
R74029 VINN.n648 VINN.n217 0.0353837
R74030 VINN.n647 VINN.n396 0.0353837
R74031 VINN.n646 VINN.n218 0.0353837
R74032 VINN.n645 VINN.n394 0.0353837
R74033 VINN.n644 VINN.n219 0.0353837
R74034 VINN.n643 VINN.n392 0.0353837
R74035 VINN.n642 VINN.n220 0.0353837
R74036 VINN.n641 VINN.n390 0.0353837
R74037 VINN.n640 VINN.n221 0.0353837
R74038 VINN.n639 VINN.n388 0.0353837
R74039 VINN.n638 VINN.n222 0.0353837
R74040 VINN.n637 VINN.n386 0.0353837
R74041 VINN.n636 VINN.n223 0.0353837
R74042 VINN.n635 VINN.n384 0.0353837
R74043 VINN.n634 VINN.n224 0.0353837
R74044 VINN.n633 VINN.n382 0.0353837
R74045 VINN.n632 VINN.n225 0.0353837
R74046 VINN.n631 VINN.n380 0.0353837
R74047 VINN.n630 VINN.n226 0.0353837
R74048 VINN.n629 VINN.n378 0.0353837
R74049 VINN.n628 VINN.n227 0.0353837
R74050 VINN.n627 VINN.n376 0.0353837
R74051 VINN.n626 VINN.n228 0.0353837
R74052 VINN.n625 VINN.n374 0.0353837
R74053 VINN.n624 VINN.n229 0.0353837
R74054 VINN.n623 VINN.n372 0.0353837
R74055 VINN.n622 VINN.n230 0.0353837
R74056 VINN.n621 VINN.n370 0.0353837
R74057 VINN.n620 VINN.n231 0.0353837
R74058 VINN.n619 VINN.n368 0.0353837
R74059 VINN.n618 VINN.n232 0.0353837
R74060 VINN.n617 VINN.n366 0.0353837
R74061 VINN.n616 VINN.n233 0.0353837
R74062 VINN.n615 VINN.n364 0.0353837
R74063 VINN.n614 VINN.n234 0.0353837
R74064 VINN.n613 VINN.n362 0.0353837
R74065 VINN.n612 VINN.n235 0.0353837
R74066 VINN.n611 VINN.n360 0.0353837
R74067 VINN.n610 VINN.n236 0.0353837
R74068 VINN.n609 VINN.n358 0.0353837
R74069 VINN.n608 VINN.n237 0.0353837
R74070 VINN.n607 VINN.n356 0.0353837
R74071 VINN.n606 VINN.n238 0.0353837
R74072 VINN.n605 VINN.n354 0.0353837
R74073 VINN.n604 VINN.n239 0.0353837
R74074 VINN.n603 VINN.n352 0.0353837
R74075 VINN.n602 VINN.n240 0.0353837
R74076 VINN.n601 VINN.n350 0.0353837
R74077 VINN.n600 VINN.n241 0.0353837
R74078 VINN.n599 VINN.n348 0.0353837
R74079 VINN.n598 VINN.n242 0.0353837
R74080 VINN.n597 VINN.n346 0.0353837
R74081 VINN.n596 VINN.n243 0.0353837
R74082 VINN.n595 VINN.n344 0.0353837
R74083 VINN.n594 VINN.n244 0.0353837
R74084 VINN.n593 VINN.n342 0.0353837
R74085 VINN.n592 VINN.n245 0.0353837
R74086 VINN.n591 VINN.n340 0.0353837
R74087 VINN.n590 VINN.n246 0.0353837
R74088 VINN.n589 VINN.n338 0.0353837
R74089 VINN.n588 VINN.n247 0.0353837
R74090 VINN.n587 VINN.n336 0.0353837
R74091 VINN.n586 VINN.n248 0.0353837
R74092 VINN.n585 VINN.n334 0.0353837
R74093 VINN.n584 VINN.n249 0.0353837
R74094 VINN.n583 VINN.n332 0.0353837
R74095 VINN.n582 VINN.n250 0.0353837
R74096 VINN.n581 VINN.n330 0.0353837
R74097 VINN.n580 VINN.n251 0.0353837
R74098 VINN.n579 VINN.n328 0.0353837
R74099 VINN.n578 VINN.n252 0.0353837
R74100 VINN.n577 VINN.n326 0.0353837
R74101 VINN.n576 VINN.n253 0.0353837
R74102 VINN.n575 VINN.n324 0.0353837
R74103 VINN.n574 VINN.n254 0.0353837
R74104 VINN.n573 VINN.n322 0.0353837
R74105 VINN.n572 VINN.n255 0.0353837
R74106 VINN.n571 VINN.n320 0.0353837
R74107 VINN.n570 VINN.n256 0.0353837
R74108 VINN.n569 VINN.n318 0.0353837
R74109 VINN.n568 VINN.n257 0.0353837
R74110 VINN.n567 VINN.n316 0.0353837
R74111 VINN.n566 VINN.n258 0.0353837
R74112 VINN.n565 VINN.n314 0.0353837
R74113 VINN.n564 VINN.n259 0.0353837
R74114 VINN.n563 VINN.n312 0.0353837
R74115 VINN.n562 VINN.n260 0.0353837
R74116 VINN.n561 VINN.n310 0.0353837
R74117 VINN.n560 VINN.n261 0.0353837
R74118 VINN.n559 VINN.n308 0.0353837
R74119 VINN.n558 VINN.n262 0.0353837
R74120 VINN.n557 VINN.n306 0.0353837
R74121 VINN.n556 VINN.n263 0.0353837
R74122 VINN.n555 VINN.n304 0.0353837
R74123 VINN.n554 VINN.n264 0.0353837
R74124 VINN.n553 VINN.n302 0.0353837
R74125 VINN.n552 VINN.n265 0.0353837
R74126 VINN.n551 VINN.n300 0.0353837
R74127 VINN.n550 VINN.n266 0.0353837
R74128 VINN.n549 VINN.n298 0.0353837
R74129 VINN.n548 VINN.n267 0.0353837
R74130 VINN.n547 VINN.n296 0.0353837
R74131 VINN.n546 VINN.n268 0.0353837
R74132 VINN.n545 VINN.n294 0.0353837
R74133 VINN.n544 VINN.n269 0.0353837
R74134 VINN.n543 VINN.n292 0.0353837
R74135 VINN.n542 VINN.n270 0.0353837
R74136 VINN.n541 VINN.n290 0.0353837
R74137 VINN.n540 VINN.n271 0.0353837
R74138 VINN.n539 VINN.n288 0.0353837
R74139 VINN.n538 VINN.n272 0.0353837
R74140 VINN.n537 VINN.n286 0.0353837
R74141 VINN.n536 VINN.n273 0.0353837
R74142 VINN.n535 VINN.n284 0.0353837
R74143 VINN.n534 VINN.n274 0.0353837
R74144 VINN.n533 VINN.n282 0.0353837
R74145 VINN.n532 VINN.n275 0.0353837
R74146 VINN.n531 VINN.n280 0.0353837
R74147 VINN.n530 VINN.n276 0.0353837
R74148 VINN.n463 VINN.n462 0.00134872
R74149 VINN.n149 VINN.n65 0.00134872
R74150 VINN.n466 VINN.n152 0.00134872
R74151 VINN.n148 VINN.n64 0.00134872
R74152 VINN.n467 VINN.n153 0.00134872
R74153 VINN.n147 VINN.n63 0.00134872
R74154 VINN.n468 VINN.n154 0.00134872
R74155 VINN.n146 VINN.n62 0.00134872
R74156 VINN.n469 VINN.n155 0.00134872
R74157 VINN.n145 VINN.n61 0.00134872
R74158 VINN.n470 VINN.n156 0.00134872
R74159 VINN.n144 VINN.n60 0.00134872
R74160 VINN.n471 VINN.n157 0.00134872
R74161 VINN.n143 VINN.n59 0.00134872
R74162 VINN.n472 VINN.n158 0.00134872
R74163 VINN.n142 VINN.n58 0.00134872
R74164 VINN.n473 VINN.n159 0.00134872
R74165 VINN.n141 VINN.n57 0.00134872
R74166 VINN.n474 VINN.n160 0.00134872
R74167 VINN.n140 VINN.n56 0.00134872
R74168 VINN.n475 VINN.n161 0.00134872
R74169 VINN.n139 VINN.n55 0.00134872
R74170 VINN.n476 VINN.n162 0.00134872
R74171 VINN.n138 VINN.n54 0.00134872
R74172 VINN.n477 VINN.n163 0.00134872
R74173 VINN.n137 VINN.n53 0.00134872
R74174 VINN.n478 VINN.n164 0.00134872
R74175 VINN.n136 VINN.n52 0.00134872
R74176 VINN.n479 VINN.n165 0.00134872
R74177 VINN.n135 VINN.n51 0.00134872
R74178 VINN.n480 VINN.n166 0.00134872
R74179 VINN.n134 VINN.n50 0.00134872
R74180 VINN.n481 VINN.n167 0.00134872
R74181 VINN.n133 VINN.n49 0.00134872
R74182 VINN.n482 VINN.n168 0.00134872
R74183 VINN.n132 VINN.n48 0.00134872
R74184 VINN.n483 VINN.n169 0.00134872
R74185 VINN.n131 VINN.n47 0.00134872
R74186 VINN.n484 VINN.n170 0.00134872
R74187 VINN.n130 VINN.n46 0.00134872
R74188 VINN.n485 VINN.n171 0.00134872
R74189 VINN.n129 VINN.n45 0.00134872
R74190 VINN.n486 VINN.n172 0.00134872
R74191 VINN.n128 VINN.n44 0.00134872
R74192 VINN.n487 VINN.n173 0.00134872
R74193 VINN.n127 VINN.n43 0.00134872
R74194 VINN.n488 VINN.n174 0.00134872
R74195 VINN.n126 VINN.n42 0.00134872
R74196 VINN.n489 VINN.n175 0.00134872
R74197 VINN.n125 VINN.n41 0.00134872
R74198 VINN.n490 VINN.n176 0.00134872
R74199 VINN.n124 VINN.n40 0.00134872
R74200 VINN.n491 VINN.n177 0.00134872
R74201 VINN.n123 VINN.n39 0.00134872
R74202 VINN.n492 VINN.n178 0.00134872
R74203 VINN.n122 VINN.n38 0.00134872
R74204 VINN.n493 VINN.n179 0.00134872
R74205 VINN.n121 VINN.n37 0.00134872
R74206 VINN.n494 VINN.n180 0.00134872
R74207 VINN.n120 VINN.n36 0.00134872
R74208 VINN.n495 VINN.n181 0.00134872
R74209 VINN.n119 VINN.n35 0.00134872
R74210 VINN.n496 VINN.n182 0.00134872
R74211 VINN.n118 VINN.n34 0.00134872
R74212 VINN.n497 VINN.n183 0.00134872
R74213 VINN.n117 VINN.n33 0.00134872
R74214 VINN.n498 VINN.n184 0.00134872
R74215 VINN.n116 VINN.n32 0.00134872
R74216 VINN.n499 VINN.n185 0.00134872
R74217 VINN.n115 VINN.n31 0.00134872
R74218 VINN.n500 VINN.n186 0.00134872
R74219 VINN.n114 VINN.n30 0.00134872
R74220 VINN.n501 VINN.n187 0.00134872
R74221 VINN.n113 VINN.n29 0.00134872
R74222 VINN.n502 VINN.n188 0.00134872
R74223 VINN.n112 VINN.n28 0.00134872
R74224 VINN.n503 VINN.n189 0.00134872
R74225 VINN.n111 VINN.n27 0.00134872
R74226 VINN.n504 VINN.n190 0.00134872
R74227 VINN.n110 VINN.n26 0.00134872
R74228 VINN.n505 VINN.n191 0.00134872
R74229 VINN.n109 VINN.n25 0.00134872
R74230 VINN.n506 VINN.n192 0.00134872
R74231 VINN.n108 VINN.n24 0.00134872
R74232 VINN.n507 VINN.n193 0.00134872
R74233 VINN.n107 VINN.n23 0.00134872
R74234 VINN.n508 VINN.n194 0.00134872
R74235 VINN.n106 VINN.n22 0.00134872
R74236 VINN.n509 VINN.n195 0.00134872
R74237 VINN.n105 VINN.n21 0.00134872
R74238 VINN.n510 VINN.n196 0.00134872
R74239 VINN.n104 VINN.n20 0.00134872
R74240 VINN.n511 VINN.n197 0.00134872
R74241 VINN.n103 VINN.n19 0.00134872
R74242 VINN.n512 VINN.n198 0.00134872
R74243 VINN.n102 VINN.n18 0.00134872
R74244 VINN.n513 VINN.n199 0.00134872
R74245 VINN.n101 VINN.n17 0.00134872
R74246 VINN.n514 VINN.n200 0.00134872
R74247 VINN.n100 VINN.n16 0.00134872
R74248 VINN.n515 VINN.n201 0.00134872
R74249 VINN.n99 VINN.n15 0.00134872
R74250 VINN.n516 VINN.n202 0.00134872
R74251 VINN.n98 VINN.n14 0.00134872
R74252 VINN.n517 VINN.n203 0.00134872
R74253 VINN.n97 VINN.n13 0.00134872
R74254 VINN.n518 VINN.n204 0.00134872
R74255 VINN.n96 VINN.n12 0.00134872
R74256 VINN.n519 VINN.n205 0.00134872
R74257 VINN.n95 VINN.n11 0.00134872
R74258 VINN.n520 VINN.n206 0.00134872
R74259 VINN.n94 VINN.n10 0.00134872
R74260 VINN.n521 VINN.n207 0.00134872
R74261 VINN.n93 VINN.n9 0.00134872
R74262 VINN.n522 VINN.n208 0.00134872
R74263 VINN.n92 VINN.n8 0.00134872
R74264 VINN.n523 VINN.n209 0.00134872
R74265 VINN.n91 VINN.n7 0.00134872
R74266 VINN.n524 VINN.n210 0.00134872
R74267 VINN.n90 VINN.n6 0.00134872
R74268 VINN.n525 VINN.n211 0.00134872
R74269 VINN.n89 VINN.n5 0.00134872
R74270 VINN.n526 VINN.n212 0.00134872
R74271 VINN.n88 VINN.n4 0.00134872
R74272 VINN.n527 VINN.n213 0.00134872
R74273 VINN.n87 VINN.n3 0.00134872
R74274 VINN.n655 VINN.n214 0.00134872
R74275 VINN.n86 VINN.n2 0.00134872
R74276 VINN.n66 VINN.n0 0.00134872
R74277 VINN.n656 VINN.n150 0.00134872
R74278 VINN.n528 VINN.n465 0.00134872
R74279 VINN.n654 VINN.n464 0.00134872
R74280 VINN.n399 VINN.n215 0.00134872
R74281 VINN.n401 VINN.n400 0.00134872
R74282 VINN.n397 VINN.n216 0.00134872
R74283 VINN.n402 VINN.n398 0.00134872
R74284 VINN.n395 VINN.n217 0.00134872
R74285 VINN.n403 VINN.n396 0.00134872
R74286 VINN.n393 VINN.n218 0.00134872
R74287 VINN.n404 VINN.n394 0.00134872
R74288 VINN.n391 VINN.n219 0.00134872
R74289 VINN.n405 VINN.n392 0.00134872
R74290 VINN.n389 VINN.n220 0.00134872
R74291 VINN.n406 VINN.n390 0.00134872
R74292 VINN.n387 VINN.n221 0.00134872
R74293 VINN.n407 VINN.n388 0.00134872
R74294 VINN.n385 VINN.n222 0.00134872
R74295 VINN.n408 VINN.n386 0.00134872
R74296 VINN.n383 VINN.n223 0.00134872
R74297 VINN.n409 VINN.n384 0.00134872
R74298 VINN.n381 VINN.n224 0.00134872
R74299 VINN.n410 VINN.n382 0.00134872
R74300 VINN.n379 VINN.n225 0.00134872
R74301 VINN.n411 VINN.n380 0.00134872
R74302 VINN.n377 VINN.n226 0.00134872
R74303 VINN.n412 VINN.n378 0.00134872
R74304 VINN.n375 VINN.n227 0.00134872
R74305 VINN.n413 VINN.n376 0.00134872
R74306 VINN.n373 VINN.n228 0.00134872
R74307 VINN.n414 VINN.n374 0.00134872
R74308 VINN.n371 VINN.n229 0.00134872
R74309 VINN.n415 VINN.n372 0.00134872
R74310 VINN.n369 VINN.n230 0.00134872
R74311 VINN.n416 VINN.n370 0.00134872
R74312 VINN.n367 VINN.n231 0.00134872
R74313 VINN.n417 VINN.n368 0.00134872
R74314 VINN.n365 VINN.n232 0.00134872
R74315 VINN.n418 VINN.n366 0.00134872
R74316 VINN.n363 VINN.n233 0.00134872
R74317 VINN.n419 VINN.n364 0.00134872
R74318 VINN.n361 VINN.n234 0.00134872
R74319 VINN.n420 VINN.n362 0.00134872
R74320 VINN.n359 VINN.n235 0.00134872
R74321 VINN.n421 VINN.n360 0.00134872
R74322 VINN.n357 VINN.n236 0.00134872
R74323 VINN.n422 VINN.n358 0.00134872
R74324 VINN.n355 VINN.n237 0.00134872
R74325 VINN.n423 VINN.n356 0.00134872
R74326 VINN.n353 VINN.n238 0.00134872
R74327 VINN.n424 VINN.n354 0.00134872
R74328 VINN.n351 VINN.n239 0.00134872
R74329 VINN.n425 VINN.n352 0.00134872
R74330 VINN.n349 VINN.n240 0.00134872
R74331 VINN.n426 VINN.n350 0.00134872
R74332 VINN.n347 VINN.n241 0.00134872
R74333 VINN.n427 VINN.n348 0.00134872
R74334 VINN.n345 VINN.n242 0.00134872
R74335 VINN.n428 VINN.n346 0.00134872
R74336 VINN.n343 VINN.n243 0.00134872
R74337 VINN.n429 VINN.n344 0.00134872
R74338 VINN.n341 VINN.n244 0.00134872
R74339 VINN.n430 VINN.n342 0.00134872
R74340 VINN.n339 VINN.n245 0.00134872
R74341 VINN.n431 VINN.n340 0.00134872
R74342 VINN.n337 VINN.n246 0.00134872
R74343 VINN.n432 VINN.n338 0.00134872
R74344 VINN.n335 VINN.n247 0.00134872
R74345 VINN.n433 VINN.n336 0.00134872
R74346 VINN.n333 VINN.n248 0.00134872
R74347 VINN.n434 VINN.n334 0.00134872
R74348 VINN.n331 VINN.n249 0.00134872
R74349 VINN.n435 VINN.n332 0.00134872
R74350 VINN.n329 VINN.n250 0.00134872
R74351 VINN.n436 VINN.n330 0.00134872
R74352 VINN.n327 VINN.n251 0.00134872
R74353 VINN.n437 VINN.n328 0.00134872
R74354 VINN.n325 VINN.n252 0.00134872
R74355 VINN.n438 VINN.n326 0.00134872
R74356 VINN.n323 VINN.n253 0.00134872
R74357 VINN.n439 VINN.n324 0.00134872
R74358 VINN.n321 VINN.n254 0.00134872
R74359 VINN.n440 VINN.n322 0.00134872
R74360 VINN.n319 VINN.n255 0.00134872
R74361 VINN.n441 VINN.n320 0.00134872
R74362 VINN.n317 VINN.n256 0.00134872
R74363 VINN.n442 VINN.n318 0.00134872
R74364 VINN.n315 VINN.n257 0.00134872
R74365 VINN.n443 VINN.n316 0.00134872
R74366 VINN.n313 VINN.n258 0.00134872
R74367 VINN.n444 VINN.n314 0.00134872
R74368 VINN.n311 VINN.n259 0.00134872
R74369 VINN.n445 VINN.n312 0.00134872
R74370 VINN.n309 VINN.n260 0.00134872
R74371 VINN.n446 VINN.n310 0.00134872
R74372 VINN.n307 VINN.n261 0.00134872
R74373 VINN.n447 VINN.n308 0.00134872
R74374 VINN.n305 VINN.n262 0.00134872
R74375 VINN.n448 VINN.n306 0.00134872
R74376 VINN.n303 VINN.n263 0.00134872
R74377 VINN.n449 VINN.n304 0.00134872
R74378 VINN.n301 VINN.n264 0.00134872
R74379 VINN.n450 VINN.n302 0.00134872
R74380 VINN.n299 VINN.n265 0.00134872
R74381 VINN.n451 VINN.n300 0.00134872
R74382 VINN.n297 VINN.n266 0.00134872
R74383 VINN.n452 VINN.n298 0.00134872
R74384 VINN.n295 VINN.n267 0.00134872
R74385 VINN.n453 VINN.n296 0.00134872
R74386 VINN.n293 VINN.n268 0.00134872
R74387 VINN.n454 VINN.n294 0.00134872
R74388 VINN.n291 VINN.n269 0.00134872
R74389 VINN.n455 VINN.n292 0.00134872
R74390 VINN.n289 VINN.n270 0.00134872
R74391 VINN.n456 VINN.n290 0.00134872
R74392 VINN.n287 VINN.n271 0.00134872
R74393 VINN.n457 VINN.n288 0.00134872
R74394 VINN.n285 VINN.n272 0.00134872
R74395 VINN.n458 VINN.n286 0.00134872
R74396 VINN.n283 VINN.n273 0.00134872
R74397 VINN.n459 VINN.n284 0.00134872
R74398 VINN.n281 VINN.n274 0.00134872
R74399 VINN.n460 VINN.n282 0.00134872
R74400 VINN.n279 VINN.n275 0.00134872
R74401 VINN.n461 VINN.n280 0.00134872
R74402 VINN.n277 VINN.n276 0.00134872
R74403 VINN.n461 VINN.n276 0.00134872
R74404 VINN.n460 VINN.n275 0.00134872
R74405 VINN.n459 VINN.n274 0.00134872
R74406 VINN.n458 VINN.n273 0.00134872
R74407 VINN.n457 VINN.n272 0.00134872
R74408 VINN.n456 VINN.n271 0.00134872
R74409 VINN.n455 VINN.n270 0.00134872
R74410 VINN.n454 VINN.n269 0.00134872
R74411 VINN.n453 VINN.n268 0.00134872
R74412 VINN.n452 VINN.n267 0.00134872
R74413 VINN.n451 VINN.n266 0.00134872
R74414 VINN.n450 VINN.n265 0.00134872
R74415 VINN.n449 VINN.n264 0.00134872
R74416 VINN.n448 VINN.n263 0.00134872
R74417 VINN.n447 VINN.n262 0.00134872
R74418 VINN.n446 VINN.n261 0.00134872
R74419 VINN.n445 VINN.n260 0.00134872
R74420 VINN.n444 VINN.n259 0.00134872
R74421 VINN.n443 VINN.n258 0.00134872
R74422 VINN.n442 VINN.n257 0.00134872
R74423 VINN.n441 VINN.n256 0.00134872
R74424 VINN.n440 VINN.n255 0.00134872
R74425 VINN.n439 VINN.n254 0.00134872
R74426 VINN.n438 VINN.n253 0.00134872
R74427 VINN.n437 VINN.n252 0.00134872
R74428 VINN.n436 VINN.n251 0.00134872
R74429 VINN.n435 VINN.n250 0.00134872
R74430 VINN.n434 VINN.n249 0.00134872
R74431 VINN.n433 VINN.n248 0.00134872
R74432 VINN.n432 VINN.n247 0.00134872
R74433 VINN.n431 VINN.n246 0.00134872
R74434 VINN.n430 VINN.n245 0.00134872
R74435 VINN.n429 VINN.n244 0.00134872
R74436 VINN.n428 VINN.n243 0.00134872
R74437 VINN.n427 VINN.n242 0.00134872
R74438 VINN.n426 VINN.n241 0.00134872
R74439 VINN.n425 VINN.n240 0.00134872
R74440 VINN.n424 VINN.n239 0.00134872
R74441 VINN.n423 VINN.n238 0.00134872
R74442 VINN.n422 VINN.n237 0.00134872
R74443 VINN.n421 VINN.n236 0.00134872
R74444 VINN.n420 VINN.n235 0.00134872
R74445 VINN.n419 VINN.n234 0.00134872
R74446 VINN.n418 VINN.n233 0.00134872
R74447 VINN.n417 VINN.n232 0.00134872
R74448 VINN.n416 VINN.n231 0.00134872
R74449 VINN.n415 VINN.n230 0.00134872
R74450 VINN.n414 VINN.n229 0.00134872
R74451 VINN.n413 VINN.n228 0.00134872
R74452 VINN.n412 VINN.n227 0.00134872
R74453 VINN.n411 VINN.n226 0.00134872
R74454 VINN.n410 VINN.n225 0.00134872
R74455 VINN.n409 VINN.n224 0.00134872
R74456 VINN.n408 VINN.n223 0.00134872
R74457 VINN.n407 VINN.n222 0.00134872
R74458 VINN.n406 VINN.n221 0.00134872
R74459 VINN.n405 VINN.n220 0.00134872
R74460 VINN.n404 VINN.n219 0.00134872
R74461 VINN.n403 VINN.n218 0.00134872
R74462 VINN.n402 VINN.n217 0.00134872
R74463 VINN.n401 VINN.n216 0.00134872
R74464 VINN.n464 VINN.n215 0.00134872
R74465 VINN.n528 VINN.n150 0.00134872
R74466 VINN.n657 VINN.n66 0.00134872
R74467 VINN.n462 VINN.n151 0.00134872
R74468 VINN.n280 VINN.n279 0.00134872
R74469 VINN.n282 VINN.n281 0.00134872
R74470 VINN.n284 VINN.n283 0.00134872
R74471 VINN.n286 VINN.n285 0.00134872
R74472 VINN.n288 VINN.n287 0.00134872
R74473 VINN.n290 VINN.n289 0.00134872
R74474 VINN.n292 VINN.n291 0.00134872
R74475 VINN.n294 VINN.n293 0.00134872
R74476 VINN.n296 VINN.n295 0.00134872
R74477 VINN.n298 VINN.n297 0.00134872
R74478 VINN.n300 VINN.n299 0.00134872
R74479 VINN.n302 VINN.n301 0.00134872
R74480 VINN.n304 VINN.n303 0.00134872
R74481 VINN.n306 VINN.n305 0.00134872
R74482 VINN.n308 VINN.n307 0.00134872
R74483 VINN.n310 VINN.n309 0.00134872
R74484 VINN.n312 VINN.n311 0.00134872
R74485 VINN.n314 VINN.n313 0.00134872
R74486 VINN.n316 VINN.n315 0.00134872
R74487 VINN.n318 VINN.n317 0.00134872
R74488 VINN.n320 VINN.n319 0.00134872
R74489 VINN.n322 VINN.n321 0.00134872
R74490 VINN.n324 VINN.n323 0.00134872
R74491 VINN.n326 VINN.n325 0.00134872
R74492 VINN.n328 VINN.n327 0.00134872
R74493 VINN.n330 VINN.n329 0.00134872
R74494 VINN.n332 VINN.n331 0.00134872
R74495 VINN.n334 VINN.n333 0.00134872
R74496 VINN.n336 VINN.n335 0.00134872
R74497 VINN.n338 VINN.n337 0.00134872
R74498 VINN.n340 VINN.n339 0.00134872
R74499 VINN.n342 VINN.n341 0.00134872
R74500 VINN.n344 VINN.n343 0.00134872
R74501 VINN.n346 VINN.n345 0.00134872
R74502 VINN.n348 VINN.n347 0.00134872
R74503 VINN.n350 VINN.n349 0.00134872
R74504 VINN.n352 VINN.n351 0.00134872
R74505 VINN.n354 VINN.n353 0.00134872
R74506 VINN.n356 VINN.n355 0.00134872
R74507 VINN.n358 VINN.n357 0.00134872
R74508 VINN.n360 VINN.n359 0.00134872
R74509 VINN.n362 VINN.n361 0.00134872
R74510 VINN.n364 VINN.n363 0.00134872
R74511 VINN.n366 VINN.n365 0.00134872
R74512 VINN.n368 VINN.n367 0.00134872
R74513 VINN.n370 VINN.n369 0.00134872
R74514 VINN.n372 VINN.n371 0.00134872
R74515 VINN.n374 VINN.n373 0.00134872
R74516 VINN.n376 VINN.n375 0.00134872
R74517 VINN.n378 VINN.n377 0.00134872
R74518 VINN.n380 VINN.n379 0.00134872
R74519 VINN.n382 VINN.n381 0.00134872
R74520 VINN.n384 VINN.n383 0.00134872
R74521 VINN.n386 VINN.n385 0.00134872
R74522 VINN.n388 VINN.n387 0.00134872
R74523 VINN.n390 VINN.n389 0.00134872
R74524 VINN.n392 VINN.n391 0.00134872
R74525 VINN.n394 VINN.n393 0.00134872
R74526 VINN.n396 VINN.n395 0.00134872
R74527 VINN.n398 VINN.n397 0.00134872
R74528 VINN.n400 VINN.n399 0.00134872
R74529 VINN.n654 VINN.n465 0.00134872
R74530 VINN.n151 VINN.n65 0.00134872
R74531 VINN.n278 VINN.n277 0.00134872
R74532 VINN.n466 VINN.n149 0.00134872
R74533 VINN.n152 VINN.n64 0.00134872
R74534 VINN.n467 VINN.n148 0.00134872
R74535 VINN.n153 VINN.n63 0.00134872
R74536 VINN.n468 VINN.n147 0.00134872
R74537 VINN.n154 VINN.n62 0.00134872
R74538 VINN.n469 VINN.n146 0.00134872
R74539 VINN.n155 VINN.n61 0.00134872
R74540 VINN.n470 VINN.n145 0.00134872
R74541 VINN.n156 VINN.n60 0.00134872
R74542 VINN.n471 VINN.n144 0.00134872
R74543 VINN.n157 VINN.n59 0.00134872
R74544 VINN.n472 VINN.n143 0.00134872
R74545 VINN.n158 VINN.n58 0.00134872
R74546 VINN.n473 VINN.n142 0.00134872
R74547 VINN.n159 VINN.n57 0.00134872
R74548 VINN.n474 VINN.n141 0.00134872
R74549 VINN.n160 VINN.n56 0.00134872
R74550 VINN.n475 VINN.n140 0.00134872
R74551 VINN.n161 VINN.n55 0.00134872
R74552 VINN.n476 VINN.n139 0.00134872
R74553 VINN.n162 VINN.n54 0.00134872
R74554 VINN.n477 VINN.n138 0.00134872
R74555 VINN.n163 VINN.n53 0.00134872
R74556 VINN.n478 VINN.n137 0.00134872
R74557 VINN.n164 VINN.n52 0.00134872
R74558 VINN.n479 VINN.n136 0.00134872
R74559 VINN.n165 VINN.n51 0.00134872
R74560 VINN.n480 VINN.n135 0.00134872
R74561 VINN.n166 VINN.n50 0.00134872
R74562 VINN.n481 VINN.n134 0.00134872
R74563 VINN.n167 VINN.n49 0.00134872
R74564 VINN.n482 VINN.n133 0.00134872
R74565 VINN.n168 VINN.n48 0.00134872
R74566 VINN.n483 VINN.n132 0.00134872
R74567 VINN.n169 VINN.n47 0.00134872
R74568 VINN.n484 VINN.n131 0.00134872
R74569 VINN.n170 VINN.n46 0.00134872
R74570 VINN.n485 VINN.n130 0.00134872
R74571 VINN.n171 VINN.n45 0.00134872
R74572 VINN.n486 VINN.n129 0.00134872
R74573 VINN.n172 VINN.n44 0.00134872
R74574 VINN.n487 VINN.n128 0.00134872
R74575 VINN.n173 VINN.n43 0.00134872
R74576 VINN.n488 VINN.n127 0.00134872
R74577 VINN.n174 VINN.n42 0.00134872
R74578 VINN.n489 VINN.n126 0.00134872
R74579 VINN.n175 VINN.n41 0.00134872
R74580 VINN.n490 VINN.n125 0.00134872
R74581 VINN.n176 VINN.n40 0.00134872
R74582 VINN.n491 VINN.n124 0.00134872
R74583 VINN.n177 VINN.n39 0.00134872
R74584 VINN.n492 VINN.n123 0.00134872
R74585 VINN.n178 VINN.n38 0.00134872
R74586 VINN.n493 VINN.n122 0.00134872
R74587 VINN.n179 VINN.n37 0.00134872
R74588 VINN.n494 VINN.n121 0.00134872
R74589 VINN.n180 VINN.n36 0.00134872
R74590 VINN.n495 VINN.n120 0.00134872
R74591 VINN.n181 VINN.n35 0.00134872
R74592 VINN.n496 VINN.n119 0.00134872
R74593 VINN.n182 VINN.n34 0.00134872
R74594 VINN.n497 VINN.n118 0.00134872
R74595 VINN.n183 VINN.n33 0.00134872
R74596 VINN.n498 VINN.n117 0.00134872
R74597 VINN.n184 VINN.n32 0.00134872
R74598 VINN.n499 VINN.n116 0.00134872
R74599 VINN.n185 VINN.n31 0.00134872
R74600 VINN.n500 VINN.n115 0.00134872
R74601 VINN.n186 VINN.n30 0.00134872
R74602 VINN.n501 VINN.n114 0.00134872
R74603 VINN.n187 VINN.n29 0.00134872
R74604 VINN.n502 VINN.n113 0.00134872
R74605 VINN.n188 VINN.n28 0.00134872
R74606 VINN.n503 VINN.n112 0.00134872
R74607 VINN.n189 VINN.n27 0.00134872
R74608 VINN.n504 VINN.n111 0.00134872
R74609 VINN.n190 VINN.n26 0.00134872
R74610 VINN.n505 VINN.n110 0.00134872
R74611 VINN.n191 VINN.n25 0.00134872
R74612 VINN.n506 VINN.n109 0.00134872
R74613 VINN.n192 VINN.n24 0.00134872
R74614 VINN.n507 VINN.n108 0.00134872
R74615 VINN.n193 VINN.n23 0.00134872
R74616 VINN.n508 VINN.n107 0.00134872
R74617 VINN.n194 VINN.n22 0.00134872
R74618 VINN.n509 VINN.n106 0.00134872
R74619 VINN.n195 VINN.n21 0.00134872
R74620 VINN.n510 VINN.n105 0.00134872
R74621 VINN.n196 VINN.n20 0.00134872
R74622 VINN.n511 VINN.n104 0.00134872
R74623 VINN.n197 VINN.n19 0.00134872
R74624 VINN.n512 VINN.n103 0.00134872
R74625 VINN.n198 VINN.n18 0.00134872
R74626 VINN.n513 VINN.n102 0.00134872
R74627 VINN.n199 VINN.n17 0.00134872
R74628 VINN.n514 VINN.n101 0.00134872
R74629 VINN.n200 VINN.n16 0.00134872
R74630 VINN.n515 VINN.n100 0.00134872
R74631 VINN.n201 VINN.n15 0.00134872
R74632 VINN.n516 VINN.n99 0.00134872
R74633 VINN.n202 VINN.n14 0.00134872
R74634 VINN.n517 VINN.n98 0.00134872
R74635 VINN.n203 VINN.n13 0.00134872
R74636 VINN.n518 VINN.n97 0.00134872
R74637 VINN.n204 VINN.n12 0.00134872
R74638 VINN.n519 VINN.n96 0.00134872
R74639 VINN.n205 VINN.n11 0.00134872
R74640 VINN.n520 VINN.n95 0.00134872
R74641 VINN.n206 VINN.n10 0.00134872
R74642 VINN.n521 VINN.n94 0.00134872
R74643 VINN.n207 VINN.n9 0.00134872
R74644 VINN.n522 VINN.n93 0.00134872
R74645 VINN.n208 VINN.n8 0.00134872
R74646 VINN.n523 VINN.n92 0.00134872
R74647 VINN.n209 VINN.n7 0.00134872
R74648 VINN.n524 VINN.n91 0.00134872
R74649 VINN.n210 VINN.n6 0.00134872
R74650 VINN.n525 VINN.n90 0.00134872
R74651 VINN.n211 VINN.n5 0.00134872
R74652 VINN.n526 VINN.n89 0.00134872
R74653 VINN.n212 VINN.n4 0.00134872
R74654 VINN.n527 VINN.n88 0.00134872
R74655 VINN.n213 VINN.n3 0.00134872
R74656 VINN.n214 VINN.n87 0.00134872
R74657 VINN.n655 VINN.n2 0.00134872
R74658 VINN.n657 VINN.n656 0.0011975
R74659 VINN.n658 VINN.n1 0.000965
R74660 VINN.n529 VINN.n1 0.000965
R74661 VINN.n653 VINN.n529 0.000965
R74662 VINN.n653 VINN.n652 0.000965
R74663 VINN.n652 VINN.n651 0.000965
R74664 VINN.n651 VINN.n650 0.000965
R74665 VINN.n650 VINN.n649 0.000965
R74666 VINN.n649 VINN.n648 0.000965
R74667 VINN.n648 VINN.n647 0.000965
R74668 VINN.n647 VINN.n646 0.000965
R74669 VINN.n646 VINN.n645 0.000965
R74670 VINN.n645 VINN.n644 0.000965
R74671 VINN.n644 VINN.n643 0.000965
R74672 VINN.n643 VINN.n642 0.000965
R74673 VINN.n642 VINN.n641 0.000965
R74674 VINN.n641 VINN.n640 0.000965
R74675 VINN.n640 VINN.n639 0.000965
R74676 VINN.n639 VINN.n638 0.000965
R74677 VINN.n638 VINN.n637 0.000965
R74678 VINN.n637 VINN.n636 0.000965
R74679 VINN.n636 VINN.n635 0.000965
R74680 VINN.n635 VINN.n634 0.000965
R74681 VINN.n634 VINN.n633 0.000965
R74682 VINN.n633 VINN.n632 0.000965
R74683 VINN.n632 VINN.n631 0.000965
R74684 VINN.n631 VINN.n630 0.000965
R74685 VINN.n630 VINN.n629 0.000965
R74686 VINN.n629 VINN.n628 0.000965
R74687 VINN.n628 VINN.n627 0.000965
R74688 VINN.n627 VINN.n626 0.000965
R74689 VINN.n626 VINN.n625 0.000965
R74690 VINN.n625 VINN.n624 0.000965
R74691 VINN.n624 VINN.n623 0.000965
R74692 VINN.n623 VINN.n622 0.000965
R74693 VINN.n622 VINN.n621 0.000965
R74694 VINN.n621 VINN.n620 0.000965
R74695 VINN.n620 VINN.n619 0.000965
R74696 VINN.n619 VINN.n618 0.000965
R74697 VINN.n618 VINN.n617 0.000965
R74698 VINN.n617 VINN.n616 0.000965
R74699 VINN.n616 VINN.n615 0.000965
R74700 VINN.n615 VINN.n614 0.000965
R74701 VINN.n614 VINN.n613 0.000965
R74702 VINN.n613 VINN.n612 0.000965
R74703 VINN.n612 VINN.n611 0.000965
R74704 VINN.n611 VINN.n610 0.000965
R74705 VINN.n610 VINN.n609 0.000965
R74706 VINN.n609 VINN.n608 0.000965
R74707 VINN.n608 VINN.n607 0.000965
R74708 VINN.n607 VINN.n606 0.000965
R74709 VINN.n606 VINN.n605 0.000965
R74710 VINN.n605 VINN.n604 0.000965
R74711 VINN.n604 VINN.n603 0.000965
R74712 VINN.n603 VINN.n602 0.000965
R74713 VINN.n602 VINN.n601 0.000965
R74714 VINN.n601 VINN.n600 0.000965
R74715 VINN.n600 VINN.n599 0.000965
R74716 VINN.n599 VINN.n598 0.000965
R74717 VINN.n598 VINN.n597 0.000965
R74718 VINN.n597 VINN.n596 0.000965
R74719 VINN.n596 VINN.n595 0.000965
R74720 VINN.n595 VINN.n594 0.000965
R74721 VINN.n594 VINN.n593 0.000965
R74722 VINN.n593 VINN.n592 0.000965
R74723 VINN.n592 VINN.n591 0.000965
R74724 VINN.n591 VINN.n590 0.000965
R74725 VINN.n590 VINN.n589 0.000965
R74726 VINN.n589 VINN.n588 0.000965
R74727 VINN.n588 VINN.n587 0.000965
R74728 VINN.n587 VINN.n586 0.000965
R74729 VINN.n586 VINN.n585 0.000965
R74730 VINN.n585 VINN.n584 0.000965
R74731 VINN.n584 VINN.n583 0.000965
R74732 VINN.n583 VINN.n582 0.000965
R74733 VINN.n582 VINN.n581 0.000965
R74734 VINN.n581 VINN.n580 0.000965
R74735 VINN.n580 VINN.n579 0.000965
R74736 VINN.n579 VINN.n578 0.000965
R74737 VINN.n578 VINN.n577 0.000965
R74738 VINN.n577 VINN.n576 0.000965
R74739 VINN.n576 VINN.n575 0.000965
R74740 VINN.n574 VINN.n573 0.000965
R74741 VINN.n573 VINN.n572 0.000965
R74742 VINN.n572 VINN.n571 0.000965
R74743 VINN.n571 VINN.n570 0.000965
R74744 VINN.n570 VINN.n569 0.000965
R74745 VINN.n569 VINN.n568 0.000965
R74746 VINN.n568 VINN.n567 0.000965
R74747 VINN.n567 VINN.n566 0.000965
R74748 VINN.n566 VINN.n565 0.000965
R74749 VINN.n565 VINN.n564 0.000965
R74750 VINN.n564 VINN.n563 0.000965
R74751 VINN.n563 VINN.n562 0.000965
R74752 VINN.n562 VINN.n561 0.000965
R74753 VINN.n561 VINN.n560 0.000965
R74754 VINN.n560 VINN.n559 0.000965
R74755 VINN.n559 VINN.n558 0.000965
R74756 VINN.n558 VINN.n557 0.000965
R74757 VINN.n557 VINN.n556 0.000965
R74758 VINN.n556 VINN.n555 0.000965
R74759 VINN.n555 VINN.n554 0.000965
R74760 VINN.n554 VINN.n553 0.000965
R74761 VINN.n553 VINN.n552 0.000965
R74762 VINN.n552 VINN.n551 0.000965
R74763 VINN.n551 VINN.n550 0.000965
R74764 VINN.n550 VINN.n549 0.000965
R74765 VINN.n549 VINN.n548 0.000965
R74766 VINN.n548 VINN.n547 0.000965
R74767 VINN.n547 VINN.n546 0.000965
R74768 VINN.n546 VINN.n545 0.000965
R74769 VINN.n545 VINN.n544 0.000965
R74770 VINN.n544 VINN.n543 0.000965
R74771 VINN.n543 VINN.n542 0.000965
R74772 VINN.n542 VINN.n541 0.000965
R74773 VINN.n541 VINN.n540 0.000965
R74774 VINN.n540 VINN.n539 0.000965
R74775 VINN.n539 VINN.n538 0.000965
R74776 VINN.n538 VINN.n537 0.000965
R74777 VINN.n537 VINN.n536 0.000965
R74778 VINN.n536 VINN.n535 0.000965
R74779 VINN.n535 VINN.n534 0.000965
R74780 VINN.n534 VINN.n533 0.000965
R74781 VINN.n533 VINN.n532 0.000965
R74782 VINN.n532 VINN.n531 0.000965
R74783 VINN.n531 VINN.n530 0.000965
R74784 VINN.n575 VINN 0.00089
R74785 VINN VINN.n574 0.000575
R74786 a_2044_n43060.n0 a_2044_n43060.t22 47.2735
R74787 a_2044_n43060.n0 a_2044_n43060.t0 45.5905
R74788 a_2044_n43060.n13 a_2044_n43060.t5 9.50526
R74789 a_2044_n43060.n0 a_2044_n43060.t1 9.36137
R74790 a_2044_n43060.n1 a_2044_n43060.t4 9.32226
R74791 a_2044_n43060.n13 a_2044_n43060.n12 7.97226
R74792 a_2044_n43060.n15 a_2044_n43060.n14 7.97226
R74793 a_2044_n43060.n17 a_2044_n43060.n16 7.97226
R74794 a_2044_n43060.n11 a_2044_n43060.n10 7.97226
R74795 a_2044_n43060.n9 a_2044_n43060.n8 7.97226
R74796 a_2044_n43060.n7 a_2044_n43060.n6 7.97226
R74797 a_2044_n43060.n5 a_2044_n43060.n4 7.97226
R74798 a_2044_n43060.n3 a_2044_n43060.n2 7.97226
R74799 a_2044_n43060.n19 a_2044_n43060.n18 7.97226
R74800 a_2044_n43060.n1 a_2044_n43060.n0 1.31354
R74801 a_2044_n43060.n12 a_2044_n43060.t17 0.6505
R74802 a_2044_n43060.n12 a_2044_n43060.t13 0.6505
R74803 a_2044_n43060.n14 a_2044_n43060.t6 0.6505
R74804 a_2044_n43060.n14 a_2044_n43060.t9 0.6505
R74805 a_2044_n43060.n16 a_2044_n43060.t2 0.6505
R74806 a_2044_n43060.n16 a_2044_n43060.t18 0.6505
R74807 a_2044_n43060.n10 a_2044_n43060.t11 0.6505
R74808 a_2044_n43060.n10 a_2044_n43060.t19 0.6505
R74809 a_2044_n43060.n8 a_2044_n43060.t20 0.6505
R74810 a_2044_n43060.n8 a_2044_n43060.t15 0.6505
R74811 a_2044_n43060.n6 a_2044_n43060.t12 0.6505
R74812 a_2044_n43060.n6 a_2044_n43060.t7 0.6505
R74813 a_2044_n43060.n4 a_2044_n43060.t8 0.6505
R74814 a_2044_n43060.n4 a_2044_n43060.t3 0.6505
R74815 a_2044_n43060.n2 a_2044_n43060.t16 0.6505
R74816 a_2044_n43060.n2 a_2044_n43060.t14 0.6505
R74817 a_2044_n43060.t21 a_2044_n43060.n19 0.6505
R74818 a_2044_n43060.n19 a_2044_n43060.t10 0.6505
R74819 a_2044_n43060.n3 a_2044_n43060.n1 0.1835
R74820 a_2044_n43060.n5 a_2044_n43060.n3 0.1625
R74821 a_2044_n43060.n7 a_2044_n43060.n5 0.1625
R74822 a_2044_n43060.n9 a_2044_n43060.n7 0.1625
R74823 a_2044_n43060.n11 a_2044_n43060.n9 0.1625
R74824 a_2044_n43060.n18 a_2044_n43060.n11 0.1625
R74825 a_2044_n43060.n18 a_2044_n43060.n17 0.1625
R74826 a_2044_n43060.n17 a_2044_n43060.n15 0.1625
R74827 a_2044_n43060.n15 a_2044_n43060.n13 0.1625
R74828 IB.n0 IB.t9 50.7028
R74829 IB.n24 IB.t21 50.638
R74830 IB.n23 IB.t13 50.638
R74831 IB.n22 IB.t22 50.638
R74832 IB.n21 IB.t11 50.638
R74833 IB.n20 IB.t6 50.638
R74834 IB.n19 IB.t28 50.638
R74835 IB.n18 IB.t8 50.638
R74836 IB.n17 IB.t4 50.638
R74837 IB.n16 IB.t14 50.638
R74838 IB.n15 IB.t19 50.638
R74839 IB.n14 IB.t7 50.638
R74840 IB.n13 IB.t20 50.638
R74841 IB.n12 IB.t12 50.638
R74842 IB.n11 IB.t23 50.638
R74843 IB.n10 IB.t25 50.638
R74844 IB.n9 IB.t17 50.638
R74845 IB.n8 IB.t26 50.638
R74846 IB.n7 IB.t18 50.638
R74847 IB.n6 IB.t15 50.638
R74848 IB.n5 IB.t5 50.638
R74849 IB.n4 IB.t27 50.638
R74850 IB.n3 IB.t10 50.638
R74851 IB.n2 IB.t29 50.638
R74852 IB.n1 IB.t24 50.638
R74853 IB.n0 IB.t16 50.638
R74854 IB.n27 IB.t2 46.138
R74855 IB.n26 IB.t0 46.138
R74856 IB IB.n28 12.0813
R74857 IB.n27 IB.t3 9.37595
R74858 IB.n26 IB.t1 9.37595
R74859 IB.n26 IB.n25 4.5005
R74860 IB.n28 IB.n27 4.5005
R74861 IB.n19 IB.n18 0.6347
R74862 IB.n23 IB.n22 0.6347
R74863 IB.n25 IB.n24 0.6053
R74864 IB.n1 IB.n0 0.0653
R74865 IB.n2 IB.n1 0.0653
R74866 IB.n3 IB.n2 0.0653
R74867 IB.n4 IB.n3 0.0653
R74868 IB.n5 IB.n4 0.0653
R74869 IB.n6 IB.n5 0.0653
R74870 IB.n7 IB.n6 0.0653
R74871 IB.n8 IB.n7 0.0653
R74872 IB.n9 IB.n8 0.0653
R74873 IB.n10 IB.n9 0.0653
R74874 IB.n11 IB.n10 0.0653
R74875 IB.n12 IB.n11 0.0653
R74876 IB.n13 IB.n12 0.0653
R74877 IB.n14 IB.n13 0.0653
R74878 IB.n15 IB.n14 0.0653
R74879 IB.n16 IB.n15 0.0653
R74880 IB.n17 IB.n16 0.0653
R74881 IB.n18 IB.n17 0.0653
R74882 IB.n20 IB.n19 0.0653
R74883 IB.n21 IB.n20 0.0653
R74884 IB.n22 IB.n21 0.0653
R74885 IB.n24 IB.n23 0.0653
R74886 IB.n28 IB.n25 0.0653
R74887 IB.n27 IB.n26 0.0513901
R74888 VDD.n766 VDD.t42 270.493
R74889 VDD.t46 VDD.n764 270.493
R74890 VDD.n733 VDD.t2 270.493
R74891 VDD.t14 VDD.n731 270.493
R74892 VDD.t28 VDD.n403 270.493
R74893 VDD.t52 VDD.n405 270.493
R74894 VDD.n720 VDD.t30 270.493
R74895 VDD.t16 VDD.n718 270.493
R74896 VDD.n766 VDD.n669 235.089
R74897 VDD.n766 VDD.n670 235.089
R74898 VDD.n764 VDD.n669 235.089
R74899 VDD.n764 VDD.n670 235.089
R74900 VDD.t42 VDD.t26 169.28
R74901 VDD.t26 VDD.t10 169.28
R74902 VDD.t10 VDD.t0 169.28
R74903 VDD.t0 VDD.t40 169.28
R74904 VDD.t40 VDD.t4 169.28
R74905 VDD.t4 VDD.t50 169.28
R74906 VDD.t50 VDD.t32 169.28
R74907 VDD.t32 VDD.t22 169.28
R74908 VDD.t22 VDD.t6 169.28
R74909 VDD.t24 VDD.t8 169.28
R74910 VDD.t8 VDD.t12 169.28
R74911 VDD.t12 VDD.t36 169.28
R74912 VDD.t36 VDD.t18 169.28
R74913 VDD.t18 VDD.t48 169.28
R74914 VDD.t48 VDD.t20 169.28
R74915 VDD.t20 VDD.t34 169.28
R74916 VDD.t34 VDD.t54 169.28
R74917 VDD.t54 VDD.t46 169.28
R74918 VDD.t2 VDD.t44 169.28
R74919 VDD.t38 VDD.t14 169.28
R74920 VDD.n731 VDD.n673 91.8479
R74921 VDD.n731 VDD.n674 91.8479
R74922 VDD.n733 VDD.n674 91.8479
R74923 VDD.n733 VDD.n673 91.8479
R74924 VDD.t6 VDD.n765 84.64
R74925 VDD.n765 VDD.t24 84.64
R74926 VDD.t44 VDD.n732 84.64
R74927 VDD.n732 VDD.t38 84.64
R74928 VDD.n951 VDD.t28 84.64
R74929 VDD.n951 VDD.t52 84.64
R74930 VDD.t30 VDD.n719 84.64
R74931 VDD.n719 VDD.t16 84.64
R74932 VDD.n720 VDD.n692 73.9426
R74933 VDD.n718 VDD.n692 73.9426
R74934 VDD.n720 VDD.n694 73.9426
R74935 VDD.n718 VDD.n694 73.9426
R74936 VDD.n950 VDD.n405 73.9426
R74937 VDD.n952 VDD.n405 73.9426
R74938 VDD.n952 VDD.n403 73.9426
R74939 VDD.n950 VDD.n403 73.9426
R74940 VDD.n1607 VDD.n1341 4.5005
R74941 VDD.n1607 VDD.n1415 4.5005
R74942 VDD.n1674 VDD.n1607 4.5005
R74943 VDD.n1416 VDD.n1342 4.5005
R74944 VDD.n1416 VDD.n1340 4.5005
R74945 VDD.n1416 VDD.n1344 4.5005
R74946 VDD.n1416 VDD.n1339 4.5005
R74947 VDD.n1416 VDD.n1345 4.5005
R74948 VDD.n1416 VDD.n1338 4.5005
R74949 VDD.n1416 VDD.n1347 4.5005
R74950 VDD.n1416 VDD.n1337 4.5005
R74951 VDD.n1416 VDD.n1348 4.5005
R74952 VDD.n1416 VDD.n1336 4.5005
R74953 VDD.n1416 VDD.n1350 4.5005
R74954 VDD.n1416 VDD.n1335 4.5005
R74955 VDD.n1416 VDD.n1351 4.5005
R74956 VDD.n1416 VDD.n1334 4.5005
R74957 VDD.n1416 VDD.n1353 4.5005
R74958 VDD.n1416 VDD.n1333 4.5005
R74959 VDD.n1416 VDD.n1354 4.5005
R74960 VDD.n1416 VDD.n1332 4.5005
R74961 VDD.n1416 VDD.n1356 4.5005
R74962 VDD.n1416 VDD.n1331 4.5005
R74963 VDD.n1416 VDD.n1357 4.5005
R74964 VDD.n1416 VDD.n1330 4.5005
R74965 VDD.n1416 VDD.n1359 4.5005
R74966 VDD.n1416 VDD.n1329 4.5005
R74967 VDD.n1416 VDD.n1360 4.5005
R74968 VDD.n1416 VDD.n1328 4.5005
R74969 VDD.n1416 VDD.n1362 4.5005
R74970 VDD.n1416 VDD.n1327 4.5005
R74971 VDD.n1416 VDD.n1363 4.5005
R74972 VDD.n1416 VDD.n1326 4.5005
R74973 VDD.n1416 VDD.n1365 4.5005
R74974 VDD.n1416 VDD.n1325 4.5005
R74975 VDD.n1416 VDD.n1366 4.5005
R74976 VDD.n1416 VDD.n1324 4.5005
R74977 VDD.n1416 VDD.n1368 4.5005
R74978 VDD.n1416 VDD.n1323 4.5005
R74979 VDD.n1416 VDD.n1369 4.5005
R74980 VDD.n1416 VDD.n1322 4.5005
R74981 VDD.n1416 VDD.n1371 4.5005
R74982 VDD.n1416 VDD.n1321 4.5005
R74983 VDD.n1416 VDD.n1372 4.5005
R74984 VDD.n1416 VDD.n1320 4.5005
R74985 VDD.n1416 VDD.n1374 4.5005
R74986 VDD.n1416 VDD.n1319 4.5005
R74987 VDD.n1416 VDD.n1375 4.5005
R74988 VDD.n1416 VDD.n1318 4.5005
R74989 VDD.n1416 VDD.n1376 4.5005
R74990 VDD.n1416 VDD.n1316 4.5005
R74991 VDD.n1416 VDD.n1377 4.5005
R74992 VDD.n1416 VDD.n1315 4.5005
R74993 VDD.n1416 VDD.n1378 4.5005
R74994 VDD.n1416 VDD.n1313 4.5005
R74995 VDD.n1416 VDD.n1379 4.5005
R74996 VDD.n1416 VDD.n1312 4.5005
R74997 VDD.n1416 VDD.n1380 4.5005
R74998 VDD.n1416 VDD.n1310 4.5005
R74999 VDD.n1416 VDD.n1381 4.5005
R75000 VDD.n1416 VDD.n1309 4.5005
R75001 VDD.n1416 VDD.n1382 4.5005
R75002 VDD.n1416 VDD.n1307 4.5005
R75003 VDD.n1416 VDD.n1383 4.5005
R75004 VDD.n1416 VDD.n1306 4.5005
R75005 VDD.n1416 VDD.n1384 4.5005
R75006 VDD.n1416 VDD.n1304 4.5005
R75007 VDD.n1416 VDD.n1385 4.5005
R75008 VDD.n1416 VDD.n1303 4.5005
R75009 VDD.n1416 VDD.n1386 4.5005
R75010 VDD.n1416 VDD.n1301 4.5005
R75011 VDD.n1416 VDD.n1387 4.5005
R75012 VDD.n1416 VDD.n1300 4.5005
R75013 VDD.n1416 VDD.n1388 4.5005
R75014 VDD.n1416 VDD.n1298 4.5005
R75015 VDD.n1416 VDD.n1389 4.5005
R75016 VDD.n1416 VDD.n1297 4.5005
R75017 VDD.n1416 VDD.n1390 4.5005
R75018 VDD.n1416 VDD.n1295 4.5005
R75019 VDD.n1416 VDD.n1391 4.5005
R75020 VDD.n1416 VDD.n1294 4.5005
R75021 VDD.n1416 VDD.n1392 4.5005
R75022 VDD.n1416 VDD.n1292 4.5005
R75023 VDD.n1416 VDD.n1393 4.5005
R75024 VDD.n1416 VDD.n1291 4.5005
R75025 VDD.n1416 VDD.n1394 4.5005
R75026 VDD.n1416 VDD.n1289 4.5005
R75027 VDD.n1416 VDD.n1395 4.5005
R75028 VDD.n1416 VDD.n1288 4.5005
R75029 VDD.n1416 VDD.n1396 4.5005
R75030 VDD.n1416 VDD.n1286 4.5005
R75031 VDD.n1416 VDD.n1397 4.5005
R75032 VDD.n1416 VDD.n1285 4.5005
R75033 VDD.n1416 VDD.n1398 4.5005
R75034 VDD.n1416 VDD.n1283 4.5005
R75035 VDD.n1416 VDD.n1399 4.5005
R75036 VDD.n1416 VDD.n1282 4.5005
R75037 VDD.n1416 VDD.n1400 4.5005
R75038 VDD.n1416 VDD.n1280 4.5005
R75039 VDD.n1416 VDD.n1401 4.5005
R75040 VDD.n1416 VDD.n1279 4.5005
R75041 VDD.n1416 VDD.n1402 4.5005
R75042 VDD.n1416 VDD.n1277 4.5005
R75043 VDD.n1416 VDD.n1403 4.5005
R75044 VDD.n1416 VDD.n1276 4.5005
R75045 VDD.n1416 VDD.n1404 4.5005
R75046 VDD.n1416 VDD.n1274 4.5005
R75047 VDD.n1416 VDD.n1405 4.5005
R75048 VDD.n1416 VDD.n1273 4.5005
R75049 VDD.n1416 VDD.n1406 4.5005
R75050 VDD.n1416 VDD.n1271 4.5005
R75051 VDD.n1416 VDD.n1407 4.5005
R75052 VDD.n1416 VDD.n1270 4.5005
R75053 VDD.n1416 VDD.n1408 4.5005
R75054 VDD.n1416 VDD.n1268 4.5005
R75055 VDD.n1416 VDD.n1409 4.5005
R75056 VDD.n1416 VDD.n1267 4.5005
R75057 VDD.n1416 VDD.n1410 4.5005
R75058 VDD.n1416 VDD.n1265 4.5005
R75059 VDD.n1416 VDD.n1411 4.5005
R75060 VDD.n1416 VDD.n1264 4.5005
R75061 VDD.n1416 VDD.n1412 4.5005
R75062 VDD.n1416 VDD.n1262 4.5005
R75063 VDD.n1416 VDD.n1413 4.5005
R75064 VDD.n1416 VDD.n1261 4.5005
R75065 VDD.n1416 VDD.n1414 4.5005
R75066 VDD.n1416 VDD.n1415 4.5005
R75067 VDD.n1674 VDD.n1416 4.5005
R75068 VDD.n1676 VDD.n1196 4.5005
R75069 VDD.n1341 VDD.n1196 4.5005
R75070 VDD.n1342 VDD.n1196 4.5005
R75071 VDD.n1340 VDD.n1196 4.5005
R75072 VDD.n1344 VDD.n1196 4.5005
R75073 VDD.n1339 VDD.n1196 4.5005
R75074 VDD.n1345 VDD.n1196 4.5005
R75075 VDD.n1338 VDD.n1196 4.5005
R75076 VDD.n1347 VDD.n1196 4.5005
R75077 VDD.n1337 VDD.n1196 4.5005
R75078 VDD.n1348 VDD.n1196 4.5005
R75079 VDD.n1336 VDD.n1196 4.5005
R75080 VDD.n1350 VDD.n1196 4.5005
R75081 VDD.n1335 VDD.n1196 4.5005
R75082 VDD.n1351 VDD.n1196 4.5005
R75083 VDD.n1334 VDD.n1196 4.5005
R75084 VDD.n1353 VDD.n1196 4.5005
R75085 VDD.n1333 VDD.n1196 4.5005
R75086 VDD.n1354 VDD.n1196 4.5005
R75087 VDD.n1332 VDD.n1196 4.5005
R75088 VDD.n1356 VDD.n1196 4.5005
R75089 VDD.n1331 VDD.n1196 4.5005
R75090 VDD.n1357 VDD.n1196 4.5005
R75091 VDD.n1330 VDD.n1196 4.5005
R75092 VDD.n1359 VDD.n1196 4.5005
R75093 VDD.n1329 VDD.n1196 4.5005
R75094 VDD.n1360 VDD.n1196 4.5005
R75095 VDD.n1328 VDD.n1196 4.5005
R75096 VDD.n1362 VDD.n1196 4.5005
R75097 VDD.n1327 VDD.n1196 4.5005
R75098 VDD.n1363 VDD.n1196 4.5005
R75099 VDD.n1326 VDD.n1196 4.5005
R75100 VDD.n1365 VDD.n1196 4.5005
R75101 VDD.n1325 VDD.n1196 4.5005
R75102 VDD.n1366 VDD.n1196 4.5005
R75103 VDD.n1324 VDD.n1196 4.5005
R75104 VDD.n1368 VDD.n1196 4.5005
R75105 VDD.n1323 VDD.n1196 4.5005
R75106 VDD.n1369 VDD.n1196 4.5005
R75107 VDD.n1322 VDD.n1196 4.5005
R75108 VDD.n1371 VDD.n1196 4.5005
R75109 VDD.n1321 VDD.n1196 4.5005
R75110 VDD.n1372 VDD.n1196 4.5005
R75111 VDD.n1320 VDD.n1196 4.5005
R75112 VDD.n1374 VDD.n1196 4.5005
R75113 VDD.n1319 VDD.n1196 4.5005
R75114 VDD.n1375 VDD.n1196 4.5005
R75115 VDD.n1318 VDD.n1196 4.5005
R75116 VDD.n1376 VDD.n1196 4.5005
R75117 VDD.n1316 VDD.n1196 4.5005
R75118 VDD.n1377 VDD.n1196 4.5005
R75119 VDD.n1315 VDD.n1196 4.5005
R75120 VDD.n1378 VDD.n1196 4.5005
R75121 VDD.n1313 VDD.n1196 4.5005
R75122 VDD.n1379 VDD.n1196 4.5005
R75123 VDD.n1312 VDD.n1196 4.5005
R75124 VDD.n1380 VDD.n1196 4.5005
R75125 VDD.n1310 VDD.n1196 4.5005
R75126 VDD.n1381 VDD.n1196 4.5005
R75127 VDD.n1309 VDD.n1196 4.5005
R75128 VDD.n1382 VDD.n1196 4.5005
R75129 VDD.n1307 VDD.n1196 4.5005
R75130 VDD.n1383 VDD.n1196 4.5005
R75131 VDD.n1306 VDD.n1196 4.5005
R75132 VDD.n1384 VDD.n1196 4.5005
R75133 VDD.n1304 VDD.n1196 4.5005
R75134 VDD.n1385 VDD.n1196 4.5005
R75135 VDD.n1303 VDD.n1196 4.5005
R75136 VDD.n1386 VDD.n1196 4.5005
R75137 VDD.n1301 VDD.n1196 4.5005
R75138 VDD.n1387 VDD.n1196 4.5005
R75139 VDD.n1300 VDD.n1196 4.5005
R75140 VDD.n1388 VDD.n1196 4.5005
R75141 VDD.n1298 VDD.n1196 4.5005
R75142 VDD.n1389 VDD.n1196 4.5005
R75143 VDD.n1297 VDD.n1196 4.5005
R75144 VDD.n1390 VDD.n1196 4.5005
R75145 VDD.n1295 VDD.n1196 4.5005
R75146 VDD.n1391 VDD.n1196 4.5005
R75147 VDD.n1294 VDD.n1196 4.5005
R75148 VDD.n1392 VDD.n1196 4.5005
R75149 VDD.n1292 VDD.n1196 4.5005
R75150 VDD.n1393 VDD.n1196 4.5005
R75151 VDD.n1291 VDD.n1196 4.5005
R75152 VDD.n1394 VDD.n1196 4.5005
R75153 VDD.n1289 VDD.n1196 4.5005
R75154 VDD.n1395 VDD.n1196 4.5005
R75155 VDD.n1288 VDD.n1196 4.5005
R75156 VDD.n1396 VDD.n1196 4.5005
R75157 VDD.n1286 VDD.n1196 4.5005
R75158 VDD.n1397 VDD.n1196 4.5005
R75159 VDD.n1285 VDD.n1196 4.5005
R75160 VDD.n1398 VDD.n1196 4.5005
R75161 VDD.n1283 VDD.n1196 4.5005
R75162 VDD.n1399 VDD.n1196 4.5005
R75163 VDD.n1282 VDD.n1196 4.5005
R75164 VDD.n1400 VDD.n1196 4.5005
R75165 VDD.n1280 VDD.n1196 4.5005
R75166 VDD.n1401 VDD.n1196 4.5005
R75167 VDD.n1279 VDD.n1196 4.5005
R75168 VDD.n1402 VDD.n1196 4.5005
R75169 VDD.n1277 VDD.n1196 4.5005
R75170 VDD.n1403 VDD.n1196 4.5005
R75171 VDD.n1276 VDD.n1196 4.5005
R75172 VDD.n1404 VDD.n1196 4.5005
R75173 VDD.n1274 VDD.n1196 4.5005
R75174 VDD.n1405 VDD.n1196 4.5005
R75175 VDD.n1273 VDD.n1196 4.5005
R75176 VDD.n1406 VDD.n1196 4.5005
R75177 VDD.n1271 VDD.n1196 4.5005
R75178 VDD.n1407 VDD.n1196 4.5005
R75179 VDD.n1270 VDD.n1196 4.5005
R75180 VDD.n1408 VDD.n1196 4.5005
R75181 VDD.n1268 VDD.n1196 4.5005
R75182 VDD.n1409 VDD.n1196 4.5005
R75183 VDD.n1267 VDD.n1196 4.5005
R75184 VDD.n1410 VDD.n1196 4.5005
R75185 VDD.n1265 VDD.n1196 4.5005
R75186 VDD.n1411 VDD.n1196 4.5005
R75187 VDD.n1264 VDD.n1196 4.5005
R75188 VDD.n1412 VDD.n1196 4.5005
R75189 VDD.n1262 VDD.n1196 4.5005
R75190 VDD.n1413 VDD.n1196 4.5005
R75191 VDD.n1261 VDD.n1196 4.5005
R75192 VDD.n1414 VDD.n1196 4.5005
R75193 VDD.n1415 VDD.n1196 4.5005
R75194 VDD.n1674 VDD.n1196 4.5005
R75195 VDD.n1676 VDD.n1193 4.5005
R75196 VDD.n1341 VDD.n1193 4.5005
R75197 VDD.n1342 VDD.n1193 4.5005
R75198 VDD.n1340 VDD.n1193 4.5005
R75199 VDD.n1344 VDD.n1193 4.5005
R75200 VDD.n1339 VDD.n1193 4.5005
R75201 VDD.n1345 VDD.n1193 4.5005
R75202 VDD.n1338 VDD.n1193 4.5005
R75203 VDD.n1347 VDD.n1193 4.5005
R75204 VDD.n1337 VDD.n1193 4.5005
R75205 VDD.n1348 VDD.n1193 4.5005
R75206 VDD.n1336 VDD.n1193 4.5005
R75207 VDD.n1350 VDD.n1193 4.5005
R75208 VDD.n1335 VDD.n1193 4.5005
R75209 VDD.n1351 VDD.n1193 4.5005
R75210 VDD.n1334 VDD.n1193 4.5005
R75211 VDD.n1353 VDD.n1193 4.5005
R75212 VDD.n1333 VDD.n1193 4.5005
R75213 VDD.n1354 VDD.n1193 4.5005
R75214 VDD.n1332 VDD.n1193 4.5005
R75215 VDD.n1356 VDD.n1193 4.5005
R75216 VDD.n1331 VDD.n1193 4.5005
R75217 VDD.n1357 VDD.n1193 4.5005
R75218 VDD.n1330 VDD.n1193 4.5005
R75219 VDD.n1359 VDD.n1193 4.5005
R75220 VDD.n1329 VDD.n1193 4.5005
R75221 VDD.n1360 VDD.n1193 4.5005
R75222 VDD.n1328 VDD.n1193 4.5005
R75223 VDD.n1362 VDD.n1193 4.5005
R75224 VDD.n1327 VDD.n1193 4.5005
R75225 VDD.n1363 VDD.n1193 4.5005
R75226 VDD.n1326 VDD.n1193 4.5005
R75227 VDD.n1365 VDD.n1193 4.5005
R75228 VDD.n1325 VDD.n1193 4.5005
R75229 VDD.n1366 VDD.n1193 4.5005
R75230 VDD.n1324 VDD.n1193 4.5005
R75231 VDD.n1368 VDD.n1193 4.5005
R75232 VDD.n1323 VDD.n1193 4.5005
R75233 VDD.n1369 VDD.n1193 4.5005
R75234 VDD.n1322 VDD.n1193 4.5005
R75235 VDD.n1371 VDD.n1193 4.5005
R75236 VDD.n1321 VDD.n1193 4.5005
R75237 VDD.n1372 VDD.n1193 4.5005
R75238 VDD.n1320 VDD.n1193 4.5005
R75239 VDD.n1374 VDD.n1193 4.5005
R75240 VDD.n1319 VDD.n1193 4.5005
R75241 VDD.n1375 VDD.n1193 4.5005
R75242 VDD.n1318 VDD.n1193 4.5005
R75243 VDD.n1376 VDD.n1193 4.5005
R75244 VDD.n1316 VDD.n1193 4.5005
R75245 VDD.n1377 VDD.n1193 4.5005
R75246 VDD.n1315 VDD.n1193 4.5005
R75247 VDD.n1378 VDD.n1193 4.5005
R75248 VDD.n1313 VDD.n1193 4.5005
R75249 VDD.n1379 VDD.n1193 4.5005
R75250 VDD.n1312 VDD.n1193 4.5005
R75251 VDD.n1380 VDD.n1193 4.5005
R75252 VDD.n1310 VDD.n1193 4.5005
R75253 VDD.n1381 VDD.n1193 4.5005
R75254 VDD.n1309 VDD.n1193 4.5005
R75255 VDD.n1382 VDD.n1193 4.5005
R75256 VDD.n1307 VDD.n1193 4.5005
R75257 VDD.n1383 VDD.n1193 4.5005
R75258 VDD.n1306 VDD.n1193 4.5005
R75259 VDD.n1384 VDD.n1193 4.5005
R75260 VDD.n1304 VDD.n1193 4.5005
R75261 VDD.n1385 VDD.n1193 4.5005
R75262 VDD.n1303 VDD.n1193 4.5005
R75263 VDD.n1386 VDD.n1193 4.5005
R75264 VDD.n1301 VDD.n1193 4.5005
R75265 VDD.n1387 VDD.n1193 4.5005
R75266 VDD.n1300 VDD.n1193 4.5005
R75267 VDD.n1388 VDD.n1193 4.5005
R75268 VDD.n1298 VDD.n1193 4.5005
R75269 VDD.n1389 VDD.n1193 4.5005
R75270 VDD.n1297 VDD.n1193 4.5005
R75271 VDD.n1390 VDD.n1193 4.5005
R75272 VDD.n1295 VDD.n1193 4.5005
R75273 VDD.n1391 VDD.n1193 4.5005
R75274 VDD.n1294 VDD.n1193 4.5005
R75275 VDD.n1392 VDD.n1193 4.5005
R75276 VDD.n1292 VDD.n1193 4.5005
R75277 VDD.n1393 VDD.n1193 4.5005
R75278 VDD.n1291 VDD.n1193 4.5005
R75279 VDD.n1394 VDD.n1193 4.5005
R75280 VDD.n1289 VDD.n1193 4.5005
R75281 VDD.n1395 VDD.n1193 4.5005
R75282 VDD.n1288 VDD.n1193 4.5005
R75283 VDD.n1396 VDD.n1193 4.5005
R75284 VDD.n1286 VDD.n1193 4.5005
R75285 VDD.n1397 VDD.n1193 4.5005
R75286 VDD.n1285 VDD.n1193 4.5005
R75287 VDD.n1398 VDD.n1193 4.5005
R75288 VDD.n1283 VDD.n1193 4.5005
R75289 VDD.n1399 VDD.n1193 4.5005
R75290 VDD.n1282 VDD.n1193 4.5005
R75291 VDD.n1400 VDD.n1193 4.5005
R75292 VDD.n1280 VDD.n1193 4.5005
R75293 VDD.n1401 VDD.n1193 4.5005
R75294 VDD.n1279 VDD.n1193 4.5005
R75295 VDD.n1402 VDD.n1193 4.5005
R75296 VDD.n1277 VDD.n1193 4.5005
R75297 VDD.n1403 VDD.n1193 4.5005
R75298 VDD.n1276 VDD.n1193 4.5005
R75299 VDD.n1404 VDD.n1193 4.5005
R75300 VDD.n1274 VDD.n1193 4.5005
R75301 VDD.n1405 VDD.n1193 4.5005
R75302 VDD.n1273 VDD.n1193 4.5005
R75303 VDD.n1406 VDD.n1193 4.5005
R75304 VDD.n1271 VDD.n1193 4.5005
R75305 VDD.n1407 VDD.n1193 4.5005
R75306 VDD.n1270 VDD.n1193 4.5005
R75307 VDD.n1408 VDD.n1193 4.5005
R75308 VDD.n1268 VDD.n1193 4.5005
R75309 VDD.n1409 VDD.n1193 4.5005
R75310 VDD.n1267 VDD.n1193 4.5005
R75311 VDD.n1410 VDD.n1193 4.5005
R75312 VDD.n1265 VDD.n1193 4.5005
R75313 VDD.n1411 VDD.n1193 4.5005
R75314 VDD.n1264 VDD.n1193 4.5005
R75315 VDD.n1412 VDD.n1193 4.5005
R75316 VDD.n1262 VDD.n1193 4.5005
R75317 VDD.n1413 VDD.n1193 4.5005
R75318 VDD.n1261 VDD.n1193 4.5005
R75319 VDD.n1414 VDD.n1193 4.5005
R75320 VDD.n1415 VDD.n1193 4.5005
R75321 VDD.n1674 VDD.n1193 4.5005
R75322 VDD.n1676 VDD.n1197 4.5005
R75323 VDD.n1341 VDD.n1197 4.5005
R75324 VDD.n1342 VDD.n1197 4.5005
R75325 VDD.n1340 VDD.n1197 4.5005
R75326 VDD.n1344 VDD.n1197 4.5005
R75327 VDD.n1339 VDD.n1197 4.5005
R75328 VDD.n1345 VDD.n1197 4.5005
R75329 VDD.n1338 VDD.n1197 4.5005
R75330 VDD.n1347 VDD.n1197 4.5005
R75331 VDD.n1337 VDD.n1197 4.5005
R75332 VDD.n1348 VDD.n1197 4.5005
R75333 VDD.n1336 VDD.n1197 4.5005
R75334 VDD.n1350 VDD.n1197 4.5005
R75335 VDD.n1335 VDD.n1197 4.5005
R75336 VDD.n1351 VDD.n1197 4.5005
R75337 VDD.n1334 VDD.n1197 4.5005
R75338 VDD.n1353 VDD.n1197 4.5005
R75339 VDD.n1333 VDD.n1197 4.5005
R75340 VDD.n1354 VDD.n1197 4.5005
R75341 VDD.n1332 VDD.n1197 4.5005
R75342 VDD.n1356 VDD.n1197 4.5005
R75343 VDD.n1331 VDD.n1197 4.5005
R75344 VDD.n1357 VDD.n1197 4.5005
R75345 VDD.n1330 VDD.n1197 4.5005
R75346 VDD.n1359 VDD.n1197 4.5005
R75347 VDD.n1329 VDD.n1197 4.5005
R75348 VDD.n1360 VDD.n1197 4.5005
R75349 VDD.n1328 VDD.n1197 4.5005
R75350 VDD.n1362 VDD.n1197 4.5005
R75351 VDD.n1327 VDD.n1197 4.5005
R75352 VDD.n1363 VDD.n1197 4.5005
R75353 VDD.n1326 VDD.n1197 4.5005
R75354 VDD.n1365 VDD.n1197 4.5005
R75355 VDD.n1325 VDD.n1197 4.5005
R75356 VDD.n1366 VDD.n1197 4.5005
R75357 VDD.n1324 VDD.n1197 4.5005
R75358 VDD.n1368 VDD.n1197 4.5005
R75359 VDD.n1323 VDD.n1197 4.5005
R75360 VDD.n1369 VDD.n1197 4.5005
R75361 VDD.n1322 VDD.n1197 4.5005
R75362 VDD.n1371 VDD.n1197 4.5005
R75363 VDD.n1321 VDD.n1197 4.5005
R75364 VDD.n1372 VDD.n1197 4.5005
R75365 VDD.n1320 VDD.n1197 4.5005
R75366 VDD.n1374 VDD.n1197 4.5005
R75367 VDD.n1319 VDD.n1197 4.5005
R75368 VDD.n1375 VDD.n1197 4.5005
R75369 VDD.n1318 VDD.n1197 4.5005
R75370 VDD.n1376 VDD.n1197 4.5005
R75371 VDD.n1316 VDD.n1197 4.5005
R75372 VDD.n1377 VDD.n1197 4.5005
R75373 VDD.n1315 VDD.n1197 4.5005
R75374 VDD.n1378 VDD.n1197 4.5005
R75375 VDD.n1313 VDD.n1197 4.5005
R75376 VDD.n1379 VDD.n1197 4.5005
R75377 VDD.n1312 VDD.n1197 4.5005
R75378 VDD.n1380 VDD.n1197 4.5005
R75379 VDD.n1310 VDD.n1197 4.5005
R75380 VDD.n1381 VDD.n1197 4.5005
R75381 VDD.n1309 VDD.n1197 4.5005
R75382 VDD.n1382 VDD.n1197 4.5005
R75383 VDD.n1307 VDD.n1197 4.5005
R75384 VDD.n1383 VDD.n1197 4.5005
R75385 VDD.n1306 VDD.n1197 4.5005
R75386 VDD.n1384 VDD.n1197 4.5005
R75387 VDD.n1304 VDD.n1197 4.5005
R75388 VDD.n1385 VDD.n1197 4.5005
R75389 VDD.n1303 VDD.n1197 4.5005
R75390 VDD.n1386 VDD.n1197 4.5005
R75391 VDD.n1301 VDD.n1197 4.5005
R75392 VDD.n1387 VDD.n1197 4.5005
R75393 VDD.n1300 VDD.n1197 4.5005
R75394 VDD.n1388 VDD.n1197 4.5005
R75395 VDD.n1298 VDD.n1197 4.5005
R75396 VDD.n1389 VDD.n1197 4.5005
R75397 VDD.n1297 VDD.n1197 4.5005
R75398 VDD.n1390 VDD.n1197 4.5005
R75399 VDD.n1295 VDD.n1197 4.5005
R75400 VDD.n1391 VDD.n1197 4.5005
R75401 VDD.n1294 VDD.n1197 4.5005
R75402 VDD.n1392 VDD.n1197 4.5005
R75403 VDD.n1292 VDD.n1197 4.5005
R75404 VDD.n1393 VDD.n1197 4.5005
R75405 VDD.n1291 VDD.n1197 4.5005
R75406 VDD.n1394 VDD.n1197 4.5005
R75407 VDD.n1289 VDD.n1197 4.5005
R75408 VDD.n1395 VDD.n1197 4.5005
R75409 VDD.n1288 VDD.n1197 4.5005
R75410 VDD.n1396 VDD.n1197 4.5005
R75411 VDD.n1286 VDD.n1197 4.5005
R75412 VDD.n1397 VDD.n1197 4.5005
R75413 VDD.n1285 VDD.n1197 4.5005
R75414 VDD.n1398 VDD.n1197 4.5005
R75415 VDD.n1283 VDD.n1197 4.5005
R75416 VDD.n1399 VDD.n1197 4.5005
R75417 VDD.n1282 VDD.n1197 4.5005
R75418 VDD.n1400 VDD.n1197 4.5005
R75419 VDD.n1280 VDD.n1197 4.5005
R75420 VDD.n1401 VDD.n1197 4.5005
R75421 VDD.n1279 VDD.n1197 4.5005
R75422 VDD.n1402 VDD.n1197 4.5005
R75423 VDD.n1277 VDD.n1197 4.5005
R75424 VDD.n1403 VDD.n1197 4.5005
R75425 VDD.n1276 VDD.n1197 4.5005
R75426 VDD.n1404 VDD.n1197 4.5005
R75427 VDD.n1274 VDD.n1197 4.5005
R75428 VDD.n1405 VDD.n1197 4.5005
R75429 VDD.n1273 VDD.n1197 4.5005
R75430 VDD.n1406 VDD.n1197 4.5005
R75431 VDD.n1271 VDD.n1197 4.5005
R75432 VDD.n1407 VDD.n1197 4.5005
R75433 VDD.n1270 VDD.n1197 4.5005
R75434 VDD.n1408 VDD.n1197 4.5005
R75435 VDD.n1268 VDD.n1197 4.5005
R75436 VDD.n1409 VDD.n1197 4.5005
R75437 VDD.n1267 VDD.n1197 4.5005
R75438 VDD.n1410 VDD.n1197 4.5005
R75439 VDD.n1265 VDD.n1197 4.5005
R75440 VDD.n1411 VDD.n1197 4.5005
R75441 VDD.n1264 VDD.n1197 4.5005
R75442 VDD.n1412 VDD.n1197 4.5005
R75443 VDD.n1262 VDD.n1197 4.5005
R75444 VDD.n1413 VDD.n1197 4.5005
R75445 VDD.n1261 VDD.n1197 4.5005
R75446 VDD.n1414 VDD.n1197 4.5005
R75447 VDD.n1415 VDD.n1197 4.5005
R75448 VDD.n1674 VDD.n1197 4.5005
R75449 VDD.n1676 VDD.n1192 4.5005
R75450 VDD.n1341 VDD.n1192 4.5005
R75451 VDD.n1342 VDD.n1192 4.5005
R75452 VDD.n1340 VDD.n1192 4.5005
R75453 VDD.n1344 VDD.n1192 4.5005
R75454 VDD.n1339 VDD.n1192 4.5005
R75455 VDD.n1345 VDD.n1192 4.5005
R75456 VDD.n1338 VDD.n1192 4.5005
R75457 VDD.n1347 VDD.n1192 4.5005
R75458 VDD.n1337 VDD.n1192 4.5005
R75459 VDD.n1348 VDD.n1192 4.5005
R75460 VDD.n1336 VDD.n1192 4.5005
R75461 VDD.n1350 VDD.n1192 4.5005
R75462 VDD.n1335 VDD.n1192 4.5005
R75463 VDD.n1351 VDD.n1192 4.5005
R75464 VDD.n1334 VDD.n1192 4.5005
R75465 VDD.n1353 VDD.n1192 4.5005
R75466 VDD.n1333 VDD.n1192 4.5005
R75467 VDD.n1354 VDD.n1192 4.5005
R75468 VDD.n1332 VDD.n1192 4.5005
R75469 VDD.n1356 VDD.n1192 4.5005
R75470 VDD.n1331 VDD.n1192 4.5005
R75471 VDD.n1357 VDD.n1192 4.5005
R75472 VDD.n1330 VDD.n1192 4.5005
R75473 VDD.n1359 VDD.n1192 4.5005
R75474 VDD.n1329 VDD.n1192 4.5005
R75475 VDD.n1360 VDD.n1192 4.5005
R75476 VDD.n1328 VDD.n1192 4.5005
R75477 VDD.n1362 VDD.n1192 4.5005
R75478 VDD.n1327 VDD.n1192 4.5005
R75479 VDD.n1363 VDD.n1192 4.5005
R75480 VDD.n1326 VDD.n1192 4.5005
R75481 VDD.n1365 VDD.n1192 4.5005
R75482 VDD.n1325 VDD.n1192 4.5005
R75483 VDD.n1366 VDD.n1192 4.5005
R75484 VDD.n1324 VDD.n1192 4.5005
R75485 VDD.n1368 VDD.n1192 4.5005
R75486 VDD.n1323 VDD.n1192 4.5005
R75487 VDD.n1369 VDD.n1192 4.5005
R75488 VDD.n1322 VDD.n1192 4.5005
R75489 VDD.n1371 VDD.n1192 4.5005
R75490 VDD.n1321 VDD.n1192 4.5005
R75491 VDD.n1372 VDD.n1192 4.5005
R75492 VDD.n1320 VDD.n1192 4.5005
R75493 VDD.n1374 VDD.n1192 4.5005
R75494 VDD.n1319 VDD.n1192 4.5005
R75495 VDD.n1375 VDD.n1192 4.5005
R75496 VDD.n1318 VDD.n1192 4.5005
R75497 VDD.n1376 VDD.n1192 4.5005
R75498 VDD.n1316 VDD.n1192 4.5005
R75499 VDD.n1377 VDD.n1192 4.5005
R75500 VDD.n1315 VDD.n1192 4.5005
R75501 VDD.n1378 VDD.n1192 4.5005
R75502 VDD.n1313 VDD.n1192 4.5005
R75503 VDD.n1379 VDD.n1192 4.5005
R75504 VDD.n1312 VDD.n1192 4.5005
R75505 VDD.n1380 VDD.n1192 4.5005
R75506 VDD.n1310 VDD.n1192 4.5005
R75507 VDD.n1381 VDD.n1192 4.5005
R75508 VDD.n1309 VDD.n1192 4.5005
R75509 VDD.n1382 VDD.n1192 4.5005
R75510 VDD.n1307 VDD.n1192 4.5005
R75511 VDD.n1383 VDD.n1192 4.5005
R75512 VDD.n1306 VDD.n1192 4.5005
R75513 VDD.n1384 VDD.n1192 4.5005
R75514 VDD.n1304 VDD.n1192 4.5005
R75515 VDD.n1385 VDD.n1192 4.5005
R75516 VDD.n1303 VDD.n1192 4.5005
R75517 VDD.n1386 VDD.n1192 4.5005
R75518 VDD.n1301 VDD.n1192 4.5005
R75519 VDD.n1387 VDD.n1192 4.5005
R75520 VDD.n1300 VDD.n1192 4.5005
R75521 VDD.n1388 VDD.n1192 4.5005
R75522 VDD.n1298 VDD.n1192 4.5005
R75523 VDD.n1389 VDD.n1192 4.5005
R75524 VDD.n1297 VDD.n1192 4.5005
R75525 VDD.n1390 VDD.n1192 4.5005
R75526 VDD.n1295 VDD.n1192 4.5005
R75527 VDD.n1391 VDD.n1192 4.5005
R75528 VDD.n1294 VDD.n1192 4.5005
R75529 VDD.n1392 VDD.n1192 4.5005
R75530 VDD.n1292 VDD.n1192 4.5005
R75531 VDD.n1393 VDD.n1192 4.5005
R75532 VDD.n1291 VDD.n1192 4.5005
R75533 VDD.n1394 VDD.n1192 4.5005
R75534 VDD.n1289 VDD.n1192 4.5005
R75535 VDD.n1395 VDD.n1192 4.5005
R75536 VDD.n1288 VDD.n1192 4.5005
R75537 VDD.n1396 VDD.n1192 4.5005
R75538 VDD.n1286 VDD.n1192 4.5005
R75539 VDD.n1397 VDD.n1192 4.5005
R75540 VDD.n1285 VDD.n1192 4.5005
R75541 VDD.n1398 VDD.n1192 4.5005
R75542 VDD.n1283 VDD.n1192 4.5005
R75543 VDD.n1399 VDD.n1192 4.5005
R75544 VDD.n1282 VDD.n1192 4.5005
R75545 VDD.n1400 VDD.n1192 4.5005
R75546 VDD.n1280 VDD.n1192 4.5005
R75547 VDD.n1401 VDD.n1192 4.5005
R75548 VDD.n1279 VDD.n1192 4.5005
R75549 VDD.n1402 VDD.n1192 4.5005
R75550 VDD.n1277 VDD.n1192 4.5005
R75551 VDD.n1403 VDD.n1192 4.5005
R75552 VDD.n1276 VDD.n1192 4.5005
R75553 VDD.n1404 VDD.n1192 4.5005
R75554 VDD.n1274 VDD.n1192 4.5005
R75555 VDD.n1405 VDD.n1192 4.5005
R75556 VDD.n1273 VDD.n1192 4.5005
R75557 VDD.n1406 VDD.n1192 4.5005
R75558 VDD.n1271 VDD.n1192 4.5005
R75559 VDD.n1407 VDD.n1192 4.5005
R75560 VDD.n1270 VDD.n1192 4.5005
R75561 VDD.n1408 VDD.n1192 4.5005
R75562 VDD.n1268 VDD.n1192 4.5005
R75563 VDD.n1409 VDD.n1192 4.5005
R75564 VDD.n1267 VDD.n1192 4.5005
R75565 VDD.n1410 VDD.n1192 4.5005
R75566 VDD.n1265 VDD.n1192 4.5005
R75567 VDD.n1411 VDD.n1192 4.5005
R75568 VDD.n1264 VDD.n1192 4.5005
R75569 VDD.n1412 VDD.n1192 4.5005
R75570 VDD.n1262 VDD.n1192 4.5005
R75571 VDD.n1413 VDD.n1192 4.5005
R75572 VDD.n1261 VDD.n1192 4.5005
R75573 VDD.n1414 VDD.n1192 4.5005
R75574 VDD.n1415 VDD.n1192 4.5005
R75575 VDD.n1674 VDD.n1192 4.5005
R75576 VDD.n1676 VDD.n1198 4.5005
R75577 VDD.n1341 VDD.n1198 4.5005
R75578 VDD.n1342 VDD.n1198 4.5005
R75579 VDD.n1340 VDD.n1198 4.5005
R75580 VDD.n1344 VDD.n1198 4.5005
R75581 VDD.n1339 VDD.n1198 4.5005
R75582 VDD.n1345 VDD.n1198 4.5005
R75583 VDD.n1338 VDD.n1198 4.5005
R75584 VDD.n1347 VDD.n1198 4.5005
R75585 VDD.n1337 VDD.n1198 4.5005
R75586 VDD.n1348 VDD.n1198 4.5005
R75587 VDD.n1336 VDD.n1198 4.5005
R75588 VDD.n1350 VDD.n1198 4.5005
R75589 VDD.n1335 VDD.n1198 4.5005
R75590 VDD.n1351 VDD.n1198 4.5005
R75591 VDD.n1334 VDD.n1198 4.5005
R75592 VDD.n1353 VDD.n1198 4.5005
R75593 VDD.n1333 VDD.n1198 4.5005
R75594 VDD.n1354 VDD.n1198 4.5005
R75595 VDD.n1332 VDD.n1198 4.5005
R75596 VDD.n1356 VDD.n1198 4.5005
R75597 VDD.n1331 VDD.n1198 4.5005
R75598 VDD.n1357 VDD.n1198 4.5005
R75599 VDD.n1330 VDD.n1198 4.5005
R75600 VDD.n1359 VDD.n1198 4.5005
R75601 VDD.n1329 VDD.n1198 4.5005
R75602 VDD.n1360 VDD.n1198 4.5005
R75603 VDD.n1328 VDD.n1198 4.5005
R75604 VDD.n1362 VDD.n1198 4.5005
R75605 VDD.n1327 VDD.n1198 4.5005
R75606 VDD.n1363 VDD.n1198 4.5005
R75607 VDD.n1326 VDD.n1198 4.5005
R75608 VDD.n1365 VDD.n1198 4.5005
R75609 VDD.n1325 VDD.n1198 4.5005
R75610 VDD.n1366 VDD.n1198 4.5005
R75611 VDD.n1324 VDD.n1198 4.5005
R75612 VDD.n1368 VDD.n1198 4.5005
R75613 VDD.n1323 VDD.n1198 4.5005
R75614 VDD.n1369 VDD.n1198 4.5005
R75615 VDD.n1322 VDD.n1198 4.5005
R75616 VDD.n1371 VDD.n1198 4.5005
R75617 VDD.n1321 VDD.n1198 4.5005
R75618 VDD.n1372 VDD.n1198 4.5005
R75619 VDD.n1320 VDD.n1198 4.5005
R75620 VDD.n1374 VDD.n1198 4.5005
R75621 VDD.n1319 VDD.n1198 4.5005
R75622 VDD.n1375 VDD.n1198 4.5005
R75623 VDD.n1318 VDD.n1198 4.5005
R75624 VDD.n1376 VDD.n1198 4.5005
R75625 VDD.n1316 VDD.n1198 4.5005
R75626 VDD.n1377 VDD.n1198 4.5005
R75627 VDD.n1315 VDD.n1198 4.5005
R75628 VDD.n1378 VDD.n1198 4.5005
R75629 VDD.n1313 VDD.n1198 4.5005
R75630 VDD.n1379 VDD.n1198 4.5005
R75631 VDD.n1312 VDD.n1198 4.5005
R75632 VDD.n1380 VDD.n1198 4.5005
R75633 VDD.n1310 VDD.n1198 4.5005
R75634 VDD.n1381 VDD.n1198 4.5005
R75635 VDD.n1309 VDD.n1198 4.5005
R75636 VDD.n1382 VDD.n1198 4.5005
R75637 VDD.n1307 VDD.n1198 4.5005
R75638 VDD.n1383 VDD.n1198 4.5005
R75639 VDD.n1306 VDD.n1198 4.5005
R75640 VDD.n1384 VDD.n1198 4.5005
R75641 VDD.n1304 VDD.n1198 4.5005
R75642 VDD.n1385 VDD.n1198 4.5005
R75643 VDD.n1303 VDD.n1198 4.5005
R75644 VDD.n1386 VDD.n1198 4.5005
R75645 VDD.n1301 VDD.n1198 4.5005
R75646 VDD.n1387 VDD.n1198 4.5005
R75647 VDD.n1300 VDD.n1198 4.5005
R75648 VDD.n1388 VDD.n1198 4.5005
R75649 VDD.n1298 VDD.n1198 4.5005
R75650 VDD.n1389 VDD.n1198 4.5005
R75651 VDD.n1297 VDD.n1198 4.5005
R75652 VDD.n1390 VDD.n1198 4.5005
R75653 VDD.n1295 VDD.n1198 4.5005
R75654 VDD.n1391 VDD.n1198 4.5005
R75655 VDD.n1294 VDD.n1198 4.5005
R75656 VDD.n1392 VDD.n1198 4.5005
R75657 VDD.n1292 VDD.n1198 4.5005
R75658 VDD.n1393 VDD.n1198 4.5005
R75659 VDD.n1291 VDD.n1198 4.5005
R75660 VDD.n1394 VDD.n1198 4.5005
R75661 VDD.n1289 VDD.n1198 4.5005
R75662 VDD.n1395 VDD.n1198 4.5005
R75663 VDD.n1288 VDD.n1198 4.5005
R75664 VDD.n1396 VDD.n1198 4.5005
R75665 VDD.n1286 VDD.n1198 4.5005
R75666 VDD.n1397 VDD.n1198 4.5005
R75667 VDD.n1285 VDD.n1198 4.5005
R75668 VDD.n1398 VDD.n1198 4.5005
R75669 VDD.n1283 VDD.n1198 4.5005
R75670 VDD.n1399 VDD.n1198 4.5005
R75671 VDD.n1282 VDD.n1198 4.5005
R75672 VDD.n1400 VDD.n1198 4.5005
R75673 VDD.n1280 VDD.n1198 4.5005
R75674 VDD.n1401 VDD.n1198 4.5005
R75675 VDD.n1279 VDD.n1198 4.5005
R75676 VDD.n1402 VDD.n1198 4.5005
R75677 VDD.n1277 VDD.n1198 4.5005
R75678 VDD.n1403 VDD.n1198 4.5005
R75679 VDD.n1276 VDD.n1198 4.5005
R75680 VDD.n1404 VDD.n1198 4.5005
R75681 VDD.n1274 VDD.n1198 4.5005
R75682 VDD.n1405 VDD.n1198 4.5005
R75683 VDD.n1273 VDD.n1198 4.5005
R75684 VDD.n1406 VDD.n1198 4.5005
R75685 VDD.n1271 VDD.n1198 4.5005
R75686 VDD.n1407 VDD.n1198 4.5005
R75687 VDD.n1270 VDD.n1198 4.5005
R75688 VDD.n1408 VDD.n1198 4.5005
R75689 VDD.n1268 VDD.n1198 4.5005
R75690 VDD.n1409 VDD.n1198 4.5005
R75691 VDD.n1267 VDD.n1198 4.5005
R75692 VDD.n1410 VDD.n1198 4.5005
R75693 VDD.n1265 VDD.n1198 4.5005
R75694 VDD.n1411 VDD.n1198 4.5005
R75695 VDD.n1264 VDD.n1198 4.5005
R75696 VDD.n1412 VDD.n1198 4.5005
R75697 VDD.n1262 VDD.n1198 4.5005
R75698 VDD.n1413 VDD.n1198 4.5005
R75699 VDD.n1261 VDD.n1198 4.5005
R75700 VDD.n1414 VDD.n1198 4.5005
R75701 VDD.n1415 VDD.n1198 4.5005
R75702 VDD.n1674 VDD.n1198 4.5005
R75703 VDD.n1676 VDD.n1191 4.5005
R75704 VDD.n1341 VDD.n1191 4.5005
R75705 VDD.n1342 VDD.n1191 4.5005
R75706 VDD.n1340 VDD.n1191 4.5005
R75707 VDD.n1344 VDD.n1191 4.5005
R75708 VDD.n1339 VDD.n1191 4.5005
R75709 VDD.n1345 VDD.n1191 4.5005
R75710 VDD.n1338 VDD.n1191 4.5005
R75711 VDD.n1347 VDD.n1191 4.5005
R75712 VDD.n1337 VDD.n1191 4.5005
R75713 VDD.n1348 VDD.n1191 4.5005
R75714 VDD.n1336 VDD.n1191 4.5005
R75715 VDD.n1350 VDD.n1191 4.5005
R75716 VDD.n1335 VDD.n1191 4.5005
R75717 VDD.n1351 VDD.n1191 4.5005
R75718 VDD.n1334 VDD.n1191 4.5005
R75719 VDD.n1353 VDD.n1191 4.5005
R75720 VDD.n1333 VDD.n1191 4.5005
R75721 VDD.n1354 VDD.n1191 4.5005
R75722 VDD.n1332 VDD.n1191 4.5005
R75723 VDD.n1356 VDD.n1191 4.5005
R75724 VDD.n1331 VDD.n1191 4.5005
R75725 VDD.n1357 VDD.n1191 4.5005
R75726 VDD.n1330 VDD.n1191 4.5005
R75727 VDD.n1359 VDD.n1191 4.5005
R75728 VDD.n1329 VDD.n1191 4.5005
R75729 VDD.n1360 VDD.n1191 4.5005
R75730 VDD.n1328 VDD.n1191 4.5005
R75731 VDD.n1362 VDD.n1191 4.5005
R75732 VDD.n1327 VDD.n1191 4.5005
R75733 VDD.n1363 VDD.n1191 4.5005
R75734 VDD.n1326 VDD.n1191 4.5005
R75735 VDD.n1365 VDD.n1191 4.5005
R75736 VDD.n1325 VDD.n1191 4.5005
R75737 VDD.n1366 VDD.n1191 4.5005
R75738 VDD.n1324 VDD.n1191 4.5005
R75739 VDD.n1368 VDD.n1191 4.5005
R75740 VDD.n1323 VDD.n1191 4.5005
R75741 VDD.n1369 VDD.n1191 4.5005
R75742 VDD.n1322 VDD.n1191 4.5005
R75743 VDD.n1371 VDD.n1191 4.5005
R75744 VDD.n1321 VDD.n1191 4.5005
R75745 VDD.n1372 VDD.n1191 4.5005
R75746 VDD.n1320 VDD.n1191 4.5005
R75747 VDD.n1374 VDD.n1191 4.5005
R75748 VDD.n1319 VDD.n1191 4.5005
R75749 VDD.n1375 VDD.n1191 4.5005
R75750 VDD.n1318 VDD.n1191 4.5005
R75751 VDD.n1376 VDD.n1191 4.5005
R75752 VDD.n1316 VDD.n1191 4.5005
R75753 VDD.n1377 VDD.n1191 4.5005
R75754 VDD.n1315 VDD.n1191 4.5005
R75755 VDD.n1378 VDD.n1191 4.5005
R75756 VDD.n1313 VDD.n1191 4.5005
R75757 VDD.n1379 VDD.n1191 4.5005
R75758 VDD.n1312 VDD.n1191 4.5005
R75759 VDD.n1380 VDD.n1191 4.5005
R75760 VDD.n1310 VDD.n1191 4.5005
R75761 VDD.n1381 VDD.n1191 4.5005
R75762 VDD.n1309 VDD.n1191 4.5005
R75763 VDD.n1382 VDD.n1191 4.5005
R75764 VDD.n1307 VDD.n1191 4.5005
R75765 VDD.n1383 VDD.n1191 4.5005
R75766 VDD.n1306 VDD.n1191 4.5005
R75767 VDD.n1384 VDD.n1191 4.5005
R75768 VDD.n1304 VDD.n1191 4.5005
R75769 VDD.n1385 VDD.n1191 4.5005
R75770 VDD.n1303 VDD.n1191 4.5005
R75771 VDD.n1386 VDD.n1191 4.5005
R75772 VDD.n1301 VDD.n1191 4.5005
R75773 VDD.n1387 VDD.n1191 4.5005
R75774 VDD.n1300 VDD.n1191 4.5005
R75775 VDD.n1388 VDD.n1191 4.5005
R75776 VDD.n1298 VDD.n1191 4.5005
R75777 VDD.n1389 VDD.n1191 4.5005
R75778 VDD.n1297 VDD.n1191 4.5005
R75779 VDD.n1390 VDD.n1191 4.5005
R75780 VDD.n1295 VDD.n1191 4.5005
R75781 VDD.n1391 VDD.n1191 4.5005
R75782 VDD.n1294 VDD.n1191 4.5005
R75783 VDD.n1392 VDD.n1191 4.5005
R75784 VDD.n1292 VDD.n1191 4.5005
R75785 VDD.n1393 VDD.n1191 4.5005
R75786 VDD.n1291 VDD.n1191 4.5005
R75787 VDD.n1394 VDD.n1191 4.5005
R75788 VDD.n1289 VDD.n1191 4.5005
R75789 VDD.n1395 VDD.n1191 4.5005
R75790 VDD.n1288 VDD.n1191 4.5005
R75791 VDD.n1396 VDD.n1191 4.5005
R75792 VDD.n1286 VDD.n1191 4.5005
R75793 VDD.n1397 VDD.n1191 4.5005
R75794 VDD.n1285 VDD.n1191 4.5005
R75795 VDD.n1398 VDD.n1191 4.5005
R75796 VDD.n1283 VDD.n1191 4.5005
R75797 VDD.n1399 VDD.n1191 4.5005
R75798 VDD.n1282 VDD.n1191 4.5005
R75799 VDD.n1400 VDD.n1191 4.5005
R75800 VDD.n1280 VDD.n1191 4.5005
R75801 VDD.n1401 VDD.n1191 4.5005
R75802 VDD.n1279 VDD.n1191 4.5005
R75803 VDD.n1402 VDD.n1191 4.5005
R75804 VDD.n1277 VDD.n1191 4.5005
R75805 VDD.n1403 VDD.n1191 4.5005
R75806 VDD.n1276 VDD.n1191 4.5005
R75807 VDD.n1404 VDD.n1191 4.5005
R75808 VDD.n1274 VDD.n1191 4.5005
R75809 VDD.n1405 VDD.n1191 4.5005
R75810 VDD.n1273 VDD.n1191 4.5005
R75811 VDD.n1406 VDD.n1191 4.5005
R75812 VDD.n1271 VDD.n1191 4.5005
R75813 VDD.n1407 VDD.n1191 4.5005
R75814 VDD.n1270 VDD.n1191 4.5005
R75815 VDD.n1408 VDD.n1191 4.5005
R75816 VDD.n1268 VDD.n1191 4.5005
R75817 VDD.n1409 VDD.n1191 4.5005
R75818 VDD.n1267 VDD.n1191 4.5005
R75819 VDD.n1410 VDD.n1191 4.5005
R75820 VDD.n1265 VDD.n1191 4.5005
R75821 VDD.n1411 VDD.n1191 4.5005
R75822 VDD.n1264 VDD.n1191 4.5005
R75823 VDD.n1412 VDD.n1191 4.5005
R75824 VDD.n1262 VDD.n1191 4.5005
R75825 VDD.n1413 VDD.n1191 4.5005
R75826 VDD.n1261 VDD.n1191 4.5005
R75827 VDD.n1414 VDD.n1191 4.5005
R75828 VDD.n1415 VDD.n1191 4.5005
R75829 VDD.n1674 VDD.n1191 4.5005
R75830 VDD.n1676 VDD.n1199 4.5005
R75831 VDD.n1341 VDD.n1199 4.5005
R75832 VDD.n1342 VDD.n1199 4.5005
R75833 VDD.n1340 VDD.n1199 4.5005
R75834 VDD.n1344 VDD.n1199 4.5005
R75835 VDD.n1339 VDD.n1199 4.5005
R75836 VDD.n1345 VDD.n1199 4.5005
R75837 VDD.n1338 VDD.n1199 4.5005
R75838 VDD.n1347 VDD.n1199 4.5005
R75839 VDD.n1337 VDD.n1199 4.5005
R75840 VDD.n1348 VDD.n1199 4.5005
R75841 VDD.n1336 VDD.n1199 4.5005
R75842 VDD.n1350 VDD.n1199 4.5005
R75843 VDD.n1335 VDD.n1199 4.5005
R75844 VDD.n1351 VDD.n1199 4.5005
R75845 VDD.n1334 VDD.n1199 4.5005
R75846 VDD.n1353 VDD.n1199 4.5005
R75847 VDD.n1333 VDD.n1199 4.5005
R75848 VDD.n1354 VDD.n1199 4.5005
R75849 VDD.n1332 VDD.n1199 4.5005
R75850 VDD.n1356 VDD.n1199 4.5005
R75851 VDD.n1331 VDD.n1199 4.5005
R75852 VDD.n1357 VDD.n1199 4.5005
R75853 VDD.n1330 VDD.n1199 4.5005
R75854 VDD.n1359 VDD.n1199 4.5005
R75855 VDD.n1329 VDD.n1199 4.5005
R75856 VDD.n1360 VDD.n1199 4.5005
R75857 VDD.n1328 VDD.n1199 4.5005
R75858 VDD.n1362 VDD.n1199 4.5005
R75859 VDD.n1327 VDD.n1199 4.5005
R75860 VDD.n1363 VDD.n1199 4.5005
R75861 VDD.n1326 VDD.n1199 4.5005
R75862 VDD.n1365 VDD.n1199 4.5005
R75863 VDD.n1325 VDD.n1199 4.5005
R75864 VDD.n1366 VDD.n1199 4.5005
R75865 VDD.n1324 VDD.n1199 4.5005
R75866 VDD.n1368 VDD.n1199 4.5005
R75867 VDD.n1323 VDD.n1199 4.5005
R75868 VDD.n1369 VDD.n1199 4.5005
R75869 VDD.n1322 VDD.n1199 4.5005
R75870 VDD.n1371 VDD.n1199 4.5005
R75871 VDD.n1321 VDD.n1199 4.5005
R75872 VDD.n1372 VDD.n1199 4.5005
R75873 VDD.n1320 VDD.n1199 4.5005
R75874 VDD.n1374 VDD.n1199 4.5005
R75875 VDD.n1319 VDD.n1199 4.5005
R75876 VDD.n1375 VDD.n1199 4.5005
R75877 VDD.n1318 VDD.n1199 4.5005
R75878 VDD.n1376 VDD.n1199 4.5005
R75879 VDD.n1316 VDD.n1199 4.5005
R75880 VDD.n1377 VDD.n1199 4.5005
R75881 VDD.n1315 VDD.n1199 4.5005
R75882 VDD.n1378 VDD.n1199 4.5005
R75883 VDD.n1313 VDD.n1199 4.5005
R75884 VDD.n1379 VDD.n1199 4.5005
R75885 VDD.n1312 VDD.n1199 4.5005
R75886 VDD.n1380 VDD.n1199 4.5005
R75887 VDD.n1310 VDD.n1199 4.5005
R75888 VDD.n1381 VDD.n1199 4.5005
R75889 VDD.n1309 VDD.n1199 4.5005
R75890 VDD.n1382 VDD.n1199 4.5005
R75891 VDD.n1307 VDD.n1199 4.5005
R75892 VDD.n1383 VDD.n1199 4.5005
R75893 VDD.n1306 VDD.n1199 4.5005
R75894 VDD.n1384 VDD.n1199 4.5005
R75895 VDD.n1304 VDD.n1199 4.5005
R75896 VDD.n1385 VDD.n1199 4.5005
R75897 VDD.n1303 VDD.n1199 4.5005
R75898 VDD.n1386 VDD.n1199 4.5005
R75899 VDD.n1301 VDD.n1199 4.5005
R75900 VDD.n1387 VDD.n1199 4.5005
R75901 VDD.n1300 VDD.n1199 4.5005
R75902 VDD.n1388 VDD.n1199 4.5005
R75903 VDD.n1298 VDD.n1199 4.5005
R75904 VDD.n1389 VDD.n1199 4.5005
R75905 VDD.n1297 VDD.n1199 4.5005
R75906 VDD.n1390 VDD.n1199 4.5005
R75907 VDD.n1295 VDD.n1199 4.5005
R75908 VDD.n1391 VDD.n1199 4.5005
R75909 VDD.n1294 VDD.n1199 4.5005
R75910 VDD.n1392 VDD.n1199 4.5005
R75911 VDD.n1292 VDD.n1199 4.5005
R75912 VDD.n1393 VDD.n1199 4.5005
R75913 VDD.n1291 VDD.n1199 4.5005
R75914 VDD.n1394 VDD.n1199 4.5005
R75915 VDD.n1289 VDD.n1199 4.5005
R75916 VDD.n1395 VDD.n1199 4.5005
R75917 VDD.n1288 VDD.n1199 4.5005
R75918 VDD.n1396 VDD.n1199 4.5005
R75919 VDD.n1286 VDD.n1199 4.5005
R75920 VDD.n1397 VDD.n1199 4.5005
R75921 VDD.n1285 VDD.n1199 4.5005
R75922 VDD.n1398 VDD.n1199 4.5005
R75923 VDD.n1283 VDD.n1199 4.5005
R75924 VDD.n1399 VDD.n1199 4.5005
R75925 VDD.n1282 VDD.n1199 4.5005
R75926 VDD.n1400 VDD.n1199 4.5005
R75927 VDD.n1280 VDD.n1199 4.5005
R75928 VDD.n1401 VDD.n1199 4.5005
R75929 VDD.n1279 VDD.n1199 4.5005
R75930 VDD.n1402 VDD.n1199 4.5005
R75931 VDD.n1277 VDD.n1199 4.5005
R75932 VDD.n1403 VDD.n1199 4.5005
R75933 VDD.n1276 VDD.n1199 4.5005
R75934 VDD.n1404 VDD.n1199 4.5005
R75935 VDD.n1274 VDD.n1199 4.5005
R75936 VDD.n1405 VDD.n1199 4.5005
R75937 VDD.n1273 VDD.n1199 4.5005
R75938 VDD.n1406 VDD.n1199 4.5005
R75939 VDD.n1271 VDD.n1199 4.5005
R75940 VDD.n1407 VDD.n1199 4.5005
R75941 VDD.n1270 VDD.n1199 4.5005
R75942 VDD.n1408 VDD.n1199 4.5005
R75943 VDD.n1268 VDD.n1199 4.5005
R75944 VDD.n1409 VDD.n1199 4.5005
R75945 VDD.n1267 VDD.n1199 4.5005
R75946 VDD.n1410 VDD.n1199 4.5005
R75947 VDD.n1265 VDD.n1199 4.5005
R75948 VDD.n1411 VDD.n1199 4.5005
R75949 VDD.n1264 VDD.n1199 4.5005
R75950 VDD.n1412 VDD.n1199 4.5005
R75951 VDD.n1262 VDD.n1199 4.5005
R75952 VDD.n1413 VDD.n1199 4.5005
R75953 VDD.n1261 VDD.n1199 4.5005
R75954 VDD.n1414 VDD.n1199 4.5005
R75955 VDD.n1415 VDD.n1199 4.5005
R75956 VDD.n1674 VDD.n1199 4.5005
R75957 VDD.n1676 VDD.n1190 4.5005
R75958 VDD.n1341 VDD.n1190 4.5005
R75959 VDD.n1342 VDD.n1190 4.5005
R75960 VDD.n1340 VDD.n1190 4.5005
R75961 VDD.n1344 VDD.n1190 4.5005
R75962 VDD.n1339 VDD.n1190 4.5005
R75963 VDD.n1345 VDD.n1190 4.5005
R75964 VDD.n1338 VDD.n1190 4.5005
R75965 VDD.n1347 VDD.n1190 4.5005
R75966 VDD.n1337 VDD.n1190 4.5005
R75967 VDD.n1348 VDD.n1190 4.5005
R75968 VDD.n1336 VDD.n1190 4.5005
R75969 VDD.n1350 VDD.n1190 4.5005
R75970 VDD.n1335 VDD.n1190 4.5005
R75971 VDD.n1351 VDD.n1190 4.5005
R75972 VDD.n1334 VDD.n1190 4.5005
R75973 VDD.n1353 VDD.n1190 4.5005
R75974 VDD.n1333 VDD.n1190 4.5005
R75975 VDD.n1354 VDD.n1190 4.5005
R75976 VDD.n1332 VDD.n1190 4.5005
R75977 VDD.n1356 VDD.n1190 4.5005
R75978 VDD.n1331 VDD.n1190 4.5005
R75979 VDD.n1357 VDD.n1190 4.5005
R75980 VDD.n1330 VDD.n1190 4.5005
R75981 VDD.n1359 VDD.n1190 4.5005
R75982 VDD.n1329 VDD.n1190 4.5005
R75983 VDD.n1360 VDD.n1190 4.5005
R75984 VDD.n1328 VDD.n1190 4.5005
R75985 VDD.n1362 VDD.n1190 4.5005
R75986 VDD.n1327 VDD.n1190 4.5005
R75987 VDD.n1363 VDD.n1190 4.5005
R75988 VDD.n1326 VDD.n1190 4.5005
R75989 VDD.n1365 VDD.n1190 4.5005
R75990 VDD.n1325 VDD.n1190 4.5005
R75991 VDD.n1366 VDD.n1190 4.5005
R75992 VDD.n1324 VDD.n1190 4.5005
R75993 VDD.n1368 VDD.n1190 4.5005
R75994 VDD.n1323 VDD.n1190 4.5005
R75995 VDD.n1369 VDD.n1190 4.5005
R75996 VDD.n1322 VDD.n1190 4.5005
R75997 VDD.n1371 VDD.n1190 4.5005
R75998 VDD.n1321 VDD.n1190 4.5005
R75999 VDD.n1372 VDD.n1190 4.5005
R76000 VDD.n1320 VDD.n1190 4.5005
R76001 VDD.n1374 VDD.n1190 4.5005
R76002 VDD.n1319 VDD.n1190 4.5005
R76003 VDD.n1375 VDD.n1190 4.5005
R76004 VDD.n1318 VDD.n1190 4.5005
R76005 VDD.n1376 VDD.n1190 4.5005
R76006 VDD.n1316 VDD.n1190 4.5005
R76007 VDD.n1377 VDD.n1190 4.5005
R76008 VDD.n1315 VDD.n1190 4.5005
R76009 VDD.n1378 VDD.n1190 4.5005
R76010 VDD.n1313 VDD.n1190 4.5005
R76011 VDD.n1379 VDD.n1190 4.5005
R76012 VDD.n1312 VDD.n1190 4.5005
R76013 VDD.n1380 VDD.n1190 4.5005
R76014 VDD.n1310 VDD.n1190 4.5005
R76015 VDD.n1381 VDD.n1190 4.5005
R76016 VDD.n1309 VDD.n1190 4.5005
R76017 VDD.n1382 VDD.n1190 4.5005
R76018 VDD.n1307 VDD.n1190 4.5005
R76019 VDD.n1383 VDD.n1190 4.5005
R76020 VDD.n1306 VDD.n1190 4.5005
R76021 VDD.n1384 VDD.n1190 4.5005
R76022 VDD.n1304 VDD.n1190 4.5005
R76023 VDD.n1385 VDD.n1190 4.5005
R76024 VDD.n1303 VDD.n1190 4.5005
R76025 VDD.n1386 VDD.n1190 4.5005
R76026 VDD.n1301 VDD.n1190 4.5005
R76027 VDD.n1387 VDD.n1190 4.5005
R76028 VDD.n1300 VDD.n1190 4.5005
R76029 VDD.n1388 VDD.n1190 4.5005
R76030 VDD.n1298 VDD.n1190 4.5005
R76031 VDD.n1389 VDD.n1190 4.5005
R76032 VDD.n1297 VDD.n1190 4.5005
R76033 VDD.n1390 VDD.n1190 4.5005
R76034 VDD.n1295 VDD.n1190 4.5005
R76035 VDD.n1391 VDD.n1190 4.5005
R76036 VDD.n1294 VDD.n1190 4.5005
R76037 VDD.n1392 VDD.n1190 4.5005
R76038 VDD.n1292 VDD.n1190 4.5005
R76039 VDD.n1393 VDD.n1190 4.5005
R76040 VDD.n1291 VDD.n1190 4.5005
R76041 VDD.n1394 VDD.n1190 4.5005
R76042 VDD.n1289 VDD.n1190 4.5005
R76043 VDD.n1395 VDD.n1190 4.5005
R76044 VDD.n1288 VDD.n1190 4.5005
R76045 VDD.n1396 VDD.n1190 4.5005
R76046 VDD.n1286 VDD.n1190 4.5005
R76047 VDD.n1397 VDD.n1190 4.5005
R76048 VDD.n1285 VDD.n1190 4.5005
R76049 VDD.n1398 VDD.n1190 4.5005
R76050 VDD.n1283 VDD.n1190 4.5005
R76051 VDD.n1399 VDD.n1190 4.5005
R76052 VDD.n1282 VDD.n1190 4.5005
R76053 VDD.n1400 VDD.n1190 4.5005
R76054 VDD.n1280 VDD.n1190 4.5005
R76055 VDD.n1401 VDD.n1190 4.5005
R76056 VDD.n1279 VDD.n1190 4.5005
R76057 VDD.n1402 VDD.n1190 4.5005
R76058 VDD.n1277 VDD.n1190 4.5005
R76059 VDD.n1403 VDD.n1190 4.5005
R76060 VDD.n1276 VDD.n1190 4.5005
R76061 VDD.n1404 VDD.n1190 4.5005
R76062 VDD.n1274 VDD.n1190 4.5005
R76063 VDD.n1405 VDD.n1190 4.5005
R76064 VDD.n1273 VDD.n1190 4.5005
R76065 VDD.n1406 VDD.n1190 4.5005
R76066 VDD.n1271 VDD.n1190 4.5005
R76067 VDD.n1407 VDD.n1190 4.5005
R76068 VDD.n1270 VDD.n1190 4.5005
R76069 VDD.n1408 VDD.n1190 4.5005
R76070 VDD.n1268 VDD.n1190 4.5005
R76071 VDD.n1409 VDD.n1190 4.5005
R76072 VDD.n1267 VDD.n1190 4.5005
R76073 VDD.n1410 VDD.n1190 4.5005
R76074 VDD.n1265 VDD.n1190 4.5005
R76075 VDD.n1411 VDD.n1190 4.5005
R76076 VDD.n1264 VDD.n1190 4.5005
R76077 VDD.n1412 VDD.n1190 4.5005
R76078 VDD.n1262 VDD.n1190 4.5005
R76079 VDD.n1413 VDD.n1190 4.5005
R76080 VDD.n1261 VDD.n1190 4.5005
R76081 VDD.n1414 VDD.n1190 4.5005
R76082 VDD.n1415 VDD.n1190 4.5005
R76083 VDD.n1674 VDD.n1190 4.5005
R76084 VDD.n1676 VDD.n1200 4.5005
R76085 VDD.n1341 VDD.n1200 4.5005
R76086 VDD.n1342 VDD.n1200 4.5005
R76087 VDD.n1340 VDD.n1200 4.5005
R76088 VDD.n1344 VDD.n1200 4.5005
R76089 VDD.n1339 VDD.n1200 4.5005
R76090 VDD.n1345 VDD.n1200 4.5005
R76091 VDD.n1338 VDD.n1200 4.5005
R76092 VDD.n1347 VDD.n1200 4.5005
R76093 VDD.n1337 VDD.n1200 4.5005
R76094 VDD.n1348 VDD.n1200 4.5005
R76095 VDD.n1336 VDD.n1200 4.5005
R76096 VDD.n1350 VDD.n1200 4.5005
R76097 VDD.n1335 VDD.n1200 4.5005
R76098 VDD.n1351 VDD.n1200 4.5005
R76099 VDD.n1334 VDD.n1200 4.5005
R76100 VDD.n1353 VDD.n1200 4.5005
R76101 VDD.n1333 VDD.n1200 4.5005
R76102 VDD.n1354 VDD.n1200 4.5005
R76103 VDD.n1332 VDD.n1200 4.5005
R76104 VDD.n1356 VDD.n1200 4.5005
R76105 VDD.n1331 VDD.n1200 4.5005
R76106 VDD.n1357 VDD.n1200 4.5005
R76107 VDD.n1330 VDD.n1200 4.5005
R76108 VDD.n1359 VDD.n1200 4.5005
R76109 VDD.n1329 VDD.n1200 4.5005
R76110 VDD.n1360 VDD.n1200 4.5005
R76111 VDD.n1328 VDD.n1200 4.5005
R76112 VDD.n1362 VDD.n1200 4.5005
R76113 VDD.n1327 VDD.n1200 4.5005
R76114 VDD.n1363 VDD.n1200 4.5005
R76115 VDD.n1326 VDD.n1200 4.5005
R76116 VDD.n1365 VDD.n1200 4.5005
R76117 VDD.n1325 VDD.n1200 4.5005
R76118 VDD.n1366 VDD.n1200 4.5005
R76119 VDD.n1324 VDD.n1200 4.5005
R76120 VDD.n1368 VDD.n1200 4.5005
R76121 VDD.n1323 VDD.n1200 4.5005
R76122 VDD.n1369 VDD.n1200 4.5005
R76123 VDD.n1322 VDD.n1200 4.5005
R76124 VDD.n1371 VDD.n1200 4.5005
R76125 VDD.n1321 VDD.n1200 4.5005
R76126 VDD.n1372 VDD.n1200 4.5005
R76127 VDD.n1320 VDD.n1200 4.5005
R76128 VDD.n1374 VDD.n1200 4.5005
R76129 VDD.n1319 VDD.n1200 4.5005
R76130 VDD.n1375 VDD.n1200 4.5005
R76131 VDD.n1318 VDD.n1200 4.5005
R76132 VDD.n1376 VDD.n1200 4.5005
R76133 VDD.n1316 VDD.n1200 4.5005
R76134 VDD.n1377 VDD.n1200 4.5005
R76135 VDD.n1315 VDD.n1200 4.5005
R76136 VDD.n1378 VDD.n1200 4.5005
R76137 VDD.n1313 VDD.n1200 4.5005
R76138 VDD.n1379 VDD.n1200 4.5005
R76139 VDD.n1312 VDD.n1200 4.5005
R76140 VDD.n1380 VDD.n1200 4.5005
R76141 VDD.n1310 VDD.n1200 4.5005
R76142 VDD.n1381 VDD.n1200 4.5005
R76143 VDD.n1309 VDD.n1200 4.5005
R76144 VDD.n1382 VDD.n1200 4.5005
R76145 VDD.n1307 VDD.n1200 4.5005
R76146 VDD.n1383 VDD.n1200 4.5005
R76147 VDD.n1306 VDD.n1200 4.5005
R76148 VDD.n1384 VDD.n1200 4.5005
R76149 VDD.n1304 VDD.n1200 4.5005
R76150 VDD.n1385 VDD.n1200 4.5005
R76151 VDD.n1303 VDD.n1200 4.5005
R76152 VDD.n1386 VDD.n1200 4.5005
R76153 VDD.n1301 VDD.n1200 4.5005
R76154 VDD.n1387 VDD.n1200 4.5005
R76155 VDD.n1300 VDD.n1200 4.5005
R76156 VDD.n1388 VDD.n1200 4.5005
R76157 VDD.n1298 VDD.n1200 4.5005
R76158 VDD.n1389 VDD.n1200 4.5005
R76159 VDD.n1297 VDD.n1200 4.5005
R76160 VDD.n1390 VDD.n1200 4.5005
R76161 VDD.n1295 VDD.n1200 4.5005
R76162 VDD.n1391 VDD.n1200 4.5005
R76163 VDD.n1294 VDD.n1200 4.5005
R76164 VDD.n1392 VDD.n1200 4.5005
R76165 VDD.n1292 VDD.n1200 4.5005
R76166 VDD.n1393 VDD.n1200 4.5005
R76167 VDD.n1291 VDD.n1200 4.5005
R76168 VDD.n1394 VDD.n1200 4.5005
R76169 VDD.n1289 VDD.n1200 4.5005
R76170 VDD.n1395 VDD.n1200 4.5005
R76171 VDD.n1288 VDD.n1200 4.5005
R76172 VDD.n1396 VDD.n1200 4.5005
R76173 VDD.n1286 VDD.n1200 4.5005
R76174 VDD.n1397 VDD.n1200 4.5005
R76175 VDD.n1285 VDD.n1200 4.5005
R76176 VDD.n1398 VDD.n1200 4.5005
R76177 VDD.n1283 VDD.n1200 4.5005
R76178 VDD.n1399 VDD.n1200 4.5005
R76179 VDD.n1282 VDD.n1200 4.5005
R76180 VDD.n1400 VDD.n1200 4.5005
R76181 VDD.n1280 VDD.n1200 4.5005
R76182 VDD.n1401 VDD.n1200 4.5005
R76183 VDD.n1279 VDD.n1200 4.5005
R76184 VDD.n1402 VDD.n1200 4.5005
R76185 VDD.n1277 VDD.n1200 4.5005
R76186 VDD.n1403 VDD.n1200 4.5005
R76187 VDD.n1276 VDD.n1200 4.5005
R76188 VDD.n1404 VDD.n1200 4.5005
R76189 VDD.n1274 VDD.n1200 4.5005
R76190 VDD.n1405 VDD.n1200 4.5005
R76191 VDD.n1273 VDD.n1200 4.5005
R76192 VDD.n1406 VDD.n1200 4.5005
R76193 VDD.n1271 VDD.n1200 4.5005
R76194 VDD.n1407 VDD.n1200 4.5005
R76195 VDD.n1270 VDD.n1200 4.5005
R76196 VDD.n1408 VDD.n1200 4.5005
R76197 VDD.n1268 VDD.n1200 4.5005
R76198 VDD.n1409 VDD.n1200 4.5005
R76199 VDD.n1267 VDD.n1200 4.5005
R76200 VDD.n1410 VDD.n1200 4.5005
R76201 VDD.n1265 VDD.n1200 4.5005
R76202 VDD.n1411 VDD.n1200 4.5005
R76203 VDD.n1264 VDD.n1200 4.5005
R76204 VDD.n1412 VDD.n1200 4.5005
R76205 VDD.n1262 VDD.n1200 4.5005
R76206 VDD.n1413 VDD.n1200 4.5005
R76207 VDD.n1261 VDD.n1200 4.5005
R76208 VDD.n1414 VDD.n1200 4.5005
R76209 VDD.n1415 VDD.n1200 4.5005
R76210 VDD.n1674 VDD.n1200 4.5005
R76211 VDD.n1676 VDD.n1189 4.5005
R76212 VDD.n1341 VDD.n1189 4.5005
R76213 VDD.n1342 VDD.n1189 4.5005
R76214 VDD.n1340 VDD.n1189 4.5005
R76215 VDD.n1344 VDD.n1189 4.5005
R76216 VDD.n1339 VDD.n1189 4.5005
R76217 VDD.n1345 VDD.n1189 4.5005
R76218 VDD.n1338 VDD.n1189 4.5005
R76219 VDD.n1347 VDD.n1189 4.5005
R76220 VDD.n1337 VDD.n1189 4.5005
R76221 VDD.n1348 VDD.n1189 4.5005
R76222 VDD.n1336 VDD.n1189 4.5005
R76223 VDD.n1350 VDD.n1189 4.5005
R76224 VDD.n1335 VDD.n1189 4.5005
R76225 VDD.n1351 VDD.n1189 4.5005
R76226 VDD.n1334 VDD.n1189 4.5005
R76227 VDD.n1353 VDD.n1189 4.5005
R76228 VDD.n1333 VDD.n1189 4.5005
R76229 VDD.n1354 VDD.n1189 4.5005
R76230 VDD.n1332 VDD.n1189 4.5005
R76231 VDD.n1356 VDD.n1189 4.5005
R76232 VDD.n1331 VDD.n1189 4.5005
R76233 VDD.n1357 VDD.n1189 4.5005
R76234 VDD.n1330 VDD.n1189 4.5005
R76235 VDD.n1359 VDD.n1189 4.5005
R76236 VDD.n1329 VDD.n1189 4.5005
R76237 VDD.n1360 VDD.n1189 4.5005
R76238 VDD.n1328 VDD.n1189 4.5005
R76239 VDD.n1362 VDD.n1189 4.5005
R76240 VDD.n1327 VDD.n1189 4.5005
R76241 VDD.n1363 VDD.n1189 4.5005
R76242 VDD.n1326 VDD.n1189 4.5005
R76243 VDD.n1365 VDD.n1189 4.5005
R76244 VDD.n1325 VDD.n1189 4.5005
R76245 VDD.n1366 VDD.n1189 4.5005
R76246 VDD.n1324 VDD.n1189 4.5005
R76247 VDD.n1368 VDD.n1189 4.5005
R76248 VDD.n1323 VDD.n1189 4.5005
R76249 VDD.n1369 VDD.n1189 4.5005
R76250 VDD.n1322 VDD.n1189 4.5005
R76251 VDD.n1371 VDD.n1189 4.5005
R76252 VDD.n1321 VDD.n1189 4.5005
R76253 VDD.n1372 VDD.n1189 4.5005
R76254 VDD.n1320 VDD.n1189 4.5005
R76255 VDD.n1374 VDD.n1189 4.5005
R76256 VDD.n1319 VDD.n1189 4.5005
R76257 VDD.n1375 VDD.n1189 4.5005
R76258 VDD.n1318 VDD.n1189 4.5005
R76259 VDD.n1376 VDD.n1189 4.5005
R76260 VDD.n1316 VDD.n1189 4.5005
R76261 VDD.n1377 VDD.n1189 4.5005
R76262 VDD.n1315 VDD.n1189 4.5005
R76263 VDD.n1378 VDD.n1189 4.5005
R76264 VDD.n1313 VDD.n1189 4.5005
R76265 VDD.n1379 VDD.n1189 4.5005
R76266 VDD.n1312 VDD.n1189 4.5005
R76267 VDD.n1380 VDD.n1189 4.5005
R76268 VDD.n1310 VDD.n1189 4.5005
R76269 VDD.n1381 VDD.n1189 4.5005
R76270 VDD.n1309 VDD.n1189 4.5005
R76271 VDD.n1382 VDD.n1189 4.5005
R76272 VDD.n1307 VDD.n1189 4.5005
R76273 VDD.n1383 VDD.n1189 4.5005
R76274 VDD.n1306 VDD.n1189 4.5005
R76275 VDD.n1384 VDD.n1189 4.5005
R76276 VDD.n1304 VDD.n1189 4.5005
R76277 VDD.n1385 VDD.n1189 4.5005
R76278 VDD.n1303 VDD.n1189 4.5005
R76279 VDD.n1386 VDD.n1189 4.5005
R76280 VDD.n1301 VDD.n1189 4.5005
R76281 VDD.n1387 VDD.n1189 4.5005
R76282 VDD.n1300 VDD.n1189 4.5005
R76283 VDD.n1388 VDD.n1189 4.5005
R76284 VDD.n1298 VDD.n1189 4.5005
R76285 VDD.n1389 VDD.n1189 4.5005
R76286 VDD.n1297 VDD.n1189 4.5005
R76287 VDD.n1390 VDD.n1189 4.5005
R76288 VDD.n1295 VDD.n1189 4.5005
R76289 VDD.n1391 VDD.n1189 4.5005
R76290 VDD.n1294 VDD.n1189 4.5005
R76291 VDD.n1392 VDD.n1189 4.5005
R76292 VDD.n1292 VDD.n1189 4.5005
R76293 VDD.n1393 VDD.n1189 4.5005
R76294 VDD.n1291 VDD.n1189 4.5005
R76295 VDD.n1394 VDD.n1189 4.5005
R76296 VDD.n1289 VDD.n1189 4.5005
R76297 VDD.n1395 VDD.n1189 4.5005
R76298 VDD.n1288 VDD.n1189 4.5005
R76299 VDD.n1396 VDD.n1189 4.5005
R76300 VDD.n1286 VDD.n1189 4.5005
R76301 VDD.n1397 VDD.n1189 4.5005
R76302 VDD.n1285 VDD.n1189 4.5005
R76303 VDD.n1398 VDD.n1189 4.5005
R76304 VDD.n1283 VDD.n1189 4.5005
R76305 VDD.n1399 VDD.n1189 4.5005
R76306 VDD.n1282 VDD.n1189 4.5005
R76307 VDD.n1400 VDD.n1189 4.5005
R76308 VDD.n1280 VDD.n1189 4.5005
R76309 VDD.n1401 VDD.n1189 4.5005
R76310 VDD.n1279 VDD.n1189 4.5005
R76311 VDD.n1402 VDD.n1189 4.5005
R76312 VDD.n1277 VDD.n1189 4.5005
R76313 VDD.n1403 VDD.n1189 4.5005
R76314 VDD.n1276 VDD.n1189 4.5005
R76315 VDD.n1404 VDD.n1189 4.5005
R76316 VDD.n1274 VDD.n1189 4.5005
R76317 VDD.n1405 VDD.n1189 4.5005
R76318 VDD.n1273 VDD.n1189 4.5005
R76319 VDD.n1406 VDD.n1189 4.5005
R76320 VDD.n1271 VDD.n1189 4.5005
R76321 VDD.n1407 VDD.n1189 4.5005
R76322 VDD.n1270 VDD.n1189 4.5005
R76323 VDD.n1408 VDD.n1189 4.5005
R76324 VDD.n1268 VDD.n1189 4.5005
R76325 VDD.n1409 VDD.n1189 4.5005
R76326 VDD.n1267 VDD.n1189 4.5005
R76327 VDD.n1410 VDD.n1189 4.5005
R76328 VDD.n1265 VDD.n1189 4.5005
R76329 VDD.n1411 VDD.n1189 4.5005
R76330 VDD.n1264 VDD.n1189 4.5005
R76331 VDD.n1412 VDD.n1189 4.5005
R76332 VDD.n1262 VDD.n1189 4.5005
R76333 VDD.n1413 VDD.n1189 4.5005
R76334 VDD.n1261 VDD.n1189 4.5005
R76335 VDD.n1414 VDD.n1189 4.5005
R76336 VDD.n1415 VDD.n1189 4.5005
R76337 VDD.n1674 VDD.n1189 4.5005
R76338 VDD.n1676 VDD.n1201 4.5005
R76339 VDD.n1341 VDD.n1201 4.5005
R76340 VDD.n1342 VDD.n1201 4.5005
R76341 VDD.n1340 VDD.n1201 4.5005
R76342 VDD.n1344 VDD.n1201 4.5005
R76343 VDD.n1339 VDD.n1201 4.5005
R76344 VDD.n1345 VDD.n1201 4.5005
R76345 VDD.n1338 VDD.n1201 4.5005
R76346 VDD.n1347 VDD.n1201 4.5005
R76347 VDD.n1337 VDD.n1201 4.5005
R76348 VDD.n1348 VDD.n1201 4.5005
R76349 VDD.n1336 VDD.n1201 4.5005
R76350 VDD.n1350 VDD.n1201 4.5005
R76351 VDD.n1335 VDD.n1201 4.5005
R76352 VDD.n1351 VDD.n1201 4.5005
R76353 VDD.n1334 VDD.n1201 4.5005
R76354 VDD.n1353 VDD.n1201 4.5005
R76355 VDD.n1333 VDD.n1201 4.5005
R76356 VDD.n1354 VDD.n1201 4.5005
R76357 VDD.n1332 VDD.n1201 4.5005
R76358 VDD.n1356 VDD.n1201 4.5005
R76359 VDD.n1331 VDD.n1201 4.5005
R76360 VDD.n1357 VDD.n1201 4.5005
R76361 VDD.n1330 VDD.n1201 4.5005
R76362 VDD.n1359 VDD.n1201 4.5005
R76363 VDD.n1329 VDD.n1201 4.5005
R76364 VDD.n1360 VDD.n1201 4.5005
R76365 VDD.n1328 VDD.n1201 4.5005
R76366 VDD.n1362 VDD.n1201 4.5005
R76367 VDD.n1327 VDD.n1201 4.5005
R76368 VDD.n1363 VDD.n1201 4.5005
R76369 VDD.n1326 VDD.n1201 4.5005
R76370 VDD.n1365 VDD.n1201 4.5005
R76371 VDD.n1325 VDD.n1201 4.5005
R76372 VDD.n1366 VDD.n1201 4.5005
R76373 VDD.n1324 VDD.n1201 4.5005
R76374 VDD.n1368 VDD.n1201 4.5005
R76375 VDD.n1323 VDD.n1201 4.5005
R76376 VDD.n1369 VDD.n1201 4.5005
R76377 VDD.n1322 VDD.n1201 4.5005
R76378 VDD.n1371 VDD.n1201 4.5005
R76379 VDD.n1321 VDD.n1201 4.5005
R76380 VDD.n1372 VDD.n1201 4.5005
R76381 VDD.n1320 VDD.n1201 4.5005
R76382 VDD.n1374 VDD.n1201 4.5005
R76383 VDD.n1319 VDD.n1201 4.5005
R76384 VDD.n1375 VDD.n1201 4.5005
R76385 VDD.n1318 VDD.n1201 4.5005
R76386 VDD.n1376 VDD.n1201 4.5005
R76387 VDD.n1316 VDD.n1201 4.5005
R76388 VDD.n1377 VDD.n1201 4.5005
R76389 VDD.n1315 VDD.n1201 4.5005
R76390 VDD.n1378 VDD.n1201 4.5005
R76391 VDD.n1313 VDD.n1201 4.5005
R76392 VDD.n1379 VDD.n1201 4.5005
R76393 VDD.n1312 VDD.n1201 4.5005
R76394 VDD.n1380 VDD.n1201 4.5005
R76395 VDD.n1310 VDD.n1201 4.5005
R76396 VDD.n1381 VDD.n1201 4.5005
R76397 VDD.n1309 VDD.n1201 4.5005
R76398 VDD.n1382 VDD.n1201 4.5005
R76399 VDD.n1307 VDD.n1201 4.5005
R76400 VDD.n1383 VDD.n1201 4.5005
R76401 VDD.n1306 VDD.n1201 4.5005
R76402 VDD.n1384 VDD.n1201 4.5005
R76403 VDD.n1304 VDD.n1201 4.5005
R76404 VDD.n1385 VDD.n1201 4.5005
R76405 VDD.n1303 VDD.n1201 4.5005
R76406 VDD.n1386 VDD.n1201 4.5005
R76407 VDD.n1301 VDD.n1201 4.5005
R76408 VDD.n1387 VDD.n1201 4.5005
R76409 VDD.n1300 VDD.n1201 4.5005
R76410 VDD.n1388 VDD.n1201 4.5005
R76411 VDD.n1298 VDD.n1201 4.5005
R76412 VDD.n1389 VDD.n1201 4.5005
R76413 VDD.n1297 VDD.n1201 4.5005
R76414 VDD.n1390 VDD.n1201 4.5005
R76415 VDD.n1295 VDD.n1201 4.5005
R76416 VDD.n1391 VDD.n1201 4.5005
R76417 VDD.n1294 VDD.n1201 4.5005
R76418 VDD.n1392 VDD.n1201 4.5005
R76419 VDD.n1292 VDD.n1201 4.5005
R76420 VDD.n1393 VDD.n1201 4.5005
R76421 VDD.n1291 VDD.n1201 4.5005
R76422 VDD.n1394 VDD.n1201 4.5005
R76423 VDD.n1289 VDD.n1201 4.5005
R76424 VDD.n1395 VDD.n1201 4.5005
R76425 VDD.n1288 VDD.n1201 4.5005
R76426 VDD.n1396 VDD.n1201 4.5005
R76427 VDD.n1286 VDD.n1201 4.5005
R76428 VDD.n1397 VDD.n1201 4.5005
R76429 VDD.n1285 VDD.n1201 4.5005
R76430 VDD.n1398 VDD.n1201 4.5005
R76431 VDD.n1283 VDD.n1201 4.5005
R76432 VDD.n1399 VDD.n1201 4.5005
R76433 VDD.n1282 VDD.n1201 4.5005
R76434 VDD.n1400 VDD.n1201 4.5005
R76435 VDD.n1280 VDD.n1201 4.5005
R76436 VDD.n1401 VDD.n1201 4.5005
R76437 VDD.n1279 VDD.n1201 4.5005
R76438 VDD.n1402 VDD.n1201 4.5005
R76439 VDD.n1277 VDD.n1201 4.5005
R76440 VDD.n1403 VDD.n1201 4.5005
R76441 VDD.n1276 VDD.n1201 4.5005
R76442 VDD.n1404 VDD.n1201 4.5005
R76443 VDD.n1274 VDD.n1201 4.5005
R76444 VDD.n1405 VDD.n1201 4.5005
R76445 VDD.n1273 VDD.n1201 4.5005
R76446 VDD.n1406 VDD.n1201 4.5005
R76447 VDD.n1271 VDD.n1201 4.5005
R76448 VDD.n1407 VDD.n1201 4.5005
R76449 VDD.n1270 VDD.n1201 4.5005
R76450 VDD.n1408 VDD.n1201 4.5005
R76451 VDD.n1268 VDD.n1201 4.5005
R76452 VDD.n1409 VDD.n1201 4.5005
R76453 VDD.n1267 VDD.n1201 4.5005
R76454 VDD.n1410 VDD.n1201 4.5005
R76455 VDD.n1265 VDD.n1201 4.5005
R76456 VDD.n1411 VDD.n1201 4.5005
R76457 VDD.n1264 VDD.n1201 4.5005
R76458 VDD.n1412 VDD.n1201 4.5005
R76459 VDD.n1262 VDD.n1201 4.5005
R76460 VDD.n1413 VDD.n1201 4.5005
R76461 VDD.n1261 VDD.n1201 4.5005
R76462 VDD.n1414 VDD.n1201 4.5005
R76463 VDD.n1415 VDD.n1201 4.5005
R76464 VDD.n1674 VDD.n1201 4.5005
R76465 VDD.n1676 VDD.n1188 4.5005
R76466 VDD.n1341 VDD.n1188 4.5005
R76467 VDD.n1342 VDD.n1188 4.5005
R76468 VDD.n1340 VDD.n1188 4.5005
R76469 VDD.n1344 VDD.n1188 4.5005
R76470 VDD.n1339 VDD.n1188 4.5005
R76471 VDD.n1345 VDD.n1188 4.5005
R76472 VDD.n1338 VDD.n1188 4.5005
R76473 VDD.n1347 VDD.n1188 4.5005
R76474 VDD.n1337 VDD.n1188 4.5005
R76475 VDD.n1348 VDD.n1188 4.5005
R76476 VDD.n1336 VDD.n1188 4.5005
R76477 VDD.n1350 VDD.n1188 4.5005
R76478 VDD.n1335 VDD.n1188 4.5005
R76479 VDD.n1351 VDD.n1188 4.5005
R76480 VDD.n1334 VDD.n1188 4.5005
R76481 VDD.n1353 VDD.n1188 4.5005
R76482 VDD.n1333 VDD.n1188 4.5005
R76483 VDD.n1354 VDD.n1188 4.5005
R76484 VDD.n1332 VDD.n1188 4.5005
R76485 VDD.n1356 VDD.n1188 4.5005
R76486 VDD.n1331 VDD.n1188 4.5005
R76487 VDD.n1357 VDD.n1188 4.5005
R76488 VDD.n1330 VDD.n1188 4.5005
R76489 VDD.n1359 VDD.n1188 4.5005
R76490 VDD.n1329 VDD.n1188 4.5005
R76491 VDD.n1360 VDD.n1188 4.5005
R76492 VDD.n1328 VDD.n1188 4.5005
R76493 VDD.n1362 VDD.n1188 4.5005
R76494 VDD.n1327 VDD.n1188 4.5005
R76495 VDD.n1363 VDD.n1188 4.5005
R76496 VDD.n1326 VDD.n1188 4.5005
R76497 VDD.n1365 VDD.n1188 4.5005
R76498 VDD.n1325 VDD.n1188 4.5005
R76499 VDD.n1366 VDD.n1188 4.5005
R76500 VDD.n1324 VDD.n1188 4.5005
R76501 VDD.n1368 VDD.n1188 4.5005
R76502 VDD.n1323 VDD.n1188 4.5005
R76503 VDD.n1369 VDD.n1188 4.5005
R76504 VDD.n1322 VDD.n1188 4.5005
R76505 VDD.n1371 VDD.n1188 4.5005
R76506 VDD.n1321 VDD.n1188 4.5005
R76507 VDD.n1372 VDD.n1188 4.5005
R76508 VDD.n1320 VDD.n1188 4.5005
R76509 VDD.n1374 VDD.n1188 4.5005
R76510 VDD.n1319 VDD.n1188 4.5005
R76511 VDD.n1375 VDD.n1188 4.5005
R76512 VDD.n1318 VDD.n1188 4.5005
R76513 VDD.n1376 VDD.n1188 4.5005
R76514 VDD.n1316 VDD.n1188 4.5005
R76515 VDD.n1377 VDD.n1188 4.5005
R76516 VDD.n1315 VDD.n1188 4.5005
R76517 VDD.n1378 VDD.n1188 4.5005
R76518 VDD.n1313 VDD.n1188 4.5005
R76519 VDD.n1379 VDD.n1188 4.5005
R76520 VDD.n1312 VDD.n1188 4.5005
R76521 VDD.n1380 VDD.n1188 4.5005
R76522 VDD.n1310 VDD.n1188 4.5005
R76523 VDD.n1381 VDD.n1188 4.5005
R76524 VDD.n1309 VDD.n1188 4.5005
R76525 VDD.n1382 VDD.n1188 4.5005
R76526 VDD.n1307 VDD.n1188 4.5005
R76527 VDD.n1383 VDD.n1188 4.5005
R76528 VDD.n1306 VDD.n1188 4.5005
R76529 VDD.n1384 VDD.n1188 4.5005
R76530 VDD.n1304 VDD.n1188 4.5005
R76531 VDD.n1385 VDD.n1188 4.5005
R76532 VDD.n1303 VDD.n1188 4.5005
R76533 VDD.n1386 VDD.n1188 4.5005
R76534 VDD.n1301 VDD.n1188 4.5005
R76535 VDD.n1387 VDD.n1188 4.5005
R76536 VDD.n1300 VDD.n1188 4.5005
R76537 VDD.n1388 VDD.n1188 4.5005
R76538 VDD.n1298 VDD.n1188 4.5005
R76539 VDD.n1389 VDD.n1188 4.5005
R76540 VDD.n1297 VDD.n1188 4.5005
R76541 VDD.n1390 VDD.n1188 4.5005
R76542 VDD.n1295 VDD.n1188 4.5005
R76543 VDD.n1391 VDD.n1188 4.5005
R76544 VDD.n1294 VDD.n1188 4.5005
R76545 VDD.n1392 VDD.n1188 4.5005
R76546 VDD.n1292 VDD.n1188 4.5005
R76547 VDD.n1393 VDD.n1188 4.5005
R76548 VDD.n1291 VDD.n1188 4.5005
R76549 VDD.n1394 VDD.n1188 4.5005
R76550 VDD.n1289 VDD.n1188 4.5005
R76551 VDD.n1395 VDD.n1188 4.5005
R76552 VDD.n1288 VDD.n1188 4.5005
R76553 VDD.n1396 VDD.n1188 4.5005
R76554 VDD.n1286 VDD.n1188 4.5005
R76555 VDD.n1397 VDD.n1188 4.5005
R76556 VDD.n1285 VDD.n1188 4.5005
R76557 VDD.n1398 VDD.n1188 4.5005
R76558 VDD.n1283 VDD.n1188 4.5005
R76559 VDD.n1399 VDD.n1188 4.5005
R76560 VDD.n1282 VDD.n1188 4.5005
R76561 VDD.n1400 VDD.n1188 4.5005
R76562 VDD.n1280 VDD.n1188 4.5005
R76563 VDD.n1401 VDD.n1188 4.5005
R76564 VDD.n1279 VDD.n1188 4.5005
R76565 VDD.n1402 VDD.n1188 4.5005
R76566 VDD.n1277 VDD.n1188 4.5005
R76567 VDD.n1403 VDD.n1188 4.5005
R76568 VDD.n1276 VDD.n1188 4.5005
R76569 VDD.n1404 VDD.n1188 4.5005
R76570 VDD.n1274 VDD.n1188 4.5005
R76571 VDD.n1405 VDD.n1188 4.5005
R76572 VDD.n1273 VDD.n1188 4.5005
R76573 VDD.n1406 VDD.n1188 4.5005
R76574 VDD.n1271 VDD.n1188 4.5005
R76575 VDD.n1407 VDD.n1188 4.5005
R76576 VDD.n1270 VDD.n1188 4.5005
R76577 VDD.n1408 VDD.n1188 4.5005
R76578 VDD.n1268 VDD.n1188 4.5005
R76579 VDD.n1409 VDD.n1188 4.5005
R76580 VDD.n1267 VDD.n1188 4.5005
R76581 VDD.n1410 VDD.n1188 4.5005
R76582 VDD.n1265 VDD.n1188 4.5005
R76583 VDD.n1411 VDD.n1188 4.5005
R76584 VDD.n1264 VDD.n1188 4.5005
R76585 VDD.n1412 VDD.n1188 4.5005
R76586 VDD.n1262 VDD.n1188 4.5005
R76587 VDD.n1413 VDD.n1188 4.5005
R76588 VDD.n1261 VDD.n1188 4.5005
R76589 VDD.n1414 VDD.n1188 4.5005
R76590 VDD.n1415 VDD.n1188 4.5005
R76591 VDD.n1674 VDD.n1188 4.5005
R76592 VDD.n1676 VDD.n1202 4.5005
R76593 VDD.n1341 VDD.n1202 4.5005
R76594 VDD.n1342 VDD.n1202 4.5005
R76595 VDD.n1340 VDD.n1202 4.5005
R76596 VDD.n1344 VDD.n1202 4.5005
R76597 VDD.n1339 VDD.n1202 4.5005
R76598 VDD.n1345 VDD.n1202 4.5005
R76599 VDD.n1338 VDD.n1202 4.5005
R76600 VDD.n1347 VDD.n1202 4.5005
R76601 VDD.n1337 VDD.n1202 4.5005
R76602 VDD.n1348 VDD.n1202 4.5005
R76603 VDD.n1336 VDD.n1202 4.5005
R76604 VDD.n1350 VDD.n1202 4.5005
R76605 VDD.n1335 VDD.n1202 4.5005
R76606 VDD.n1351 VDD.n1202 4.5005
R76607 VDD.n1334 VDD.n1202 4.5005
R76608 VDD.n1353 VDD.n1202 4.5005
R76609 VDD.n1333 VDD.n1202 4.5005
R76610 VDD.n1354 VDD.n1202 4.5005
R76611 VDD.n1332 VDD.n1202 4.5005
R76612 VDD.n1356 VDD.n1202 4.5005
R76613 VDD.n1331 VDD.n1202 4.5005
R76614 VDD.n1357 VDD.n1202 4.5005
R76615 VDD.n1330 VDD.n1202 4.5005
R76616 VDD.n1359 VDD.n1202 4.5005
R76617 VDD.n1329 VDD.n1202 4.5005
R76618 VDD.n1360 VDD.n1202 4.5005
R76619 VDD.n1328 VDD.n1202 4.5005
R76620 VDD.n1362 VDD.n1202 4.5005
R76621 VDD.n1327 VDD.n1202 4.5005
R76622 VDD.n1363 VDD.n1202 4.5005
R76623 VDD.n1326 VDD.n1202 4.5005
R76624 VDD.n1365 VDD.n1202 4.5005
R76625 VDD.n1325 VDD.n1202 4.5005
R76626 VDD.n1366 VDD.n1202 4.5005
R76627 VDD.n1324 VDD.n1202 4.5005
R76628 VDD.n1368 VDD.n1202 4.5005
R76629 VDD.n1323 VDD.n1202 4.5005
R76630 VDD.n1369 VDD.n1202 4.5005
R76631 VDD.n1322 VDD.n1202 4.5005
R76632 VDD.n1371 VDD.n1202 4.5005
R76633 VDD.n1321 VDD.n1202 4.5005
R76634 VDD.n1372 VDD.n1202 4.5005
R76635 VDD.n1320 VDD.n1202 4.5005
R76636 VDD.n1374 VDD.n1202 4.5005
R76637 VDD.n1319 VDD.n1202 4.5005
R76638 VDD.n1375 VDD.n1202 4.5005
R76639 VDD.n1318 VDD.n1202 4.5005
R76640 VDD.n1376 VDD.n1202 4.5005
R76641 VDD.n1316 VDD.n1202 4.5005
R76642 VDD.n1377 VDD.n1202 4.5005
R76643 VDD.n1315 VDD.n1202 4.5005
R76644 VDD.n1378 VDD.n1202 4.5005
R76645 VDD.n1313 VDD.n1202 4.5005
R76646 VDD.n1379 VDD.n1202 4.5005
R76647 VDD.n1312 VDD.n1202 4.5005
R76648 VDD.n1380 VDD.n1202 4.5005
R76649 VDD.n1310 VDD.n1202 4.5005
R76650 VDD.n1381 VDD.n1202 4.5005
R76651 VDD.n1309 VDD.n1202 4.5005
R76652 VDD.n1382 VDD.n1202 4.5005
R76653 VDD.n1307 VDD.n1202 4.5005
R76654 VDD.n1383 VDD.n1202 4.5005
R76655 VDD.n1306 VDD.n1202 4.5005
R76656 VDD.n1384 VDD.n1202 4.5005
R76657 VDD.n1304 VDD.n1202 4.5005
R76658 VDD.n1385 VDD.n1202 4.5005
R76659 VDD.n1303 VDD.n1202 4.5005
R76660 VDD.n1386 VDD.n1202 4.5005
R76661 VDD.n1301 VDD.n1202 4.5005
R76662 VDD.n1387 VDD.n1202 4.5005
R76663 VDD.n1300 VDD.n1202 4.5005
R76664 VDD.n1388 VDD.n1202 4.5005
R76665 VDD.n1298 VDD.n1202 4.5005
R76666 VDD.n1389 VDD.n1202 4.5005
R76667 VDD.n1297 VDD.n1202 4.5005
R76668 VDD.n1390 VDD.n1202 4.5005
R76669 VDD.n1295 VDD.n1202 4.5005
R76670 VDD.n1391 VDD.n1202 4.5005
R76671 VDD.n1294 VDD.n1202 4.5005
R76672 VDD.n1392 VDD.n1202 4.5005
R76673 VDD.n1292 VDD.n1202 4.5005
R76674 VDD.n1393 VDD.n1202 4.5005
R76675 VDD.n1291 VDD.n1202 4.5005
R76676 VDD.n1394 VDD.n1202 4.5005
R76677 VDD.n1289 VDD.n1202 4.5005
R76678 VDD.n1395 VDD.n1202 4.5005
R76679 VDD.n1288 VDD.n1202 4.5005
R76680 VDD.n1396 VDD.n1202 4.5005
R76681 VDD.n1286 VDD.n1202 4.5005
R76682 VDD.n1397 VDD.n1202 4.5005
R76683 VDD.n1285 VDD.n1202 4.5005
R76684 VDD.n1398 VDD.n1202 4.5005
R76685 VDD.n1283 VDD.n1202 4.5005
R76686 VDD.n1399 VDD.n1202 4.5005
R76687 VDD.n1282 VDD.n1202 4.5005
R76688 VDD.n1400 VDD.n1202 4.5005
R76689 VDD.n1280 VDD.n1202 4.5005
R76690 VDD.n1401 VDD.n1202 4.5005
R76691 VDD.n1279 VDD.n1202 4.5005
R76692 VDD.n1402 VDD.n1202 4.5005
R76693 VDD.n1277 VDD.n1202 4.5005
R76694 VDD.n1403 VDD.n1202 4.5005
R76695 VDD.n1276 VDD.n1202 4.5005
R76696 VDD.n1404 VDD.n1202 4.5005
R76697 VDD.n1274 VDD.n1202 4.5005
R76698 VDD.n1405 VDD.n1202 4.5005
R76699 VDD.n1273 VDD.n1202 4.5005
R76700 VDD.n1406 VDD.n1202 4.5005
R76701 VDD.n1271 VDD.n1202 4.5005
R76702 VDD.n1407 VDD.n1202 4.5005
R76703 VDD.n1270 VDD.n1202 4.5005
R76704 VDD.n1408 VDD.n1202 4.5005
R76705 VDD.n1268 VDD.n1202 4.5005
R76706 VDD.n1409 VDD.n1202 4.5005
R76707 VDD.n1267 VDD.n1202 4.5005
R76708 VDD.n1410 VDD.n1202 4.5005
R76709 VDD.n1265 VDD.n1202 4.5005
R76710 VDD.n1411 VDD.n1202 4.5005
R76711 VDD.n1264 VDD.n1202 4.5005
R76712 VDD.n1412 VDD.n1202 4.5005
R76713 VDD.n1262 VDD.n1202 4.5005
R76714 VDD.n1413 VDD.n1202 4.5005
R76715 VDD.n1261 VDD.n1202 4.5005
R76716 VDD.n1414 VDD.n1202 4.5005
R76717 VDD.n1415 VDD.n1202 4.5005
R76718 VDD.n1674 VDD.n1202 4.5005
R76719 VDD.n1676 VDD.n1187 4.5005
R76720 VDD.n1341 VDD.n1187 4.5005
R76721 VDD.n1342 VDD.n1187 4.5005
R76722 VDD.n1340 VDD.n1187 4.5005
R76723 VDD.n1344 VDD.n1187 4.5005
R76724 VDD.n1339 VDD.n1187 4.5005
R76725 VDD.n1345 VDD.n1187 4.5005
R76726 VDD.n1338 VDD.n1187 4.5005
R76727 VDD.n1347 VDD.n1187 4.5005
R76728 VDD.n1337 VDD.n1187 4.5005
R76729 VDD.n1348 VDD.n1187 4.5005
R76730 VDD.n1336 VDD.n1187 4.5005
R76731 VDD.n1350 VDD.n1187 4.5005
R76732 VDD.n1335 VDD.n1187 4.5005
R76733 VDD.n1351 VDD.n1187 4.5005
R76734 VDD.n1334 VDD.n1187 4.5005
R76735 VDD.n1353 VDD.n1187 4.5005
R76736 VDD.n1333 VDD.n1187 4.5005
R76737 VDD.n1354 VDD.n1187 4.5005
R76738 VDD.n1332 VDD.n1187 4.5005
R76739 VDD.n1356 VDD.n1187 4.5005
R76740 VDD.n1331 VDD.n1187 4.5005
R76741 VDD.n1357 VDD.n1187 4.5005
R76742 VDD.n1330 VDD.n1187 4.5005
R76743 VDD.n1359 VDD.n1187 4.5005
R76744 VDD.n1329 VDD.n1187 4.5005
R76745 VDD.n1360 VDD.n1187 4.5005
R76746 VDD.n1328 VDD.n1187 4.5005
R76747 VDD.n1362 VDD.n1187 4.5005
R76748 VDD.n1327 VDD.n1187 4.5005
R76749 VDD.n1363 VDD.n1187 4.5005
R76750 VDD.n1326 VDD.n1187 4.5005
R76751 VDD.n1365 VDD.n1187 4.5005
R76752 VDD.n1325 VDD.n1187 4.5005
R76753 VDD.n1366 VDD.n1187 4.5005
R76754 VDD.n1324 VDD.n1187 4.5005
R76755 VDD.n1368 VDD.n1187 4.5005
R76756 VDD.n1323 VDD.n1187 4.5005
R76757 VDD.n1369 VDD.n1187 4.5005
R76758 VDD.n1322 VDD.n1187 4.5005
R76759 VDD.n1371 VDD.n1187 4.5005
R76760 VDD.n1321 VDD.n1187 4.5005
R76761 VDD.n1372 VDD.n1187 4.5005
R76762 VDD.n1320 VDD.n1187 4.5005
R76763 VDD.n1374 VDD.n1187 4.5005
R76764 VDD.n1319 VDD.n1187 4.5005
R76765 VDD.n1375 VDD.n1187 4.5005
R76766 VDD.n1318 VDD.n1187 4.5005
R76767 VDD.n1376 VDD.n1187 4.5005
R76768 VDD.n1316 VDD.n1187 4.5005
R76769 VDD.n1377 VDD.n1187 4.5005
R76770 VDD.n1315 VDD.n1187 4.5005
R76771 VDD.n1378 VDD.n1187 4.5005
R76772 VDD.n1313 VDD.n1187 4.5005
R76773 VDD.n1379 VDD.n1187 4.5005
R76774 VDD.n1312 VDD.n1187 4.5005
R76775 VDD.n1380 VDD.n1187 4.5005
R76776 VDD.n1310 VDD.n1187 4.5005
R76777 VDD.n1381 VDD.n1187 4.5005
R76778 VDD.n1309 VDD.n1187 4.5005
R76779 VDD.n1382 VDD.n1187 4.5005
R76780 VDD.n1307 VDD.n1187 4.5005
R76781 VDD.n1383 VDD.n1187 4.5005
R76782 VDD.n1306 VDD.n1187 4.5005
R76783 VDD.n1384 VDD.n1187 4.5005
R76784 VDD.n1304 VDD.n1187 4.5005
R76785 VDD.n1385 VDD.n1187 4.5005
R76786 VDD.n1303 VDD.n1187 4.5005
R76787 VDD.n1386 VDD.n1187 4.5005
R76788 VDD.n1301 VDD.n1187 4.5005
R76789 VDD.n1387 VDD.n1187 4.5005
R76790 VDD.n1300 VDD.n1187 4.5005
R76791 VDD.n1388 VDD.n1187 4.5005
R76792 VDD.n1298 VDD.n1187 4.5005
R76793 VDD.n1389 VDD.n1187 4.5005
R76794 VDD.n1297 VDD.n1187 4.5005
R76795 VDD.n1390 VDD.n1187 4.5005
R76796 VDD.n1295 VDD.n1187 4.5005
R76797 VDD.n1391 VDD.n1187 4.5005
R76798 VDD.n1294 VDD.n1187 4.5005
R76799 VDD.n1392 VDD.n1187 4.5005
R76800 VDD.n1292 VDD.n1187 4.5005
R76801 VDD.n1393 VDD.n1187 4.5005
R76802 VDD.n1291 VDD.n1187 4.5005
R76803 VDD.n1394 VDD.n1187 4.5005
R76804 VDD.n1289 VDD.n1187 4.5005
R76805 VDD.n1395 VDD.n1187 4.5005
R76806 VDD.n1288 VDD.n1187 4.5005
R76807 VDD.n1396 VDD.n1187 4.5005
R76808 VDD.n1286 VDD.n1187 4.5005
R76809 VDD.n1397 VDD.n1187 4.5005
R76810 VDD.n1285 VDD.n1187 4.5005
R76811 VDD.n1398 VDD.n1187 4.5005
R76812 VDD.n1283 VDD.n1187 4.5005
R76813 VDD.n1399 VDD.n1187 4.5005
R76814 VDD.n1282 VDD.n1187 4.5005
R76815 VDD.n1400 VDD.n1187 4.5005
R76816 VDD.n1280 VDD.n1187 4.5005
R76817 VDD.n1401 VDD.n1187 4.5005
R76818 VDD.n1279 VDD.n1187 4.5005
R76819 VDD.n1402 VDD.n1187 4.5005
R76820 VDD.n1277 VDD.n1187 4.5005
R76821 VDD.n1403 VDD.n1187 4.5005
R76822 VDD.n1276 VDD.n1187 4.5005
R76823 VDD.n1404 VDD.n1187 4.5005
R76824 VDD.n1274 VDD.n1187 4.5005
R76825 VDD.n1405 VDD.n1187 4.5005
R76826 VDD.n1273 VDD.n1187 4.5005
R76827 VDD.n1406 VDD.n1187 4.5005
R76828 VDD.n1271 VDD.n1187 4.5005
R76829 VDD.n1407 VDD.n1187 4.5005
R76830 VDD.n1270 VDD.n1187 4.5005
R76831 VDD.n1408 VDD.n1187 4.5005
R76832 VDD.n1268 VDD.n1187 4.5005
R76833 VDD.n1409 VDD.n1187 4.5005
R76834 VDD.n1267 VDD.n1187 4.5005
R76835 VDD.n1410 VDD.n1187 4.5005
R76836 VDD.n1265 VDD.n1187 4.5005
R76837 VDD.n1411 VDD.n1187 4.5005
R76838 VDD.n1264 VDD.n1187 4.5005
R76839 VDD.n1412 VDD.n1187 4.5005
R76840 VDD.n1262 VDD.n1187 4.5005
R76841 VDD.n1413 VDD.n1187 4.5005
R76842 VDD.n1261 VDD.n1187 4.5005
R76843 VDD.n1414 VDD.n1187 4.5005
R76844 VDD.n1415 VDD.n1187 4.5005
R76845 VDD.n1674 VDD.n1187 4.5005
R76846 VDD.n1676 VDD.n1203 4.5005
R76847 VDD.n1341 VDD.n1203 4.5005
R76848 VDD.n1342 VDD.n1203 4.5005
R76849 VDD.n1340 VDD.n1203 4.5005
R76850 VDD.n1344 VDD.n1203 4.5005
R76851 VDD.n1339 VDD.n1203 4.5005
R76852 VDD.n1345 VDD.n1203 4.5005
R76853 VDD.n1338 VDD.n1203 4.5005
R76854 VDD.n1347 VDD.n1203 4.5005
R76855 VDD.n1337 VDD.n1203 4.5005
R76856 VDD.n1348 VDD.n1203 4.5005
R76857 VDD.n1336 VDD.n1203 4.5005
R76858 VDD.n1350 VDD.n1203 4.5005
R76859 VDD.n1335 VDD.n1203 4.5005
R76860 VDD.n1351 VDD.n1203 4.5005
R76861 VDD.n1334 VDD.n1203 4.5005
R76862 VDD.n1353 VDD.n1203 4.5005
R76863 VDD.n1333 VDD.n1203 4.5005
R76864 VDD.n1354 VDD.n1203 4.5005
R76865 VDD.n1332 VDD.n1203 4.5005
R76866 VDD.n1356 VDD.n1203 4.5005
R76867 VDD.n1331 VDD.n1203 4.5005
R76868 VDD.n1357 VDD.n1203 4.5005
R76869 VDD.n1330 VDD.n1203 4.5005
R76870 VDD.n1359 VDD.n1203 4.5005
R76871 VDD.n1329 VDD.n1203 4.5005
R76872 VDD.n1360 VDD.n1203 4.5005
R76873 VDD.n1328 VDD.n1203 4.5005
R76874 VDD.n1362 VDD.n1203 4.5005
R76875 VDD.n1327 VDD.n1203 4.5005
R76876 VDD.n1363 VDD.n1203 4.5005
R76877 VDD.n1326 VDD.n1203 4.5005
R76878 VDD.n1365 VDD.n1203 4.5005
R76879 VDD.n1325 VDD.n1203 4.5005
R76880 VDD.n1366 VDD.n1203 4.5005
R76881 VDD.n1324 VDD.n1203 4.5005
R76882 VDD.n1368 VDD.n1203 4.5005
R76883 VDD.n1323 VDD.n1203 4.5005
R76884 VDD.n1369 VDD.n1203 4.5005
R76885 VDD.n1322 VDD.n1203 4.5005
R76886 VDD.n1371 VDD.n1203 4.5005
R76887 VDD.n1321 VDD.n1203 4.5005
R76888 VDD.n1372 VDD.n1203 4.5005
R76889 VDD.n1320 VDD.n1203 4.5005
R76890 VDD.n1374 VDD.n1203 4.5005
R76891 VDD.n1319 VDD.n1203 4.5005
R76892 VDD.n1375 VDD.n1203 4.5005
R76893 VDD.n1318 VDD.n1203 4.5005
R76894 VDD.n1376 VDD.n1203 4.5005
R76895 VDD.n1316 VDD.n1203 4.5005
R76896 VDD.n1377 VDD.n1203 4.5005
R76897 VDD.n1315 VDD.n1203 4.5005
R76898 VDD.n1378 VDD.n1203 4.5005
R76899 VDD.n1313 VDD.n1203 4.5005
R76900 VDD.n1379 VDD.n1203 4.5005
R76901 VDD.n1312 VDD.n1203 4.5005
R76902 VDD.n1380 VDD.n1203 4.5005
R76903 VDD.n1310 VDD.n1203 4.5005
R76904 VDD.n1381 VDD.n1203 4.5005
R76905 VDD.n1309 VDD.n1203 4.5005
R76906 VDD.n1382 VDD.n1203 4.5005
R76907 VDD.n1307 VDD.n1203 4.5005
R76908 VDD.n1383 VDD.n1203 4.5005
R76909 VDD.n1306 VDD.n1203 4.5005
R76910 VDD.n1384 VDD.n1203 4.5005
R76911 VDD.n1304 VDD.n1203 4.5005
R76912 VDD.n1385 VDD.n1203 4.5005
R76913 VDD.n1303 VDD.n1203 4.5005
R76914 VDD.n1386 VDD.n1203 4.5005
R76915 VDD.n1301 VDD.n1203 4.5005
R76916 VDD.n1387 VDD.n1203 4.5005
R76917 VDD.n1300 VDD.n1203 4.5005
R76918 VDD.n1388 VDD.n1203 4.5005
R76919 VDD.n1298 VDD.n1203 4.5005
R76920 VDD.n1389 VDD.n1203 4.5005
R76921 VDD.n1297 VDD.n1203 4.5005
R76922 VDD.n1390 VDD.n1203 4.5005
R76923 VDD.n1295 VDD.n1203 4.5005
R76924 VDD.n1391 VDD.n1203 4.5005
R76925 VDD.n1294 VDD.n1203 4.5005
R76926 VDD.n1392 VDD.n1203 4.5005
R76927 VDD.n1292 VDD.n1203 4.5005
R76928 VDD.n1393 VDD.n1203 4.5005
R76929 VDD.n1291 VDD.n1203 4.5005
R76930 VDD.n1394 VDD.n1203 4.5005
R76931 VDD.n1289 VDD.n1203 4.5005
R76932 VDD.n1395 VDD.n1203 4.5005
R76933 VDD.n1288 VDD.n1203 4.5005
R76934 VDD.n1396 VDD.n1203 4.5005
R76935 VDD.n1286 VDD.n1203 4.5005
R76936 VDD.n1397 VDD.n1203 4.5005
R76937 VDD.n1285 VDD.n1203 4.5005
R76938 VDD.n1398 VDD.n1203 4.5005
R76939 VDD.n1283 VDD.n1203 4.5005
R76940 VDD.n1399 VDD.n1203 4.5005
R76941 VDD.n1282 VDD.n1203 4.5005
R76942 VDD.n1400 VDD.n1203 4.5005
R76943 VDD.n1280 VDD.n1203 4.5005
R76944 VDD.n1401 VDD.n1203 4.5005
R76945 VDD.n1279 VDD.n1203 4.5005
R76946 VDD.n1402 VDD.n1203 4.5005
R76947 VDD.n1277 VDD.n1203 4.5005
R76948 VDD.n1403 VDD.n1203 4.5005
R76949 VDD.n1276 VDD.n1203 4.5005
R76950 VDD.n1404 VDD.n1203 4.5005
R76951 VDD.n1274 VDD.n1203 4.5005
R76952 VDD.n1405 VDD.n1203 4.5005
R76953 VDD.n1273 VDD.n1203 4.5005
R76954 VDD.n1406 VDD.n1203 4.5005
R76955 VDD.n1271 VDD.n1203 4.5005
R76956 VDD.n1407 VDD.n1203 4.5005
R76957 VDD.n1270 VDD.n1203 4.5005
R76958 VDD.n1408 VDD.n1203 4.5005
R76959 VDD.n1268 VDD.n1203 4.5005
R76960 VDD.n1409 VDD.n1203 4.5005
R76961 VDD.n1267 VDD.n1203 4.5005
R76962 VDD.n1410 VDD.n1203 4.5005
R76963 VDD.n1265 VDD.n1203 4.5005
R76964 VDD.n1411 VDD.n1203 4.5005
R76965 VDD.n1264 VDD.n1203 4.5005
R76966 VDD.n1412 VDD.n1203 4.5005
R76967 VDD.n1262 VDD.n1203 4.5005
R76968 VDD.n1413 VDD.n1203 4.5005
R76969 VDD.n1261 VDD.n1203 4.5005
R76970 VDD.n1414 VDD.n1203 4.5005
R76971 VDD.n1415 VDD.n1203 4.5005
R76972 VDD.n1674 VDD.n1203 4.5005
R76973 VDD.n1676 VDD.n1186 4.5005
R76974 VDD.n1341 VDD.n1186 4.5005
R76975 VDD.n1342 VDD.n1186 4.5005
R76976 VDD.n1340 VDD.n1186 4.5005
R76977 VDD.n1344 VDD.n1186 4.5005
R76978 VDD.n1339 VDD.n1186 4.5005
R76979 VDD.n1345 VDD.n1186 4.5005
R76980 VDD.n1338 VDD.n1186 4.5005
R76981 VDD.n1347 VDD.n1186 4.5005
R76982 VDD.n1337 VDD.n1186 4.5005
R76983 VDD.n1348 VDD.n1186 4.5005
R76984 VDD.n1336 VDD.n1186 4.5005
R76985 VDD.n1350 VDD.n1186 4.5005
R76986 VDD.n1335 VDD.n1186 4.5005
R76987 VDD.n1351 VDD.n1186 4.5005
R76988 VDD.n1334 VDD.n1186 4.5005
R76989 VDD.n1353 VDD.n1186 4.5005
R76990 VDD.n1333 VDD.n1186 4.5005
R76991 VDD.n1354 VDD.n1186 4.5005
R76992 VDD.n1332 VDD.n1186 4.5005
R76993 VDD.n1356 VDD.n1186 4.5005
R76994 VDD.n1331 VDD.n1186 4.5005
R76995 VDD.n1357 VDD.n1186 4.5005
R76996 VDD.n1330 VDD.n1186 4.5005
R76997 VDD.n1359 VDD.n1186 4.5005
R76998 VDD.n1329 VDD.n1186 4.5005
R76999 VDD.n1360 VDD.n1186 4.5005
R77000 VDD.n1328 VDD.n1186 4.5005
R77001 VDD.n1362 VDD.n1186 4.5005
R77002 VDD.n1327 VDD.n1186 4.5005
R77003 VDD.n1363 VDD.n1186 4.5005
R77004 VDD.n1326 VDD.n1186 4.5005
R77005 VDD.n1365 VDD.n1186 4.5005
R77006 VDD.n1325 VDD.n1186 4.5005
R77007 VDD.n1366 VDD.n1186 4.5005
R77008 VDD.n1324 VDD.n1186 4.5005
R77009 VDD.n1368 VDD.n1186 4.5005
R77010 VDD.n1323 VDD.n1186 4.5005
R77011 VDD.n1369 VDD.n1186 4.5005
R77012 VDD.n1322 VDD.n1186 4.5005
R77013 VDD.n1371 VDD.n1186 4.5005
R77014 VDD.n1321 VDD.n1186 4.5005
R77015 VDD.n1372 VDD.n1186 4.5005
R77016 VDD.n1320 VDD.n1186 4.5005
R77017 VDD.n1374 VDD.n1186 4.5005
R77018 VDD.n1319 VDD.n1186 4.5005
R77019 VDD.n1375 VDD.n1186 4.5005
R77020 VDD.n1318 VDD.n1186 4.5005
R77021 VDD.n1376 VDD.n1186 4.5005
R77022 VDD.n1316 VDD.n1186 4.5005
R77023 VDD.n1377 VDD.n1186 4.5005
R77024 VDD.n1315 VDD.n1186 4.5005
R77025 VDD.n1378 VDD.n1186 4.5005
R77026 VDD.n1313 VDD.n1186 4.5005
R77027 VDD.n1379 VDD.n1186 4.5005
R77028 VDD.n1312 VDD.n1186 4.5005
R77029 VDD.n1380 VDD.n1186 4.5005
R77030 VDD.n1310 VDD.n1186 4.5005
R77031 VDD.n1381 VDD.n1186 4.5005
R77032 VDD.n1309 VDD.n1186 4.5005
R77033 VDD.n1382 VDD.n1186 4.5005
R77034 VDD.n1307 VDD.n1186 4.5005
R77035 VDD.n1383 VDD.n1186 4.5005
R77036 VDD.n1306 VDD.n1186 4.5005
R77037 VDD.n1384 VDD.n1186 4.5005
R77038 VDD.n1304 VDD.n1186 4.5005
R77039 VDD.n1385 VDD.n1186 4.5005
R77040 VDD.n1303 VDD.n1186 4.5005
R77041 VDD.n1386 VDD.n1186 4.5005
R77042 VDD.n1301 VDD.n1186 4.5005
R77043 VDD.n1387 VDD.n1186 4.5005
R77044 VDD.n1300 VDD.n1186 4.5005
R77045 VDD.n1388 VDD.n1186 4.5005
R77046 VDD.n1298 VDD.n1186 4.5005
R77047 VDD.n1389 VDD.n1186 4.5005
R77048 VDD.n1297 VDD.n1186 4.5005
R77049 VDD.n1390 VDD.n1186 4.5005
R77050 VDD.n1295 VDD.n1186 4.5005
R77051 VDD.n1391 VDD.n1186 4.5005
R77052 VDD.n1294 VDD.n1186 4.5005
R77053 VDD.n1392 VDD.n1186 4.5005
R77054 VDD.n1292 VDD.n1186 4.5005
R77055 VDD.n1393 VDD.n1186 4.5005
R77056 VDD.n1291 VDD.n1186 4.5005
R77057 VDD.n1394 VDD.n1186 4.5005
R77058 VDD.n1289 VDD.n1186 4.5005
R77059 VDD.n1395 VDD.n1186 4.5005
R77060 VDD.n1288 VDD.n1186 4.5005
R77061 VDD.n1396 VDD.n1186 4.5005
R77062 VDD.n1286 VDD.n1186 4.5005
R77063 VDD.n1397 VDD.n1186 4.5005
R77064 VDD.n1285 VDD.n1186 4.5005
R77065 VDD.n1398 VDD.n1186 4.5005
R77066 VDD.n1283 VDD.n1186 4.5005
R77067 VDD.n1399 VDD.n1186 4.5005
R77068 VDD.n1282 VDD.n1186 4.5005
R77069 VDD.n1400 VDD.n1186 4.5005
R77070 VDD.n1280 VDD.n1186 4.5005
R77071 VDD.n1401 VDD.n1186 4.5005
R77072 VDD.n1279 VDD.n1186 4.5005
R77073 VDD.n1402 VDD.n1186 4.5005
R77074 VDD.n1277 VDD.n1186 4.5005
R77075 VDD.n1403 VDD.n1186 4.5005
R77076 VDD.n1276 VDD.n1186 4.5005
R77077 VDD.n1404 VDD.n1186 4.5005
R77078 VDD.n1274 VDD.n1186 4.5005
R77079 VDD.n1405 VDD.n1186 4.5005
R77080 VDD.n1273 VDD.n1186 4.5005
R77081 VDD.n1406 VDD.n1186 4.5005
R77082 VDD.n1271 VDD.n1186 4.5005
R77083 VDD.n1407 VDD.n1186 4.5005
R77084 VDD.n1270 VDD.n1186 4.5005
R77085 VDD.n1408 VDD.n1186 4.5005
R77086 VDD.n1268 VDD.n1186 4.5005
R77087 VDD.n1409 VDD.n1186 4.5005
R77088 VDD.n1267 VDD.n1186 4.5005
R77089 VDD.n1410 VDD.n1186 4.5005
R77090 VDD.n1265 VDD.n1186 4.5005
R77091 VDD.n1411 VDD.n1186 4.5005
R77092 VDD.n1264 VDD.n1186 4.5005
R77093 VDD.n1412 VDD.n1186 4.5005
R77094 VDD.n1262 VDD.n1186 4.5005
R77095 VDD.n1413 VDD.n1186 4.5005
R77096 VDD.n1261 VDD.n1186 4.5005
R77097 VDD.n1414 VDD.n1186 4.5005
R77098 VDD.n1415 VDD.n1186 4.5005
R77099 VDD.n1674 VDD.n1186 4.5005
R77100 VDD.n1676 VDD.n1204 4.5005
R77101 VDD.n1341 VDD.n1204 4.5005
R77102 VDD.n1342 VDD.n1204 4.5005
R77103 VDD.n1340 VDD.n1204 4.5005
R77104 VDD.n1344 VDD.n1204 4.5005
R77105 VDD.n1339 VDD.n1204 4.5005
R77106 VDD.n1345 VDD.n1204 4.5005
R77107 VDD.n1338 VDD.n1204 4.5005
R77108 VDD.n1347 VDD.n1204 4.5005
R77109 VDD.n1337 VDD.n1204 4.5005
R77110 VDD.n1348 VDD.n1204 4.5005
R77111 VDD.n1336 VDD.n1204 4.5005
R77112 VDD.n1350 VDD.n1204 4.5005
R77113 VDD.n1335 VDD.n1204 4.5005
R77114 VDD.n1351 VDD.n1204 4.5005
R77115 VDD.n1334 VDD.n1204 4.5005
R77116 VDD.n1353 VDD.n1204 4.5005
R77117 VDD.n1333 VDD.n1204 4.5005
R77118 VDD.n1354 VDD.n1204 4.5005
R77119 VDD.n1332 VDD.n1204 4.5005
R77120 VDD.n1356 VDD.n1204 4.5005
R77121 VDD.n1331 VDD.n1204 4.5005
R77122 VDD.n1357 VDD.n1204 4.5005
R77123 VDD.n1330 VDD.n1204 4.5005
R77124 VDD.n1359 VDD.n1204 4.5005
R77125 VDD.n1329 VDD.n1204 4.5005
R77126 VDD.n1360 VDD.n1204 4.5005
R77127 VDD.n1328 VDD.n1204 4.5005
R77128 VDD.n1362 VDD.n1204 4.5005
R77129 VDD.n1327 VDD.n1204 4.5005
R77130 VDD.n1363 VDD.n1204 4.5005
R77131 VDD.n1326 VDD.n1204 4.5005
R77132 VDD.n1365 VDD.n1204 4.5005
R77133 VDD.n1325 VDD.n1204 4.5005
R77134 VDD.n1366 VDD.n1204 4.5005
R77135 VDD.n1324 VDD.n1204 4.5005
R77136 VDD.n1368 VDD.n1204 4.5005
R77137 VDD.n1323 VDD.n1204 4.5005
R77138 VDD.n1369 VDD.n1204 4.5005
R77139 VDD.n1322 VDD.n1204 4.5005
R77140 VDD.n1371 VDD.n1204 4.5005
R77141 VDD.n1321 VDD.n1204 4.5005
R77142 VDD.n1372 VDD.n1204 4.5005
R77143 VDD.n1320 VDD.n1204 4.5005
R77144 VDD.n1374 VDD.n1204 4.5005
R77145 VDD.n1319 VDD.n1204 4.5005
R77146 VDD.n1375 VDD.n1204 4.5005
R77147 VDD.n1318 VDD.n1204 4.5005
R77148 VDD.n1376 VDD.n1204 4.5005
R77149 VDD.n1316 VDD.n1204 4.5005
R77150 VDD.n1377 VDD.n1204 4.5005
R77151 VDD.n1315 VDD.n1204 4.5005
R77152 VDD.n1378 VDD.n1204 4.5005
R77153 VDD.n1313 VDD.n1204 4.5005
R77154 VDD.n1379 VDD.n1204 4.5005
R77155 VDD.n1312 VDD.n1204 4.5005
R77156 VDD.n1380 VDD.n1204 4.5005
R77157 VDD.n1310 VDD.n1204 4.5005
R77158 VDD.n1381 VDD.n1204 4.5005
R77159 VDD.n1309 VDD.n1204 4.5005
R77160 VDD.n1382 VDD.n1204 4.5005
R77161 VDD.n1307 VDD.n1204 4.5005
R77162 VDD.n1383 VDD.n1204 4.5005
R77163 VDD.n1306 VDD.n1204 4.5005
R77164 VDD.n1384 VDD.n1204 4.5005
R77165 VDD.n1304 VDD.n1204 4.5005
R77166 VDD.n1385 VDD.n1204 4.5005
R77167 VDD.n1303 VDD.n1204 4.5005
R77168 VDD.n1386 VDD.n1204 4.5005
R77169 VDD.n1301 VDD.n1204 4.5005
R77170 VDD.n1387 VDD.n1204 4.5005
R77171 VDD.n1300 VDD.n1204 4.5005
R77172 VDD.n1388 VDD.n1204 4.5005
R77173 VDD.n1298 VDD.n1204 4.5005
R77174 VDD.n1389 VDD.n1204 4.5005
R77175 VDD.n1297 VDD.n1204 4.5005
R77176 VDD.n1390 VDD.n1204 4.5005
R77177 VDD.n1295 VDD.n1204 4.5005
R77178 VDD.n1391 VDD.n1204 4.5005
R77179 VDD.n1294 VDD.n1204 4.5005
R77180 VDD.n1392 VDD.n1204 4.5005
R77181 VDD.n1292 VDD.n1204 4.5005
R77182 VDD.n1393 VDD.n1204 4.5005
R77183 VDD.n1291 VDD.n1204 4.5005
R77184 VDD.n1394 VDD.n1204 4.5005
R77185 VDD.n1289 VDD.n1204 4.5005
R77186 VDD.n1395 VDD.n1204 4.5005
R77187 VDD.n1288 VDD.n1204 4.5005
R77188 VDD.n1396 VDD.n1204 4.5005
R77189 VDD.n1286 VDD.n1204 4.5005
R77190 VDD.n1397 VDD.n1204 4.5005
R77191 VDD.n1285 VDD.n1204 4.5005
R77192 VDD.n1398 VDD.n1204 4.5005
R77193 VDD.n1283 VDD.n1204 4.5005
R77194 VDD.n1399 VDD.n1204 4.5005
R77195 VDD.n1282 VDD.n1204 4.5005
R77196 VDD.n1400 VDD.n1204 4.5005
R77197 VDD.n1280 VDD.n1204 4.5005
R77198 VDD.n1401 VDD.n1204 4.5005
R77199 VDD.n1279 VDD.n1204 4.5005
R77200 VDD.n1402 VDD.n1204 4.5005
R77201 VDD.n1277 VDD.n1204 4.5005
R77202 VDD.n1403 VDD.n1204 4.5005
R77203 VDD.n1276 VDD.n1204 4.5005
R77204 VDD.n1404 VDD.n1204 4.5005
R77205 VDD.n1274 VDD.n1204 4.5005
R77206 VDD.n1405 VDD.n1204 4.5005
R77207 VDD.n1273 VDD.n1204 4.5005
R77208 VDD.n1406 VDD.n1204 4.5005
R77209 VDD.n1271 VDD.n1204 4.5005
R77210 VDD.n1407 VDD.n1204 4.5005
R77211 VDD.n1270 VDD.n1204 4.5005
R77212 VDD.n1408 VDD.n1204 4.5005
R77213 VDD.n1268 VDD.n1204 4.5005
R77214 VDD.n1409 VDD.n1204 4.5005
R77215 VDD.n1267 VDD.n1204 4.5005
R77216 VDD.n1410 VDD.n1204 4.5005
R77217 VDD.n1265 VDD.n1204 4.5005
R77218 VDD.n1411 VDD.n1204 4.5005
R77219 VDD.n1264 VDD.n1204 4.5005
R77220 VDD.n1412 VDD.n1204 4.5005
R77221 VDD.n1262 VDD.n1204 4.5005
R77222 VDD.n1413 VDD.n1204 4.5005
R77223 VDD.n1261 VDD.n1204 4.5005
R77224 VDD.n1414 VDD.n1204 4.5005
R77225 VDD.n1415 VDD.n1204 4.5005
R77226 VDD.n1674 VDD.n1204 4.5005
R77227 VDD.n1676 VDD.n1185 4.5005
R77228 VDD.n1341 VDD.n1185 4.5005
R77229 VDD.n1342 VDD.n1185 4.5005
R77230 VDD.n1340 VDD.n1185 4.5005
R77231 VDD.n1344 VDD.n1185 4.5005
R77232 VDD.n1339 VDD.n1185 4.5005
R77233 VDD.n1345 VDD.n1185 4.5005
R77234 VDD.n1338 VDD.n1185 4.5005
R77235 VDD.n1347 VDD.n1185 4.5005
R77236 VDD.n1337 VDD.n1185 4.5005
R77237 VDD.n1348 VDD.n1185 4.5005
R77238 VDD.n1336 VDD.n1185 4.5005
R77239 VDD.n1350 VDD.n1185 4.5005
R77240 VDD.n1335 VDD.n1185 4.5005
R77241 VDD.n1351 VDD.n1185 4.5005
R77242 VDD.n1334 VDD.n1185 4.5005
R77243 VDD.n1353 VDD.n1185 4.5005
R77244 VDD.n1333 VDD.n1185 4.5005
R77245 VDD.n1354 VDD.n1185 4.5005
R77246 VDD.n1332 VDD.n1185 4.5005
R77247 VDD.n1356 VDD.n1185 4.5005
R77248 VDD.n1331 VDD.n1185 4.5005
R77249 VDD.n1357 VDD.n1185 4.5005
R77250 VDD.n1330 VDD.n1185 4.5005
R77251 VDD.n1359 VDD.n1185 4.5005
R77252 VDD.n1329 VDD.n1185 4.5005
R77253 VDD.n1360 VDD.n1185 4.5005
R77254 VDD.n1328 VDD.n1185 4.5005
R77255 VDD.n1362 VDD.n1185 4.5005
R77256 VDD.n1327 VDD.n1185 4.5005
R77257 VDD.n1363 VDD.n1185 4.5005
R77258 VDD.n1326 VDD.n1185 4.5005
R77259 VDD.n1365 VDD.n1185 4.5005
R77260 VDD.n1325 VDD.n1185 4.5005
R77261 VDD.n1366 VDD.n1185 4.5005
R77262 VDD.n1324 VDD.n1185 4.5005
R77263 VDD.n1368 VDD.n1185 4.5005
R77264 VDD.n1323 VDD.n1185 4.5005
R77265 VDD.n1369 VDD.n1185 4.5005
R77266 VDD.n1322 VDD.n1185 4.5005
R77267 VDD.n1371 VDD.n1185 4.5005
R77268 VDD.n1321 VDD.n1185 4.5005
R77269 VDD.n1372 VDD.n1185 4.5005
R77270 VDD.n1320 VDD.n1185 4.5005
R77271 VDD.n1374 VDD.n1185 4.5005
R77272 VDD.n1319 VDD.n1185 4.5005
R77273 VDD.n1375 VDD.n1185 4.5005
R77274 VDD.n1318 VDD.n1185 4.5005
R77275 VDD.n1376 VDD.n1185 4.5005
R77276 VDD.n1316 VDD.n1185 4.5005
R77277 VDD.n1377 VDD.n1185 4.5005
R77278 VDD.n1315 VDD.n1185 4.5005
R77279 VDD.n1378 VDD.n1185 4.5005
R77280 VDD.n1313 VDD.n1185 4.5005
R77281 VDD.n1379 VDD.n1185 4.5005
R77282 VDD.n1312 VDD.n1185 4.5005
R77283 VDD.n1380 VDD.n1185 4.5005
R77284 VDD.n1310 VDD.n1185 4.5005
R77285 VDD.n1381 VDD.n1185 4.5005
R77286 VDD.n1309 VDD.n1185 4.5005
R77287 VDD.n1382 VDD.n1185 4.5005
R77288 VDD.n1307 VDD.n1185 4.5005
R77289 VDD.n1383 VDD.n1185 4.5005
R77290 VDD.n1306 VDD.n1185 4.5005
R77291 VDD.n1384 VDD.n1185 4.5005
R77292 VDD.n1304 VDD.n1185 4.5005
R77293 VDD.n1385 VDD.n1185 4.5005
R77294 VDD.n1303 VDD.n1185 4.5005
R77295 VDD.n1386 VDD.n1185 4.5005
R77296 VDD.n1301 VDD.n1185 4.5005
R77297 VDD.n1387 VDD.n1185 4.5005
R77298 VDD.n1300 VDD.n1185 4.5005
R77299 VDD.n1388 VDD.n1185 4.5005
R77300 VDD.n1298 VDD.n1185 4.5005
R77301 VDD.n1389 VDD.n1185 4.5005
R77302 VDD.n1297 VDD.n1185 4.5005
R77303 VDD.n1390 VDD.n1185 4.5005
R77304 VDD.n1295 VDD.n1185 4.5005
R77305 VDD.n1391 VDD.n1185 4.5005
R77306 VDD.n1294 VDD.n1185 4.5005
R77307 VDD.n1392 VDD.n1185 4.5005
R77308 VDD.n1292 VDD.n1185 4.5005
R77309 VDD.n1393 VDD.n1185 4.5005
R77310 VDD.n1291 VDD.n1185 4.5005
R77311 VDD.n1394 VDD.n1185 4.5005
R77312 VDD.n1289 VDD.n1185 4.5005
R77313 VDD.n1395 VDD.n1185 4.5005
R77314 VDD.n1288 VDD.n1185 4.5005
R77315 VDD.n1396 VDD.n1185 4.5005
R77316 VDD.n1286 VDD.n1185 4.5005
R77317 VDD.n1397 VDD.n1185 4.5005
R77318 VDD.n1285 VDD.n1185 4.5005
R77319 VDD.n1398 VDD.n1185 4.5005
R77320 VDD.n1283 VDD.n1185 4.5005
R77321 VDD.n1399 VDD.n1185 4.5005
R77322 VDD.n1282 VDD.n1185 4.5005
R77323 VDD.n1400 VDD.n1185 4.5005
R77324 VDD.n1280 VDD.n1185 4.5005
R77325 VDD.n1401 VDD.n1185 4.5005
R77326 VDD.n1279 VDD.n1185 4.5005
R77327 VDD.n1402 VDD.n1185 4.5005
R77328 VDD.n1277 VDD.n1185 4.5005
R77329 VDD.n1403 VDD.n1185 4.5005
R77330 VDD.n1276 VDD.n1185 4.5005
R77331 VDD.n1404 VDD.n1185 4.5005
R77332 VDD.n1274 VDD.n1185 4.5005
R77333 VDD.n1405 VDD.n1185 4.5005
R77334 VDD.n1273 VDD.n1185 4.5005
R77335 VDD.n1406 VDD.n1185 4.5005
R77336 VDD.n1271 VDD.n1185 4.5005
R77337 VDD.n1407 VDD.n1185 4.5005
R77338 VDD.n1270 VDD.n1185 4.5005
R77339 VDD.n1408 VDD.n1185 4.5005
R77340 VDD.n1268 VDD.n1185 4.5005
R77341 VDD.n1409 VDD.n1185 4.5005
R77342 VDD.n1267 VDD.n1185 4.5005
R77343 VDD.n1410 VDD.n1185 4.5005
R77344 VDD.n1265 VDD.n1185 4.5005
R77345 VDD.n1411 VDD.n1185 4.5005
R77346 VDD.n1264 VDD.n1185 4.5005
R77347 VDD.n1412 VDD.n1185 4.5005
R77348 VDD.n1262 VDD.n1185 4.5005
R77349 VDD.n1413 VDD.n1185 4.5005
R77350 VDD.n1261 VDD.n1185 4.5005
R77351 VDD.n1414 VDD.n1185 4.5005
R77352 VDD.n1415 VDD.n1185 4.5005
R77353 VDD.n1674 VDD.n1185 4.5005
R77354 VDD.n1676 VDD.n1205 4.5005
R77355 VDD.n1341 VDD.n1205 4.5005
R77356 VDD.n1342 VDD.n1205 4.5005
R77357 VDD.n1340 VDD.n1205 4.5005
R77358 VDD.n1344 VDD.n1205 4.5005
R77359 VDD.n1339 VDD.n1205 4.5005
R77360 VDD.n1345 VDD.n1205 4.5005
R77361 VDD.n1338 VDD.n1205 4.5005
R77362 VDD.n1347 VDD.n1205 4.5005
R77363 VDD.n1337 VDD.n1205 4.5005
R77364 VDD.n1348 VDD.n1205 4.5005
R77365 VDD.n1336 VDD.n1205 4.5005
R77366 VDD.n1350 VDD.n1205 4.5005
R77367 VDD.n1335 VDD.n1205 4.5005
R77368 VDD.n1351 VDD.n1205 4.5005
R77369 VDD.n1334 VDD.n1205 4.5005
R77370 VDD.n1353 VDD.n1205 4.5005
R77371 VDD.n1333 VDD.n1205 4.5005
R77372 VDD.n1354 VDD.n1205 4.5005
R77373 VDD.n1332 VDD.n1205 4.5005
R77374 VDD.n1356 VDD.n1205 4.5005
R77375 VDD.n1331 VDD.n1205 4.5005
R77376 VDD.n1357 VDD.n1205 4.5005
R77377 VDD.n1330 VDD.n1205 4.5005
R77378 VDD.n1359 VDD.n1205 4.5005
R77379 VDD.n1329 VDD.n1205 4.5005
R77380 VDD.n1360 VDD.n1205 4.5005
R77381 VDD.n1328 VDD.n1205 4.5005
R77382 VDD.n1362 VDD.n1205 4.5005
R77383 VDD.n1327 VDD.n1205 4.5005
R77384 VDD.n1363 VDD.n1205 4.5005
R77385 VDD.n1326 VDD.n1205 4.5005
R77386 VDD.n1365 VDD.n1205 4.5005
R77387 VDD.n1325 VDD.n1205 4.5005
R77388 VDD.n1366 VDD.n1205 4.5005
R77389 VDD.n1324 VDD.n1205 4.5005
R77390 VDD.n1368 VDD.n1205 4.5005
R77391 VDD.n1323 VDD.n1205 4.5005
R77392 VDD.n1369 VDD.n1205 4.5005
R77393 VDD.n1322 VDD.n1205 4.5005
R77394 VDD.n1371 VDD.n1205 4.5005
R77395 VDD.n1321 VDD.n1205 4.5005
R77396 VDD.n1372 VDD.n1205 4.5005
R77397 VDD.n1320 VDD.n1205 4.5005
R77398 VDD.n1374 VDD.n1205 4.5005
R77399 VDD.n1319 VDD.n1205 4.5005
R77400 VDD.n1375 VDD.n1205 4.5005
R77401 VDD.n1318 VDD.n1205 4.5005
R77402 VDD.n1376 VDD.n1205 4.5005
R77403 VDD.n1316 VDD.n1205 4.5005
R77404 VDD.n1377 VDD.n1205 4.5005
R77405 VDD.n1315 VDD.n1205 4.5005
R77406 VDD.n1378 VDD.n1205 4.5005
R77407 VDD.n1313 VDD.n1205 4.5005
R77408 VDD.n1379 VDD.n1205 4.5005
R77409 VDD.n1312 VDD.n1205 4.5005
R77410 VDD.n1380 VDD.n1205 4.5005
R77411 VDD.n1310 VDD.n1205 4.5005
R77412 VDD.n1381 VDD.n1205 4.5005
R77413 VDD.n1309 VDD.n1205 4.5005
R77414 VDD.n1382 VDD.n1205 4.5005
R77415 VDD.n1307 VDD.n1205 4.5005
R77416 VDD.n1383 VDD.n1205 4.5005
R77417 VDD.n1306 VDD.n1205 4.5005
R77418 VDD.n1384 VDD.n1205 4.5005
R77419 VDD.n1304 VDD.n1205 4.5005
R77420 VDD.n1385 VDD.n1205 4.5005
R77421 VDD.n1303 VDD.n1205 4.5005
R77422 VDD.n1386 VDD.n1205 4.5005
R77423 VDD.n1301 VDD.n1205 4.5005
R77424 VDD.n1387 VDD.n1205 4.5005
R77425 VDD.n1300 VDD.n1205 4.5005
R77426 VDD.n1388 VDD.n1205 4.5005
R77427 VDD.n1298 VDD.n1205 4.5005
R77428 VDD.n1389 VDD.n1205 4.5005
R77429 VDD.n1297 VDD.n1205 4.5005
R77430 VDD.n1390 VDD.n1205 4.5005
R77431 VDD.n1295 VDD.n1205 4.5005
R77432 VDD.n1391 VDD.n1205 4.5005
R77433 VDD.n1294 VDD.n1205 4.5005
R77434 VDD.n1392 VDD.n1205 4.5005
R77435 VDD.n1292 VDD.n1205 4.5005
R77436 VDD.n1393 VDD.n1205 4.5005
R77437 VDD.n1291 VDD.n1205 4.5005
R77438 VDD.n1394 VDD.n1205 4.5005
R77439 VDD.n1289 VDD.n1205 4.5005
R77440 VDD.n1395 VDD.n1205 4.5005
R77441 VDD.n1288 VDD.n1205 4.5005
R77442 VDD.n1396 VDD.n1205 4.5005
R77443 VDD.n1286 VDD.n1205 4.5005
R77444 VDD.n1397 VDD.n1205 4.5005
R77445 VDD.n1285 VDD.n1205 4.5005
R77446 VDD.n1398 VDD.n1205 4.5005
R77447 VDD.n1283 VDD.n1205 4.5005
R77448 VDD.n1399 VDD.n1205 4.5005
R77449 VDD.n1282 VDD.n1205 4.5005
R77450 VDD.n1400 VDD.n1205 4.5005
R77451 VDD.n1280 VDD.n1205 4.5005
R77452 VDD.n1401 VDD.n1205 4.5005
R77453 VDD.n1279 VDD.n1205 4.5005
R77454 VDD.n1402 VDD.n1205 4.5005
R77455 VDD.n1277 VDD.n1205 4.5005
R77456 VDD.n1403 VDD.n1205 4.5005
R77457 VDD.n1276 VDD.n1205 4.5005
R77458 VDD.n1404 VDD.n1205 4.5005
R77459 VDD.n1274 VDD.n1205 4.5005
R77460 VDD.n1405 VDD.n1205 4.5005
R77461 VDD.n1273 VDD.n1205 4.5005
R77462 VDD.n1406 VDD.n1205 4.5005
R77463 VDD.n1271 VDD.n1205 4.5005
R77464 VDD.n1407 VDD.n1205 4.5005
R77465 VDD.n1270 VDD.n1205 4.5005
R77466 VDD.n1408 VDD.n1205 4.5005
R77467 VDD.n1268 VDD.n1205 4.5005
R77468 VDD.n1409 VDD.n1205 4.5005
R77469 VDD.n1267 VDD.n1205 4.5005
R77470 VDD.n1410 VDD.n1205 4.5005
R77471 VDD.n1265 VDD.n1205 4.5005
R77472 VDD.n1411 VDD.n1205 4.5005
R77473 VDD.n1264 VDD.n1205 4.5005
R77474 VDD.n1412 VDD.n1205 4.5005
R77475 VDD.n1262 VDD.n1205 4.5005
R77476 VDD.n1413 VDD.n1205 4.5005
R77477 VDD.n1261 VDD.n1205 4.5005
R77478 VDD.n1414 VDD.n1205 4.5005
R77479 VDD.n1415 VDD.n1205 4.5005
R77480 VDD.n1674 VDD.n1205 4.5005
R77481 VDD.n1676 VDD.n1184 4.5005
R77482 VDD.n1341 VDD.n1184 4.5005
R77483 VDD.n1342 VDD.n1184 4.5005
R77484 VDD.n1340 VDD.n1184 4.5005
R77485 VDD.n1344 VDD.n1184 4.5005
R77486 VDD.n1339 VDD.n1184 4.5005
R77487 VDD.n1345 VDD.n1184 4.5005
R77488 VDD.n1338 VDD.n1184 4.5005
R77489 VDD.n1347 VDD.n1184 4.5005
R77490 VDD.n1337 VDD.n1184 4.5005
R77491 VDD.n1348 VDD.n1184 4.5005
R77492 VDD.n1336 VDD.n1184 4.5005
R77493 VDD.n1350 VDD.n1184 4.5005
R77494 VDD.n1335 VDD.n1184 4.5005
R77495 VDD.n1351 VDD.n1184 4.5005
R77496 VDD.n1334 VDD.n1184 4.5005
R77497 VDD.n1353 VDD.n1184 4.5005
R77498 VDD.n1333 VDD.n1184 4.5005
R77499 VDD.n1354 VDD.n1184 4.5005
R77500 VDD.n1332 VDD.n1184 4.5005
R77501 VDD.n1356 VDD.n1184 4.5005
R77502 VDD.n1331 VDD.n1184 4.5005
R77503 VDD.n1357 VDD.n1184 4.5005
R77504 VDD.n1330 VDD.n1184 4.5005
R77505 VDD.n1359 VDD.n1184 4.5005
R77506 VDD.n1329 VDD.n1184 4.5005
R77507 VDD.n1360 VDD.n1184 4.5005
R77508 VDD.n1328 VDD.n1184 4.5005
R77509 VDD.n1362 VDD.n1184 4.5005
R77510 VDD.n1327 VDD.n1184 4.5005
R77511 VDD.n1363 VDD.n1184 4.5005
R77512 VDD.n1326 VDD.n1184 4.5005
R77513 VDD.n1365 VDD.n1184 4.5005
R77514 VDD.n1325 VDD.n1184 4.5005
R77515 VDD.n1366 VDD.n1184 4.5005
R77516 VDD.n1324 VDD.n1184 4.5005
R77517 VDD.n1368 VDD.n1184 4.5005
R77518 VDD.n1323 VDD.n1184 4.5005
R77519 VDD.n1369 VDD.n1184 4.5005
R77520 VDD.n1322 VDD.n1184 4.5005
R77521 VDD.n1371 VDD.n1184 4.5005
R77522 VDD.n1321 VDD.n1184 4.5005
R77523 VDD.n1372 VDD.n1184 4.5005
R77524 VDD.n1320 VDD.n1184 4.5005
R77525 VDD.n1374 VDD.n1184 4.5005
R77526 VDD.n1319 VDD.n1184 4.5005
R77527 VDD.n1375 VDD.n1184 4.5005
R77528 VDD.n1318 VDD.n1184 4.5005
R77529 VDD.n1376 VDD.n1184 4.5005
R77530 VDD.n1316 VDD.n1184 4.5005
R77531 VDD.n1377 VDD.n1184 4.5005
R77532 VDD.n1315 VDD.n1184 4.5005
R77533 VDD.n1378 VDD.n1184 4.5005
R77534 VDD.n1313 VDD.n1184 4.5005
R77535 VDD.n1379 VDD.n1184 4.5005
R77536 VDD.n1312 VDD.n1184 4.5005
R77537 VDD.n1380 VDD.n1184 4.5005
R77538 VDD.n1310 VDD.n1184 4.5005
R77539 VDD.n1381 VDD.n1184 4.5005
R77540 VDD.n1309 VDD.n1184 4.5005
R77541 VDD.n1382 VDD.n1184 4.5005
R77542 VDD.n1307 VDD.n1184 4.5005
R77543 VDD.n1383 VDD.n1184 4.5005
R77544 VDD.n1306 VDD.n1184 4.5005
R77545 VDD.n1384 VDD.n1184 4.5005
R77546 VDD.n1304 VDD.n1184 4.5005
R77547 VDD.n1385 VDD.n1184 4.5005
R77548 VDD.n1303 VDD.n1184 4.5005
R77549 VDD.n1386 VDD.n1184 4.5005
R77550 VDD.n1301 VDD.n1184 4.5005
R77551 VDD.n1387 VDD.n1184 4.5005
R77552 VDD.n1300 VDD.n1184 4.5005
R77553 VDD.n1388 VDD.n1184 4.5005
R77554 VDD.n1298 VDD.n1184 4.5005
R77555 VDD.n1389 VDD.n1184 4.5005
R77556 VDD.n1297 VDD.n1184 4.5005
R77557 VDD.n1390 VDD.n1184 4.5005
R77558 VDD.n1295 VDD.n1184 4.5005
R77559 VDD.n1391 VDD.n1184 4.5005
R77560 VDD.n1294 VDD.n1184 4.5005
R77561 VDD.n1392 VDD.n1184 4.5005
R77562 VDD.n1292 VDD.n1184 4.5005
R77563 VDD.n1393 VDD.n1184 4.5005
R77564 VDD.n1291 VDD.n1184 4.5005
R77565 VDD.n1394 VDD.n1184 4.5005
R77566 VDD.n1289 VDD.n1184 4.5005
R77567 VDD.n1395 VDD.n1184 4.5005
R77568 VDD.n1288 VDD.n1184 4.5005
R77569 VDD.n1396 VDD.n1184 4.5005
R77570 VDD.n1286 VDD.n1184 4.5005
R77571 VDD.n1397 VDD.n1184 4.5005
R77572 VDD.n1285 VDD.n1184 4.5005
R77573 VDD.n1398 VDD.n1184 4.5005
R77574 VDD.n1283 VDD.n1184 4.5005
R77575 VDD.n1399 VDD.n1184 4.5005
R77576 VDD.n1282 VDD.n1184 4.5005
R77577 VDD.n1400 VDD.n1184 4.5005
R77578 VDD.n1280 VDD.n1184 4.5005
R77579 VDD.n1401 VDD.n1184 4.5005
R77580 VDD.n1279 VDD.n1184 4.5005
R77581 VDD.n1402 VDD.n1184 4.5005
R77582 VDD.n1277 VDD.n1184 4.5005
R77583 VDD.n1403 VDD.n1184 4.5005
R77584 VDD.n1276 VDD.n1184 4.5005
R77585 VDD.n1404 VDD.n1184 4.5005
R77586 VDD.n1274 VDD.n1184 4.5005
R77587 VDD.n1405 VDD.n1184 4.5005
R77588 VDD.n1273 VDD.n1184 4.5005
R77589 VDD.n1406 VDD.n1184 4.5005
R77590 VDD.n1271 VDD.n1184 4.5005
R77591 VDD.n1407 VDD.n1184 4.5005
R77592 VDD.n1270 VDD.n1184 4.5005
R77593 VDD.n1408 VDD.n1184 4.5005
R77594 VDD.n1268 VDD.n1184 4.5005
R77595 VDD.n1409 VDD.n1184 4.5005
R77596 VDD.n1267 VDD.n1184 4.5005
R77597 VDD.n1410 VDD.n1184 4.5005
R77598 VDD.n1265 VDD.n1184 4.5005
R77599 VDD.n1411 VDD.n1184 4.5005
R77600 VDD.n1264 VDD.n1184 4.5005
R77601 VDD.n1412 VDD.n1184 4.5005
R77602 VDD.n1262 VDD.n1184 4.5005
R77603 VDD.n1413 VDD.n1184 4.5005
R77604 VDD.n1261 VDD.n1184 4.5005
R77605 VDD.n1414 VDD.n1184 4.5005
R77606 VDD.n1415 VDD.n1184 4.5005
R77607 VDD.n1674 VDD.n1184 4.5005
R77608 VDD.n1676 VDD.n1206 4.5005
R77609 VDD.n1341 VDD.n1206 4.5005
R77610 VDD.n1342 VDD.n1206 4.5005
R77611 VDD.n1340 VDD.n1206 4.5005
R77612 VDD.n1344 VDD.n1206 4.5005
R77613 VDD.n1339 VDD.n1206 4.5005
R77614 VDD.n1345 VDD.n1206 4.5005
R77615 VDD.n1338 VDD.n1206 4.5005
R77616 VDD.n1347 VDD.n1206 4.5005
R77617 VDD.n1337 VDD.n1206 4.5005
R77618 VDD.n1348 VDD.n1206 4.5005
R77619 VDD.n1336 VDD.n1206 4.5005
R77620 VDD.n1350 VDD.n1206 4.5005
R77621 VDD.n1335 VDD.n1206 4.5005
R77622 VDD.n1351 VDD.n1206 4.5005
R77623 VDD.n1334 VDD.n1206 4.5005
R77624 VDD.n1353 VDD.n1206 4.5005
R77625 VDD.n1333 VDD.n1206 4.5005
R77626 VDD.n1354 VDD.n1206 4.5005
R77627 VDD.n1332 VDD.n1206 4.5005
R77628 VDD.n1356 VDD.n1206 4.5005
R77629 VDD.n1331 VDD.n1206 4.5005
R77630 VDD.n1357 VDD.n1206 4.5005
R77631 VDD.n1330 VDD.n1206 4.5005
R77632 VDD.n1359 VDD.n1206 4.5005
R77633 VDD.n1329 VDD.n1206 4.5005
R77634 VDD.n1360 VDD.n1206 4.5005
R77635 VDD.n1328 VDD.n1206 4.5005
R77636 VDD.n1362 VDD.n1206 4.5005
R77637 VDD.n1327 VDD.n1206 4.5005
R77638 VDD.n1363 VDD.n1206 4.5005
R77639 VDD.n1326 VDD.n1206 4.5005
R77640 VDD.n1365 VDD.n1206 4.5005
R77641 VDD.n1325 VDD.n1206 4.5005
R77642 VDD.n1366 VDD.n1206 4.5005
R77643 VDD.n1324 VDD.n1206 4.5005
R77644 VDD.n1368 VDD.n1206 4.5005
R77645 VDD.n1323 VDD.n1206 4.5005
R77646 VDD.n1369 VDD.n1206 4.5005
R77647 VDD.n1322 VDD.n1206 4.5005
R77648 VDD.n1371 VDD.n1206 4.5005
R77649 VDD.n1321 VDD.n1206 4.5005
R77650 VDD.n1372 VDD.n1206 4.5005
R77651 VDD.n1320 VDD.n1206 4.5005
R77652 VDD.n1374 VDD.n1206 4.5005
R77653 VDD.n1319 VDD.n1206 4.5005
R77654 VDD.n1375 VDD.n1206 4.5005
R77655 VDD.n1318 VDD.n1206 4.5005
R77656 VDD.n1376 VDD.n1206 4.5005
R77657 VDD.n1316 VDD.n1206 4.5005
R77658 VDD.n1377 VDD.n1206 4.5005
R77659 VDD.n1315 VDD.n1206 4.5005
R77660 VDD.n1378 VDD.n1206 4.5005
R77661 VDD.n1313 VDD.n1206 4.5005
R77662 VDD.n1379 VDD.n1206 4.5005
R77663 VDD.n1312 VDD.n1206 4.5005
R77664 VDD.n1380 VDD.n1206 4.5005
R77665 VDD.n1310 VDD.n1206 4.5005
R77666 VDD.n1381 VDD.n1206 4.5005
R77667 VDD.n1309 VDD.n1206 4.5005
R77668 VDD.n1382 VDD.n1206 4.5005
R77669 VDD.n1307 VDD.n1206 4.5005
R77670 VDD.n1383 VDD.n1206 4.5005
R77671 VDD.n1306 VDD.n1206 4.5005
R77672 VDD.n1384 VDD.n1206 4.5005
R77673 VDD.n1304 VDD.n1206 4.5005
R77674 VDD.n1385 VDD.n1206 4.5005
R77675 VDD.n1303 VDD.n1206 4.5005
R77676 VDD.n1386 VDD.n1206 4.5005
R77677 VDD.n1301 VDD.n1206 4.5005
R77678 VDD.n1387 VDD.n1206 4.5005
R77679 VDD.n1300 VDD.n1206 4.5005
R77680 VDD.n1388 VDD.n1206 4.5005
R77681 VDD.n1298 VDD.n1206 4.5005
R77682 VDD.n1389 VDD.n1206 4.5005
R77683 VDD.n1297 VDD.n1206 4.5005
R77684 VDD.n1390 VDD.n1206 4.5005
R77685 VDD.n1295 VDD.n1206 4.5005
R77686 VDD.n1391 VDD.n1206 4.5005
R77687 VDD.n1294 VDD.n1206 4.5005
R77688 VDD.n1392 VDD.n1206 4.5005
R77689 VDD.n1292 VDD.n1206 4.5005
R77690 VDD.n1393 VDD.n1206 4.5005
R77691 VDD.n1291 VDD.n1206 4.5005
R77692 VDD.n1394 VDD.n1206 4.5005
R77693 VDD.n1289 VDD.n1206 4.5005
R77694 VDD.n1395 VDD.n1206 4.5005
R77695 VDD.n1288 VDD.n1206 4.5005
R77696 VDD.n1396 VDD.n1206 4.5005
R77697 VDD.n1286 VDD.n1206 4.5005
R77698 VDD.n1397 VDD.n1206 4.5005
R77699 VDD.n1285 VDD.n1206 4.5005
R77700 VDD.n1398 VDD.n1206 4.5005
R77701 VDD.n1283 VDD.n1206 4.5005
R77702 VDD.n1399 VDD.n1206 4.5005
R77703 VDD.n1282 VDD.n1206 4.5005
R77704 VDD.n1400 VDD.n1206 4.5005
R77705 VDD.n1280 VDD.n1206 4.5005
R77706 VDD.n1401 VDD.n1206 4.5005
R77707 VDD.n1279 VDD.n1206 4.5005
R77708 VDD.n1402 VDD.n1206 4.5005
R77709 VDD.n1277 VDD.n1206 4.5005
R77710 VDD.n1403 VDD.n1206 4.5005
R77711 VDD.n1276 VDD.n1206 4.5005
R77712 VDD.n1404 VDD.n1206 4.5005
R77713 VDD.n1274 VDD.n1206 4.5005
R77714 VDD.n1405 VDD.n1206 4.5005
R77715 VDD.n1273 VDD.n1206 4.5005
R77716 VDD.n1406 VDD.n1206 4.5005
R77717 VDD.n1271 VDD.n1206 4.5005
R77718 VDD.n1407 VDD.n1206 4.5005
R77719 VDD.n1270 VDD.n1206 4.5005
R77720 VDD.n1408 VDD.n1206 4.5005
R77721 VDD.n1268 VDD.n1206 4.5005
R77722 VDD.n1409 VDD.n1206 4.5005
R77723 VDD.n1267 VDD.n1206 4.5005
R77724 VDD.n1410 VDD.n1206 4.5005
R77725 VDD.n1265 VDD.n1206 4.5005
R77726 VDD.n1411 VDD.n1206 4.5005
R77727 VDD.n1264 VDD.n1206 4.5005
R77728 VDD.n1412 VDD.n1206 4.5005
R77729 VDD.n1262 VDD.n1206 4.5005
R77730 VDD.n1413 VDD.n1206 4.5005
R77731 VDD.n1261 VDD.n1206 4.5005
R77732 VDD.n1414 VDD.n1206 4.5005
R77733 VDD.n1415 VDD.n1206 4.5005
R77734 VDD.n1674 VDD.n1206 4.5005
R77735 VDD.n1676 VDD.n1183 4.5005
R77736 VDD.n1341 VDD.n1183 4.5005
R77737 VDD.n1342 VDD.n1183 4.5005
R77738 VDD.n1340 VDD.n1183 4.5005
R77739 VDD.n1344 VDD.n1183 4.5005
R77740 VDD.n1339 VDD.n1183 4.5005
R77741 VDD.n1345 VDD.n1183 4.5005
R77742 VDD.n1338 VDD.n1183 4.5005
R77743 VDD.n1347 VDD.n1183 4.5005
R77744 VDD.n1337 VDD.n1183 4.5005
R77745 VDD.n1348 VDD.n1183 4.5005
R77746 VDD.n1336 VDD.n1183 4.5005
R77747 VDD.n1350 VDD.n1183 4.5005
R77748 VDD.n1335 VDD.n1183 4.5005
R77749 VDD.n1351 VDD.n1183 4.5005
R77750 VDD.n1334 VDD.n1183 4.5005
R77751 VDD.n1353 VDD.n1183 4.5005
R77752 VDD.n1333 VDD.n1183 4.5005
R77753 VDD.n1354 VDD.n1183 4.5005
R77754 VDD.n1332 VDD.n1183 4.5005
R77755 VDD.n1356 VDD.n1183 4.5005
R77756 VDD.n1331 VDD.n1183 4.5005
R77757 VDD.n1357 VDD.n1183 4.5005
R77758 VDD.n1330 VDD.n1183 4.5005
R77759 VDD.n1359 VDD.n1183 4.5005
R77760 VDD.n1329 VDD.n1183 4.5005
R77761 VDD.n1360 VDD.n1183 4.5005
R77762 VDD.n1328 VDD.n1183 4.5005
R77763 VDD.n1362 VDD.n1183 4.5005
R77764 VDD.n1327 VDD.n1183 4.5005
R77765 VDD.n1363 VDD.n1183 4.5005
R77766 VDD.n1326 VDD.n1183 4.5005
R77767 VDD.n1365 VDD.n1183 4.5005
R77768 VDD.n1325 VDD.n1183 4.5005
R77769 VDD.n1366 VDD.n1183 4.5005
R77770 VDD.n1324 VDD.n1183 4.5005
R77771 VDD.n1368 VDD.n1183 4.5005
R77772 VDD.n1323 VDD.n1183 4.5005
R77773 VDD.n1369 VDD.n1183 4.5005
R77774 VDD.n1322 VDD.n1183 4.5005
R77775 VDD.n1371 VDD.n1183 4.5005
R77776 VDD.n1321 VDD.n1183 4.5005
R77777 VDD.n1372 VDD.n1183 4.5005
R77778 VDD.n1320 VDD.n1183 4.5005
R77779 VDD.n1374 VDD.n1183 4.5005
R77780 VDD.n1319 VDD.n1183 4.5005
R77781 VDD.n1375 VDD.n1183 4.5005
R77782 VDD.n1318 VDD.n1183 4.5005
R77783 VDD.n1376 VDD.n1183 4.5005
R77784 VDD.n1316 VDD.n1183 4.5005
R77785 VDD.n1377 VDD.n1183 4.5005
R77786 VDD.n1315 VDD.n1183 4.5005
R77787 VDD.n1378 VDD.n1183 4.5005
R77788 VDD.n1313 VDD.n1183 4.5005
R77789 VDD.n1379 VDD.n1183 4.5005
R77790 VDD.n1312 VDD.n1183 4.5005
R77791 VDD.n1380 VDD.n1183 4.5005
R77792 VDD.n1310 VDD.n1183 4.5005
R77793 VDD.n1381 VDD.n1183 4.5005
R77794 VDD.n1309 VDD.n1183 4.5005
R77795 VDD.n1382 VDD.n1183 4.5005
R77796 VDD.n1307 VDD.n1183 4.5005
R77797 VDD.n1383 VDD.n1183 4.5005
R77798 VDD.n1306 VDD.n1183 4.5005
R77799 VDD.n1384 VDD.n1183 4.5005
R77800 VDD.n1304 VDD.n1183 4.5005
R77801 VDD.n1385 VDD.n1183 4.5005
R77802 VDD.n1303 VDD.n1183 4.5005
R77803 VDD.n1386 VDD.n1183 4.5005
R77804 VDD.n1301 VDD.n1183 4.5005
R77805 VDD.n1387 VDD.n1183 4.5005
R77806 VDD.n1300 VDD.n1183 4.5005
R77807 VDD.n1388 VDD.n1183 4.5005
R77808 VDD.n1298 VDD.n1183 4.5005
R77809 VDD.n1389 VDD.n1183 4.5005
R77810 VDD.n1297 VDD.n1183 4.5005
R77811 VDD.n1390 VDD.n1183 4.5005
R77812 VDD.n1295 VDD.n1183 4.5005
R77813 VDD.n1391 VDD.n1183 4.5005
R77814 VDD.n1294 VDD.n1183 4.5005
R77815 VDD.n1392 VDD.n1183 4.5005
R77816 VDD.n1292 VDD.n1183 4.5005
R77817 VDD.n1393 VDD.n1183 4.5005
R77818 VDD.n1291 VDD.n1183 4.5005
R77819 VDD.n1394 VDD.n1183 4.5005
R77820 VDD.n1289 VDD.n1183 4.5005
R77821 VDD.n1395 VDD.n1183 4.5005
R77822 VDD.n1288 VDD.n1183 4.5005
R77823 VDD.n1396 VDD.n1183 4.5005
R77824 VDD.n1286 VDD.n1183 4.5005
R77825 VDD.n1397 VDD.n1183 4.5005
R77826 VDD.n1285 VDD.n1183 4.5005
R77827 VDD.n1398 VDD.n1183 4.5005
R77828 VDD.n1283 VDD.n1183 4.5005
R77829 VDD.n1399 VDD.n1183 4.5005
R77830 VDD.n1282 VDD.n1183 4.5005
R77831 VDD.n1400 VDD.n1183 4.5005
R77832 VDD.n1280 VDD.n1183 4.5005
R77833 VDD.n1401 VDD.n1183 4.5005
R77834 VDD.n1279 VDD.n1183 4.5005
R77835 VDD.n1402 VDD.n1183 4.5005
R77836 VDD.n1277 VDD.n1183 4.5005
R77837 VDD.n1403 VDD.n1183 4.5005
R77838 VDD.n1276 VDD.n1183 4.5005
R77839 VDD.n1404 VDD.n1183 4.5005
R77840 VDD.n1274 VDD.n1183 4.5005
R77841 VDD.n1405 VDD.n1183 4.5005
R77842 VDD.n1273 VDD.n1183 4.5005
R77843 VDD.n1406 VDD.n1183 4.5005
R77844 VDD.n1271 VDD.n1183 4.5005
R77845 VDD.n1407 VDD.n1183 4.5005
R77846 VDD.n1270 VDD.n1183 4.5005
R77847 VDD.n1408 VDD.n1183 4.5005
R77848 VDD.n1268 VDD.n1183 4.5005
R77849 VDD.n1409 VDD.n1183 4.5005
R77850 VDD.n1267 VDD.n1183 4.5005
R77851 VDD.n1410 VDD.n1183 4.5005
R77852 VDD.n1265 VDD.n1183 4.5005
R77853 VDD.n1411 VDD.n1183 4.5005
R77854 VDD.n1264 VDD.n1183 4.5005
R77855 VDD.n1412 VDD.n1183 4.5005
R77856 VDD.n1262 VDD.n1183 4.5005
R77857 VDD.n1413 VDD.n1183 4.5005
R77858 VDD.n1261 VDD.n1183 4.5005
R77859 VDD.n1414 VDD.n1183 4.5005
R77860 VDD.n1415 VDD.n1183 4.5005
R77861 VDD.n1674 VDD.n1183 4.5005
R77862 VDD.n1676 VDD.n1207 4.5005
R77863 VDD.n1341 VDD.n1207 4.5005
R77864 VDD.n1342 VDD.n1207 4.5005
R77865 VDD.n1340 VDD.n1207 4.5005
R77866 VDD.n1344 VDD.n1207 4.5005
R77867 VDD.n1339 VDD.n1207 4.5005
R77868 VDD.n1345 VDD.n1207 4.5005
R77869 VDD.n1338 VDD.n1207 4.5005
R77870 VDD.n1347 VDD.n1207 4.5005
R77871 VDD.n1337 VDD.n1207 4.5005
R77872 VDD.n1348 VDD.n1207 4.5005
R77873 VDD.n1336 VDD.n1207 4.5005
R77874 VDD.n1350 VDD.n1207 4.5005
R77875 VDD.n1335 VDD.n1207 4.5005
R77876 VDD.n1351 VDD.n1207 4.5005
R77877 VDD.n1334 VDD.n1207 4.5005
R77878 VDD.n1353 VDD.n1207 4.5005
R77879 VDD.n1333 VDD.n1207 4.5005
R77880 VDD.n1354 VDD.n1207 4.5005
R77881 VDD.n1332 VDD.n1207 4.5005
R77882 VDD.n1356 VDD.n1207 4.5005
R77883 VDD.n1331 VDD.n1207 4.5005
R77884 VDD.n1357 VDD.n1207 4.5005
R77885 VDD.n1330 VDD.n1207 4.5005
R77886 VDD.n1359 VDD.n1207 4.5005
R77887 VDD.n1329 VDD.n1207 4.5005
R77888 VDD.n1360 VDD.n1207 4.5005
R77889 VDD.n1328 VDD.n1207 4.5005
R77890 VDD.n1362 VDD.n1207 4.5005
R77891 VDD.n1327 VDD.n1207 4.5005
R77892 VDD.n1363 VDD.n1207 4.5005
R77893 VDD.n1326 VDD.n1207 4.5005
R77894 VDD.n1365 VDD.n1207 4.5005
R77895 VDD.n1325 VDD.n1207 4.5005
R77896 VDD.n1366 VDD.n1207 4.5005
R77897 VDD.n1324 VDD.n1207 4.5005
R77898 VDD.n1368 VDD.n1207 4.5005
R77899 VDD.n1323 VDD.n1207 4.5005
R77900 VDD.n1369 VDD.n1207 4.5005
R77901 VDD.n1322 VDD.n1207 4.5005
R77902 VDD.n1371 VDD.n1207 4.5005
R77903 VDD.n1321 VDD.n1207 4.5005
R77904 VDD.n1372 VDD.n1207 4.5005
R77905 VDD.n1320 VDD.n1207 4.5005
R77906 VDD.n1374 VDD.n1207 4.5005
R77907 VDD.n1319 VDD.n1207 4.5005
R77908 VDD.n1375 VDD.n1207 4.5005
R77909 VDD.n1318 VDD.n1207 4.5005
R77910 VDD.n1376 VDD.n1207 4.5005
R77911 VDD.n1316 VDD.n1207 4.5005
R77912 VDD.n1377 VDD.n1207 4.5005
R77913 VDD.n1315 VDD.n1207 4.5005
R77914 VDD.n1378 VDD.n1207 4.5005
R77915 VDD.n1313 VDD.n1207 4.5005
R77916 VDD.n1379 VDD.n1207 4.5005
R77917 VDD.n1312 VDD.n1207 4.5005
R77918 VDD.n1380 VDD.n1207 4.5005
R77919 VDD.n1310 VDD.n1207 4.5005
R77920 VDD.n1381 VDD.n1207 4.5005
R77921 VDD.n1309 VDD.n1207 4.5005
R77922 VDD.n1382 VDD.n1207 4.5005
R77923 VDD.n1307 VDD.n1207 4.5005
R77924 VDD.n1383 VDD.n1207 4.5005
R77925 VDD.n1306 VDD.n1207 4.5005
R77926 VDD.n1384 VDD.n1207 4.5005
R77927 VDD.n1304 VDD.n1207 4.5005
R77928 VDD.n1385 VDD.n1207 4.5005
R77929 VDD.n1303 VDD.n1207 4.5005
R77930 VDD.n1386 VDD.n1207 4.5005
R77931 VDD.n1301 VDD.n1207 4.5005
R77932 VDD.n1387 VDD.n1207 4.5005
R77933 VDD.n1300 VDD.n1207 4.5005
R77934 VDD.n1388 VDD.n1207 4.5005
R77935 VDD.n1298 VDD.n1207 4.5005
R77936 VDD.n1389 VDD.n1207 4.5005
R77937 VDD.n1297 VDD.n1207 4.5005
R77938 VDD.n1390 VDD.n1207 4.5005
R77939 VDD.n1295 VDD.n1207 4.5005
R77940 VDD.n1391 VDD.n1207 4.5005
R77941 VDD.n1294 VDD.n1207 4.5005
R77942 VDD.n1392 VDD.n1207 4.5005
R77943 VDD.n1292 VDD.n1207 4.5005
R77944 VDD.n1393 VDD.n1207 4.5005
R77945 VDD.n1291 VDD.n1207 4.5005
R77946 VDD.n1394 VDD.n1207 4.5005
R77947 VDD.n1289 VDD.n1207 4.5005
R77948 VDD.n1395 VDD.n1207 4.5005
R77949 VDD.n1288 VDD.n1207 4.5005
R77950 VDD.n1396 VDD.n1207 4.5005
R77951 VDD.n1286 VDD.n1207 4.5005
R77952 VDD.n1397 VDD.n1207 4.5005
R77953 VDD.n1285 VDD.n1207 4.5005
R77954 VDD.n1398 VDD.n1207 4.5005
R77955 VDD.n1283 VDD.n1207 4.5005
R77956 VDD.n1399 VDD.n1207 4.5005
R77957 VDD.n1282 VDD.n1207 4.5005
R77958 VDD.n1400 VDD.n1207 4.5005
R77959 VDD.n1280 VDD.n1207 4.5005
R77960 VDD.n1401 VDD.n1207 4.5005
R77961 VDD.n1279 VDD.n1207 4.5005
R77962 VDD.n1402 VDD.n1207 4.5005
R77963 VDD.n1277 VDD.n1207 4.5005
R77964 VDD.n1403 VDD.n1207 4.5005
R77965 VDD.n1276 VDD.n1207 4.5005
R77966 VDD.n1404 VDD.n1207 4.5005
R77967 VDD.n1274 VDD.n1207 4.5005
R77968 VDD.n1405 VDD.n1207 4.5005
R77969 VDD.n1273 VDD.n1207 4.5005
R77970 VDD.n1406 VDD.n1207 4.5005
R77971 VDD.n1271 VDD.n1207 4.5005
R77972 VDD.n1407 VDD.n1207 4.5005
R77973 VDD.n1270 VDD.n1207 4.5005
R77974 VDD.n1408 VDD.n1207 4.5005
R77975 VDD.n1268 VDD.n1207 4.5005
R77976 VDD.n1409 VDD.n1207 4.5005
R77977 VDD.n1267 VDD.n1207 4.5005
R77978 VDD.n1410 VDD.n1207 4.5005
R77979 VDD.n1265 VDD.n1207 4.5005
R77980 VDD.n1411 VDD.n1207 4.5005
R77981 VDD.n1264 VDD.n1207 4.5005
R77982 VDD.n1412 VDD.n1207 4.5005
R77983 VDD.n1262 VDD.n1207 4.5005
R77984 VDD.n1413 VDD.n1207 4.5005
R77985 VDD.n1261 VDD.n1207 4.5005
R77986 VDD.n1414 VDD.n1207 4.5005
R77987 VDD.n1415 VDD.n1207 4.5005
R77988 VDD.n1674 VDD.n1207 4.5005
R77989 VDD.n1676 VDD.n1182 4.5005
R77990 VDD.n1341 VDD.n1182 4.5005
R77991 VDD.n1342 VDD.n1182 4.5005
R77992 VDD.n1340 VDD.n1182 4.5005
R77993 VDD.n1344 VDD.n1182 4.5005
R77994 VDD.n1339 VDD.n1182 4.5005
R77995 VDD.n1345 VDD.n1182 4.5005
R77996 VDD.n1338 VDD.n1182 4.5005
R77997 VDD.n1347 VDD.n1182 4.5005
R77998 VDD.n1337 VDD.n1182 4.5005
R77999 VDD.n1348 VDD.n1182 4.5005
R78000 VDD.n1336 VDD.n1182 4.5005
R78001 VDD.n1350 VDD.n1182 4.5005
R78002 VDD.n1335 VDD.n1182 4.5005
R78003 VDD.n1351 VDD.n1182 4.5005
R78004 VDD.n1334 VDD.n1182 4.5005
R78005 VDD.n1353 VDD.n1182 4.5005
R78006 VDD.n1333 VDD.n1182 4.5005
R78007 VDD.n1354 VDD.n1182 4.5005
R78008 VDD.n1332 VDD.n1182 4.5005
R78009 VDD.n1356 VDD.n1182 4.5005
R78010 VDD.n1331 VDD.n1182 4.5005
R78011 VDD.n1357 VDD.n1182 4.5005
R78012 VDD.n1330 VDD.n1182 4.5005
R78013 VDD.n1359 VDD.n1182 4.5005
R78014 VDD.n1329 VDD.n1182 4.5005
R78015 VDD.n1360 VDD.n1182 4.5005
R78016 VDD.n1328 VDD.n1182 4.5005
R78017 VDD.n1362 VDD.n1182 4.5005
R78018 VDD.n1327 VDD.n1182 4.5005
R78019 VDD.n1363 VDD.n1182 4.5005
R78020 VDD.n1326 VDD.n1182 4.5005
R78021 VDD.n1365 VDD.n1182 4.5005
R78022 VDD.n1325 VDD.n1182 4.5005
R78023 VDD.n1366 VDD.n1182 4.5005
R78024 VDD.n1324 VDD.n1182 4.5005
R78025 VDD.n1368 VDD.n1182 4.5005
R78026 VDD.n1323 VDD.n1182 4.5005
R78027 VDD.n1369 VDD.n1182 4.5005
R78028 VDD.n1322 VDD.n1182 4.5005
R78029 VDD.n1371 VDD.n1182 4.5005
R78030 VDD.n1321 VDD.n1182 4.5005
R78031 VDD.n1372 VDD.n1182 4.5005
R78032 VDD.n1320 VDD.n1182 4.5005
R78033 VDD.n1374 VDD.n1182 4.5005
R78034 VDD.n1319 VDD.n1182 4.5005
R78035 VDD.n1375 VDD.n1182 4.5005
R78036 VDD.n1318 VDD.n1182 4.5005
R78037 VDD.n1376 VDD.n1182 4.5005
R78038 VDD.n1316 VDD.n1182 4.5005
R78039 VDD.n1377 VDD.n1182 4.5005
R78040 VDD.n1315 VDD.n1182 4.5005
R78041 VDD.n1378 VDD.n1182 4.5005
R78042 VDD.n1313 VDD.n1182 4.5005
R78043 VDD.n1379 VDD.n1182 4.5005
R78044 VDD.n1312 VDD.n1182 4.5005
R78045 VDD.n1380 VDD.n1182 4.5005
R78046 VDD.n1310 VDD.n1182 4.5005
R78047 VDD.n1381 VDD.n1182 4.5005
R78048 VDD.n1309 VDD.n1182 4.5005
R78049 VDD.n1382 VDD.n1182 4.5005
R78050 VDD.n1307 VDD.n1182 4.5005
R78051 VDD.n1383 VDD.n1182 4.5005
R78052 VDD.n1306 VDD.n1182 4.5005
R78053 VDD.n1384 VDD.n1182 4.5005
R78054 VDD.n1304 VDD.n1182 4.5005
R78055 VDD.n1385 VDD.n1182 4.5005
R78056 VDD.n1303 VDD.n1182 4.5005
R78057 VDD.n1386 VDD.n1182 4.5005
R78058 VDD.n1301 VDD.n1182 4.5005
R78059 VDD.n1387 VDD.n1182 4.5005
R78060 VDD.n1300 VDD.n1182 4.5005
R78061 VDD.n1388 VDD.n1182 4.5005
R78062 VDD.n1298 VDD.n1182 4.5005
R78063 VDD.n1389 VDD.n1182 4.5005
R78064 VDD.n1297 VDD.n1182 4.5005
R78065 VDD.n1390 VDD.n1182 4.5005
R78066 VDD.n1295 VDD.n1182 4.5005
R78067 VDD.n1391 VDD.n1182 4.5005
R78068 VDD.n1294 VDD.n1182 4.5005
R78069 VDD.n1392 VDD.n1182 4.5005
R78070 VDD.n1292 VDD.n1182 4.5005
R78071 VDD.n1393 VDD.n1182 4.5005
R78072 VDD.n1291 VDD.n1182 4.5005
R78073 VDD.n1394 VDD.n1182 4.5005
R78074 VDD.n1289 VDD.n1182 4.5005
R78075 VDD.n1395 VDD.n1182 4.5005
R78076 VDD.n1288 VDD.n1182 4.5005
R78077 VDD.n1396 VDD.n1182 4.5005
R78078 VDD.n1286 VDD.n1182 4.5005
R78079 VDD.n1397 VDD.n1182 4.5005
R78080 VDD.n1285 VDD.n1182 4.5005
R78081 VDD.n1398 VDD.n1182 4.5005
R78082 VDD.n1283 VDD.n1182 4.5005
R78083 VDD.n1399 VDD.n1182 4.5005
R78084 VDD.n1282 VDD.n1182 4.5005
R78085 VDD.n1400 VDD.n1182 4.5005
R78086 VDD.n1280 VDD.n1182 4.5005
R78087 VDD.n1401 VDD.n1182 4.5005
R78088 VDD.n1279 VDD.n1182 4.5005
R78089 VDD.n1402 VDD.n1182 4.5005
R78090 VDD.n1277 VDD.n1182 4.5005
R78091 VDD.n1403 VDD.n1182 4.5005
R78092 VDD.n1276 VDD.n1182 4.5005
R78093 VDD.n1404 VDD.n1182 4.5005
R78094 VDD.n1274 VDD.n1182 4.5005
R78095 VDD.n1405 VDD.n1182 4.5005
R78096 VDD.n1273 VDD.n1182 4.5005
R78097 VDD.n1406 VDD.n1182 4.5005
R78098 VDD.n1271 VDD.n1182 4.5005
R78099 VDD.n1407 VDD.n1182 4.5005
R78100 VDD.n1270 VDD.n1182 4.5005
R78101 VDD.n1408 VDD.n1182 4.5005
R78102 VDD.n1268 VDD.n1182 4.5005
R78103 VDD.n1409 VDD.n1182 4.5005
R78104 VDD.n1267 VDD.n1182 4.5005
R78105 VDD.n1410 VDD.n1182 4.5005
R78106 VDD.n1265 VDD.n1182 4.5005
R78107 VDD.n1411 VDD.n1182 4.5005
R78108 VDD.n1264 VDD.n1182 4.5005
R78109 VDD.n1412 VDD.n1182 4.5005
R78110 VDD.n1262 VDD.n1182 4.5005
R78111 VDD.n1413 VDD.n1182 4.5005
R78112 VDD.n1261 VDD.n1182 4.5005
R78113 VDD.n1414 VDD.n1182 4.5005
R78114 VDD.n1415 VDD.n1182 4.5005
R78115 VDD.n1674 VDD.n1182 4.5005
R78116 VDD.n1676 VDD.n1208 4.5005
R78117 VDD.n1341 VDD.n1208 4.5005
R78118 VDD.n1342 VDD.n1208 4.5005
R78119 VDD.n1340 VDD.n1208 4.5005
R78120 VDD.n1344 VDD.n1208 4.5005
R78121 VDD.n1339 VDD.n1208 4.5005
R78122 VDD.n1345 VDD.n1208 4.5005
R78123 VDD.n1338 VDD.n1208 4.5005
R78124 VDD.n1347 VDD.n1208 4.5005
R78125 VDD.n1337 VDD.n1208 4.5005
R78126 VDD.n1348 VDD.n1208 4.5005
R78127 VDD.n1336 VDD.n1208 4.5005
R78128 VDD.n1350 VDD.n1208 4.5005
R78129 VDD.n1335 VDD.n1208 4.5005
R78130 VDD.n1351 VDD.n1208 4.5005
R78131 VDD.n1334 VDD.n1208 4.5005
R78132 VDD.n1353 VDD.n1208 4.5005
R78133 VDD.n1333 VDD.n1208 4.5005
R78134 VDD.n1354 VDD.n1208 4.5005
R78135 VDD.n1332 VDD.n1208 4.5005
R78136 VDD.n1356 VDD.n1208 4.5005
R78137 VDD.n1331 VDD.n1208 4.5005
R78138 VDD.n1357 VDD.n1208 4.5005
R78139 VDD.n1330 VDD.n1208 4.5005
R78140 VDD.n1359 VDD.n1208 4.5005
R78141 VDD.n1329 VDD.n1208 4.5005
R78142 VDD.n1360 VDD.n1208 4.5005
R78143 VDD.n1328 VDD.n1208 4.5005
R78144 VDD.n1362 VDD.n1208 4.5005
R78145 VDD.n1327 VDD.n1208 4.5005
R78146 VDD.n1363 VDD.n1208 4.5005
R78147 VDD.n1326 VDD.n1208 4.5005
R78148 VDD.n1365 VDD.n1208 4.5005
R78149 VDD.n1325 VDD.n1208 4.5005
R78150 VDD.n1366 VDD.n1208 4.5005
R78151 VDD.n1324 VDD.n1208 4.5005
R78152 VDD.n1368 VDD.n1208 4.5005
R78153 VDD.n1323 VDD.n1208 4.5005
R78154 VDD.n1369 VDD.n1208 4.5005
R78155 VDD.n1322 VDD.n1208 4.5005
R78156 VDD.n1371 VDD.n1208 4.5005
R78157 VDD.n1321 VDD.n1208 4.5005
R78158 VDD.n1372 VDD.n1208 4.5005
R78159 VDD.n1320 VDD.n1208 4.5005
R78160 VDD.n1374 VDD.n1208 4.5005
R78161 VDD.n1319 VDD.n1208 4.5005
R78162 VDD.n1375 VDD.n1208 4.5005
R78163 VDD.n1318 VDD.n1208 4.5005
R78164 VDD.n1376 VDD.n1208 4.5005
R78165 VDD.n1316 VDD.n1208 4.5005
R78166 VDD.n1377 VDD.n1208 4.5005
R78167 VDD.n1315 VDD.n1208 4.5005
R78168 VDD.n1378 VDD.n1208 4.5005
R78169 VDD.n1313 VDD.n1208 4.5005
R78170 VDD.n1379 VDD.n1208 4.5005
R78171 VDD.n1312 VDD.n1208 4.5005
R78172 VDD.n1380 VDD.n1208 4.5005
R78173 VDD.n1310 VDD.n1208 4.5005
R78174 VDD.n1381 VDD.n1208 4.5005
R78175 VDD.n1309 VDD.n1208 4.5005
R78176 VDD.n1382 VDD.n1208 4.5005
R78177 VDD.n1307 VDD.n1208 4.5005
R78178 VDD.n1383 VDD.n1208 4.5005
R78179 VDD.n1306 VDD.n1208 4.5005
R78180 VDD.n1384 VDD.n1208 4.5005
R78181 VDD.n1304 VDD.n1208 4.5005
R78182 VDD.n1385 VDD.n1208 4.5005
R78183 VDD.n1303 VDD.n1208 4.5005
R78184 VDD.n1386 VDD.n1208 4.5005
R78185 VDD.n1301 VDD.n1208 4.5005
R78186 VDD.n1387 VDD.n1208 4.5005
R78187 VDD.n1300 VDD.n1208 4.5005
R78188 VDD.n1388 VDD.n1208 4.5005
R78189 VDD.n1298 VDD.n1208 4.5005
R78190 VDD.n1389 VDD.n1208 4.5005
R78191 VDD.n1297 VDD.n1208 4.5005
R78192 VDD.n1390 VDD.n1208 4.5005
R78193 VDD.n1295 VDD.n1208 4.5005
R78194 VDD.n1391 VDD.n1208 4.5005
R78195 VDD.n1294 VDD.n1208 4.5005
R78196 VDD.n1392 VDD.n1208 4.5005
R78197 VDD.n1292 VDD.n1208 4.5005
R78198 VDD.n1393 VDD.n1208 4.5005
R78199 VDD.n1291 VDD.n1208 4.5005
R78200 VDD.n1394 VDD.n1208 4.5005
R78201 VDD.n1289 VDD.n1208 4.5005
R78202 VDD.n1395 VDD.n1208 4.5005
R78203 VDD.n1288 VDD.n1208 4.5005
R78204 VDD.n1396 VDD.n1208 4.5005
R78205 VDD.n1286 VDD.n1208 4.5005
R78206 VDD.n1397 VDD.n1208 4.5005
R78207 VDD.n1285 VDD.n1208 4.5005
R78208 VDD.n1398 VDD.n1208 4.5005
R78209 VDD.n1283 VDD.n1208 4.5005
R78210 VDD.n1399 VDD.n1208 4.5005
R78211 VDD.n1282 VDD.n1208 4.5005
R78212 VDD.n1400 VDD.n1208 4.5005
R78213 VDD.n1280 VDD.n1208 4.5005
R78214 VDD.n1401 VDD.n1208 4.5005
R78215 VDD.n1279 VDD.n1208 4.5005
R78216 VDD.n1402 VDD.n1208 4.5005
R78217 VDD.n1277 VDD.n1208 4.5005
R78218 VDD.n1403 VDD.n1208 4.5005
R78219 VDD.n1276 VDD.n1208 4.5005
R78220 VDD.n1404 VDD.n1208 4.5005
R78221 VDD.n1274 VDD.n1208 4.5005
R78222 VDD.n1405 VDD.n1208 4.5005
R78223 VDD.n1273 VDD.n1208 4.5005
R78224 VDD.n1406 VDD.n1208 4.5005
R78225 VDD.n1271 VDD.n1208 4.5005
R78226 VDD.n1407 VDD.n1208 4.5005
R78227 VDD.n1270 VDD.n1208 4.5005
R78228 VDD.n1408 VDD.n1208 4.5005
R78229 VDD.n1268 VDD.n1208 4.5005
R78230 VDD.n1409 VDD.n1208 4.5005
R78231 VDD.n1267 VDD.n1208 4.5005
R78232 VDD.n1410 VDD.n1208 4.5005
R78233 VDD.n1265 VDD.n1208 4.5005
R78234 VDD.n1411 VDD.n1208 4.5005
R78235 VDD.n1264 VDD.n1208 4.5005
R78236 VDD.n1412 VDD.n1208 4.5005
R78237 VDD.n1262 VDD.n1208 4.5005
R78238 VDD.n1413 VDD.n1208 4.5005
R78239 VDD.n1261 VDD.n1208 4.5005
R78240 VDD.n1414 VDD.n1208 4.5005
R78241 VDD.n1415 VDD.n1208 4.5005
R78242 VDD.n1674 VDD.n1208 4.5005
R78243 VDD.n1676 VDD.n1181 4.5005
R78244 VDD.n1341 VDD.n1181 4.5005
R78245 VDD.n1342 VDD.n1181 4.5005
R78246 VDD.n1340 VDD.n1181 4.5005
R78247 VDD.n1344 VDD.n1181 4.5005
R78248 VDD.n1339 VDD.n1181 4.5005
R78249 VDD.n1345 VDD.n1181 4.5005
R78250 VDD.n1338 VDD.n1181 4.5005
R78251 VDD.n1347 VDD.n1181 4.5005
R78252 VDD.n1337 VDD.n1181 4.5005
R78253 VDD.n1348 VDD.n1181 4.5005
R78254 VDD.n1336 VDD.n1181 4.5005
R78255 VDD.n1350 VDD.n1181 4.5005
R78256 VDD.n1335 VDD.n1181 4.5005
R78257 VDD.n1351 VDD.n1181 4.5005
R78258 VDD.n1334 VDD.n1181 4.5005
R78259 VDD.n1353 VDD.n1181 4.5005
R78260 VDD.n1333 VDD.n1181 4.5005
R78261 VDD.n1354 VDD.n1181 4.5005
R78262 VDD.n1332 VDD.n1181 4.5005
R78263 VDD.n1356 VDD.n1181 4.5005
R78264 VDD.n1331 VDD.n1181 4.5005
R78265 VDD.n1357 VDD.n1181 4.5005
R78266 VDD.n1330 VDD.n1181 4.5005
R78267 VDD.n1359 VDD.n1181 4.5005
R78268 VDD.n1329 VDD.n1181 4.5005
R78269 VDD.n1360 VDD.n1181 4.5005
R78270 VDD.n1328 VDD.n1181 4.5005
R78271 VDD.n1362 VDD.n1181 4.5005
R78272 VDD.n1327 VDD.n1181 4.5005
R78273 VDD.n1363 VDD.n1181 4.5005
R78274 VDD.n1326 VDD.n1181 4.5005
R78275 VDD.n1365 VDD.n1181 4.5005
R78276 VDD.n1325 VDD.n1181 4.5005
R78277 VDD.n1366 VDD.n1181 4.5005
R78278 VDD.n1324 VDD.n1181 4.5005
R78279 VDD.n1368 VDD.n1181 4.5005
R78280 VDD.n1323 VDD.n1181 4.5005
R78281 VDD.n1369 VDD.n1181 4.5005
R78282 VDD.n1322 VDD.n1181 4.5005
R78283 VDD.n1371 VDD.n1181 4.5005
R78284 VDD.n1321 VDD.n1181 4.5005
R78285 VDD.n1372 VDD.n1181 4.5005
R78286 VDD.n1320 VDD.n1181 4.5005
R78287 VDD.n1374 VDD.n1181 4.5005
R78288 VDD.n1319 VDD.n1181 4.5005
R78289 VDD.n1375 VDD.n1181 4.5005
R78290 VDD.n1318 VDD.n1181 4.5005
R78291 VDD.n1376 VDD.n1181 4.5005
R78292 VDD.n1316 VDD.n1181 4.5005
R78293 VDD.n1377 VDD.n1181 4.5005
R78294 VDD.n1315 VDD.n1181 4.5005
R78295 VDD.n1378 VDD.n1181 4.5005
R78296 VDD.n1313 VDD.n1181 4.5005
R78297 VDD.n1379 VDD.n1181 4.5005
R78298 VDD.n1312 VDD.n1181 4.5005
R78299 VDD.n1380 VDD.n1181 4.5005
R78300 VDD.n1310 VDD.n1181 4.5005
R78301 VDD.n1381 VDD.n1181 4.5005
R78302 VDD.n1309 VDD.n1181 4.5005
R78303 VDD.n1382 VDD.n1181 4.5005
R78304 VDD.n1307 VDD.n1181 4.5005
R78305 VDD.n1383 VDD.n1181 4.5005
R78306 VDD.n1306 VDD.n1181 4.5005
R78307 VDD.n1384 VDD.n1181 4.5005
R78308 VDD.n1304 VDD.n1181 4.5005
R78309 VDD.n1385 VDD.n1181 4.5005
R78310 VDD.n1303 VDD.n1181 4.5005
R78311 VDD.n1386 VDD.n1181 4.5005
R78312 VDD.n1301 VDD.n1181 4.5005
R78313 VDD.n1387 VDD.n1181 4.5005
R78314 VDD.n1300 VDD.n1181 4.5005
R78315 VDD.n1388 VDD.n1181 4.5005
R78316 VDD.n1298 VDD.n1181 4.5005
R78317 VDD.n1389 VDD.n1181 4.5005
R78318 VDD.n1297 VDD.n1181 4.5005
R78319 VDD.n1390 VDD.n1181 4.5005
R78320 VDD.n1295 VDD.n1181 4.5005
R78321 VDD.n1391 VDD.n1181 4.5005
R78322 VDD.n1294 VDD.n1181 4.5005
R78323 VDD.n1392 VDD.n1181 4.5005
R78324 VDD.n1292 VDD.n1181 4.5005
R78325 VDD.n1393 VDD.n1181 4.5005
R78326 VDD.n1291 VDD.n1181 4.5005
R78327 VDD.n1394 VDD.n1181 4.5005
R78328 VDD.n1289 VDD.n1181 4.5005
R78329 VDD.n1395 VDD.n1181 4.5005
R78330 VDD.n1288 VDD.n1181 4.5005
R78331 VDD.n1396 VDD.n1181 4.5005
R78332 VDD.n1286 VDD.n1181 4.5005
R78333 VDD.n1397 VDD.n1181 4.5005
R78334 VDD.n1285 VDD.n1181 4.5005
R78335 VDD.n1398 VDD.n1181 4.5005
R78336 VDD.n1283 VDD.n1181 4.5005
R78337 VDD.n1399 VDD.n1181 4.5005
R78338 VDD.n1282 VDD.n1181 4.5005
R78339 VDD.n1400 VDD.n1181 4.5005
R78340 VDD.n1280 VDD.n1181 4.5005
R78341 VDD.n1401 VDD.n1181 4.5005
R78342 VDD.n1279 VDD.n1181 4.5005
R78343 VDD.n1402 VDD.n1181 4.5005
R78344 VDD.n1277 VDD.n1181 4.5005
R78345 VDD.n1403 VDD.n1181 4.5005
R78346 VDD.n1276 VDD.n1181 4.5005
R78347 VDD.n1404 VDD.n1181 4.5005
R78348 VDD.n1274 VDD.n1181 4.5005
R78349 VDD.n1405 VDD.n1181 4.5005
R78350 VDD.n1273 VDD.n1181 4.5005
R78351 VDD.n1406 VDD.n1181 4.5005
R78352 VDD.n1271 VDD.n1181 4.5005
R78353 VDD.n1407 VDD.n1181 4.5005
R78354 VDD.n1270 VDD.n1181 4.5005
R78355 VDD.n1408 VDD.n1181 4.5005
R78356 VDD.n1268 VDD.n1181 4.5005
R78357 VDD.n1409 VDD.n1181 4.5005
R78358 VDD.n1267 VDD.n1181 4.5005
R78359 VDD.n1410 VDD.n1181 4.5005
R78360 VDD.n1265 VDD.n1181 4.5005
R78361 VDD.n1411 VDD.n1181 4.5005
R78362 VDD.n1264 VDD.n1181 4.5005
R78363 VDD.n1412 VDD.n1181 4.5005
R78364 VDD.n1262 VDD.n1181 4.5005
R78365 VDD.n1413 VDD.n1181 4.5005
R78366 VDD.n1261 VDD.n1181 4.5005
R78367 VDD.n1414 VDD.n1181 4.5005
R78368 VDD.n1415 VDD.n1181 4.5005
R78369 VDD.n1674 VDD.n1181 4.5005
R78370 VDD.n1676 VDD.n1209 4.5005
R78371 VDD.n1341 VDD.n1209 4.5005
R78372 VDD.n1342 VDD.n1209 4.5005
R78373 VDD.n1340 VDD.n1209 4.5005
R78374 VDD.n1344 VDD.n1209 4.5005
R78375 VDD.n1339 VDD.n1209 4.5005
R78376 VDD.n1345 VDD.n1209 4.5005
R78377 VDD.n1338 VDD.n1209 4.5005
R78378 VDD.n1347 VDD.n1209 4.5005
R78379 VDD.n1337 VDD.n1209 4.5005
R78380 VDD.n1348 VDD.n1209 4.5005
R78381 VDD.n1336 VDD.n1209 4.5005
R78382 VDD.n1350 VDD.n1209 4.5005
R78383 VDD.n1335 VDD.n1209 4.5005
R78384 VDD.n1351 VDD.n1209 4.5005
R78385 VDD.n1334 VDD.n1209 4.5005
R78386 VDD.n1353 VDD.n1209 4.5005
R78387 VDD.n1333 VDD.n1209 4.5005
R78388 VDD.n1354 VDD.n1209 4.5005
R78389 VDD.n1332 VDD.n1209 4.5005
R78390 VDD.n1356 VDD.n1209 4.5005
R78391 VDD.n1331 VDD.n1209 4.5005
R78392 VDD.n1357 VDD.n1209 4.5005
R78393 VDD.n1330 VDD.n1209 4.5005
R78394 VDD.n1359 VDD.n1209 4.5005
R78395 VDD.n1329 VDD.n1209 4.5005
R78396 VDD.n1360 VDD.n1209 4.5005
R78397 VDD.n1328 VDD.n1209 4.5005
R78398 VDD.n1362 VDD.n1209 4.5005
R78399 VDD.n1327 VDD.n1209 4.5005
R78400 VDD.n1363 VDD.n1209 4.5005
R78401 VDD.n1326 VDD.n1209 4.5005
R78402 VDD.n1365 VDD.n1209 4.5005
R78403 VDD.n1325 VDD.n1209 4.5005
R78404 VDD.n1366 VDD.n1209 4.5005
R78405 VDD.n1324 VDD.n1209 4.5005
R78406 VDD.n1368 VDD.n1209 4.5005
R78407 VDD.n1323 VDD.n1209 4.5005
R78408 VDD.n1369 VDD.n1209 4.5005
R78409 VDD.n1322 VDD.n1209 4.5005
R78410 VDD.n1371 VDD.n1209 4.5005
R78411 VDD.n1321 VDD.n1209 4.5005
R78412 VDD.n1372 VDD.n1209 4.5005
R78413 VDD.n1320 VDD.n1209 4.5005
R78414 VDD.n1374 VDD.n1209 4.5005
R78415 VDD.n1319 VDD.n1209 4.5005
R78416 VDD.n1375 VDD.n1209 4.5005
R78417 VDD.n1318 VDD.n1209 4.5005
R78418 VDD.n1376 VDD.n1209 4.5005
R78419 VDD.n1316 VDD.n1209 4.5005
R78420 VDD.n1377 VDD.n1209 4.5005
R78421 VDD.n1315 VDD.n1209 4.5005
R78422 VDD.n1378 VDD.n1209 4.5005
R78423 VDD.n1313 VDD.n1209 4.5005
R78424 VDD.n1379 VDD.n1209 4.5005
R78425 VDD.n1312 VDD.n1209 4.5005
R78426 VDD.n1380 VDD.n1209 4.5005
R78427 VDD.n1310 VDD.n1209 4.5005
R78428 VDD.n1381 VDD.n1209 4.5005
R78429 VDD.n1309 VDD.n1209 4.5005
R78430 VDD.n1382 VDD.n1209 4.5005
R78431 VDD.n1307 VDD.n1209 4.5005
R78432 VDD.n1383 VDD.n1209 4.5005
R78433 VDD.n1306 VDD.n1209 4.5005
R78434 VDD.n1384 VDD.n1209 4.5005
R78435 VDD.n1304 VDD.n1209 4.5005
R78436 VDD.n1385 VDD.n1209 4.5005
R78437 VDD.n1303 VDD.n1209 4.5005
R78438 VDD.n1386 VDD.n1209 4.5005
R78439 VDD.n1301 VDD.n1209 4.5005
R78440 VDD.n1387 VDD.n1209 4.5005
R78441 VDD.n1300 VDD.n1209 4.5005
R78442 VDD.n1388 VDD.n1209 4.5005
R78443 VDD.n1298 VDD.n1209 4.5005
R78444 VDD.n1389 VDD.n1209 4.5005
R78445 VDD.n1297 VDD.n1209 4.5005
R78446 VDD.n1390 VDD.n1209 4.5005
R78447 VDD.n1295 VDD.n1209 4.5005
R78448 VDD.n1391 VDD.n1209 4.5005
R78449 VDD.n1294 VDD.n1209 4.5005
R78450 VDD.n1392 VDD.n1209 4.5005
R78451 VDD.n1292 VDD.n1209 4.5005
R78452 VDD.n1393 VDD.n1209 4.5005
R78453 VDD.n1291 VDD.n1209 4.5005
R78454 VDD.n1394 VDD.n1209 4.5005
R78455 VDD.n1289 VDD.n1209 4.5005
R78456 VDD.n1395 VDD.n1209 4.5005
R78457 VDD.n1288 VDD.n1209 4.5005
R78458 VDD.n1396 VDD.n1209 4.5005
R78459 VDD.n1286 VDD.n1209 4.5005
R78460 VDD.n1397 VDD.n1209 4.5005
R78461 VDD.n1285 VDD.n1209 4.5005
R78462 VDD.n1398 VDD.n1209 4.5005
R78463 VDD.n1283 VDD.n1209 4.5005
R78464 VDD.n1399 VDD.n1209 4.5005
R78465 VDD.n1282 VDD.n1209 4.5005
R78466 VDD.n1400 VDD.n1209 4.5005
R78467 VDD.n1280 VDD.n1209 4.5005
R78468 VDD.n1401 VDD.n1209 4.5005
R78469 VDD.n1279 VDD.n1209 4.5005
R78470 VDD.n1402 VDD.n1209 4.5005
R78471 VDD.n1277 VDD.n1209 4.5005
R78472 VDD.n1403 VDD.n1209 4.5005
R78473 VDD.n1276 VDD.n1209 4.5005
R78474 VDD.n1404 VDD.n1209 4.5005
R78475 VDD.n1274 VDD.n1209 4.5005
R78476 VDD.n1405 VDD.n1209 4.5005
R78477 VDD.n1273 VDD.n1209 4.5005
R78478 VDD.n1406 VDD.n1209 4.5005
R78479 VDD.n1271 VDD.n1209 4.5005
R78480 VDD.n1407 VDD.n1209 4.5005
R78481 VDD.n1270 VDD.n1209 4.5005
R78482 VDD.n1408 VDD.n1209 4.5005
R78483 VDD.n1268 VDD.n1209 4.5005
R78484 VDD.n1409 VDD.n1209 4.5005
R78485 VDD.n1267 VDD.n1209 4.5005
R78486 VDD.n1410 VDD.n1209 4.5005
R78487 VDD.n1265 VDD.n1209 4.5005
R78488 VDD.n1411 VDD.n1209 4.5005
R78489 VDD.n1264 VDD.n1209 4.5005
R78490 VDD.n1412 VDD.n1209 4.5005
R78491 VDD.n1262 VDD.n1209 4.5005
R78492 VDD.n1413 VDD.n1209 4.5005
R78493 VDD.n1261 VDD.n1209 4.5005
R78494 VDD.n1414 VDD.n1209 4.5005
R78495 VDD.n1415 VDD.n1209 4.5005
R78496 VDD.n1674 VDD.n1209 4.5005
R78497 VDD.n1676 VDD.n1180 4.5005
R78498 VDD.n1341 VDD.n1180 4.5005
R78499 VDD.n1342 VDD.n1180 4.5005
R78500 VDD.n1340 VDD.n1180 4.5005
R78501 VDD.n1344 VDD.n1180 4.5005
R78502 VDD.n1339 VDD.n1180 4.5005
R78503 VDD.n1345 VDD.n1180 4.5005
R78504 VDD.n1338 VDD.n1180 4.5005
R78505 VDD.n1347 VDD.n1180 4.5005
R78506 VDD.n1337 VDD.n1180 4.5005
R78507 VDD.n1348 VDD.n1180 4.5005
R78508 VDD.n1336 VDD.n1180 4.5005
R78509 VDD.n1350 VDD.n1180 4.5005
R78510 VDD.n1335 VDD.n1180 4.5005
R78511 VDD.n1351 VDD.n1180 4.5005
R78512 VDD.n1334 VDD.n1180 4.5005
R78513 VDD.n1353 VDD.n1180 4.5005
R78514 VDD.n1333 VDD.n1180 4.5005
R78515 VDD.n1354 VDD.n1180 4.5005
R78516 VDD.n1332 VDD.n1180 4.5005
R78517 VDD.n1356 VDD.n1180 4.5005
R78518 VDD.n1331 VDD.n1180 4.5005
R78519 VDD.n1357 VDD.n1180 4.5005
R78520 VDD.n1330 VDD.n1180 4.5005
R78521 VDD.n1359 VDD.n1180 4.5005
R78522 VDD.n1329 VDD.n1180 4.5005
R78523 VDD.n1360 VDD.n1180 4.5005
R78524 VDD.n1328 VDD.n1180 4.5005
R78525 VDD.n1362 VDD.n1180 4.5005
R78526 VDD.n1327 VDD.n1180 4.5005
R78527 VDD.n1363 VDD.n1180 4.5005
R78528 VDD.n1326 VDD.n1180 4.5005
R78529 VDD.n1365 VDD.n1180 4.5005
R78530 VDD.n1325 VDD.n1180 4.5005
R78531 VDD.n1366 VDD.n1180 4.5005
R78532 VDD.n1324 VDD.n1180 4.5005
R78533 VDD.n1368 VDD.n1180 4.5005
R78534 VDD.n1323 VDD.n1180 4.5005
R78535 VDD.n1369 VDD.n1180 4.5005
R78536 VDD.n1322 VDD.n1180 4.5005
R78537 VDD.n1371 VDD.n1180 4.5005
R78538 VDD.n1321 VDD.n1180 4.5005
R78539 VDD.n1372 VDD.n1180 4.5005
R78540 VDD.n1320 VDD.n1180 4.5005
R78541 VDD.n1374 VDD.n1180 4.5005
R78542 VDD.n1319 VDD.n1180 4.5005
R78543 VDD.n1375 VDD.n1180 4.5005
R78544 VDD.n1318 VDD.n1180 4.5005
R78545 VDD.n1376 VDD.n1180 4.5005
R78546 VDD.n1316 VDD.n1180 4.5005
R78547 VDD.n1377 VDD.n1180 4.5005
R78548 VDD.n1315 VDD.n1180 4.5005
R78549 VDD.n1378 VDD.n1180 4.5005
R78550 VDD.n1313 VDD.n1180 4.5005
R78551 VDD.n1379 VDD.n1180 4.5005
R78552 VDD.n1312 VDD.n1180 4.5005
R78553 VDD.n1380 VDD.n1180 4.5005
R78554 VDD.n1310 VDD.n1180 4.5005
R78555 VDD.n1381 VDD.n1180 4.5005
R78556 VDD.n1309 VDD.n1180 4.5005
R78557 VDD.n1382 VDD.n1180 4.5005
R78558 VDD.n1307 VDD.n1180 4.5005
R78559 VDD.n1383 VDD.n1180 4.5005
R78560 VDD.n1306 VDD.n1180 4.5005
R78561 VDD.n1384 VDD.n1180 4.5005
R78562 VDD.n1304 VDD.n1180 4.5005
R78563 VDD.n1385 VDD.n1180 4.5005
R78564 VDD.n1303 VDD.n1180 4.5005
R78565 VDD.n1386 VDD.n1180 4.5005
R78566 VDD.n1301 VDD.n1180 4.5005
R78567 VDD.n1387 VDD.n1180 4.5005
R78568 VDD.n1300 VDD.n1180 4.5005
R78569 VDD.n1388 VDD.n1180 4.5005
R78570 VDD.n1298 VDD.n1180 4.5005
R78571 VDD.n1389 VDD.n1180 4.5005
R78572 VDD.n1297 VDD.n1180 4.5005
R78573 VDD.n1390 VDD.n1180 4.5005
R78574 VDD.n1295 VDD.n1180 4.5005
R78575 VDD.n1391 VDD.n1180 4.5005
R78576 VDD.n1294 VDD.n1180 4.5005
R78577 VDD.n1392 VDD.n1180 4.5005
R78578 VDD.n1292 VDD.n1180 4.5005
R78579 VDD.n1393 VDD.n1180 4.5005
R78580 VDD.n1291 VDD.n1180 4.5005
R78581 VDD.n1394 VDD.n1180 4.5005
R78582 VDD.n1289 VDD.n1180 4.5005
R78583 VDD.n1395 VDD.n1180 4.5005
R78584 VDD.n1288 VDD.n1180 4.5005
R78585 VDD.n1396 VDD.n1180 4.5005
R78586 VDD.n1286 VDD.n1180 4.5005
R78587 VDD.n1397 VDD.n1180 4.5005
R78588 VDD.n1285 VDD.n1180 4.5005
R78589 VDD.n1398 VDD.n1180 4.5005
R78590 VDD.n1283 VDD.n1180 4.5005
R78591 VDD.n1399 VDD.n1180 4.5005
R78592 VDD.n1282 VDD.n1180 4.5005
R78593 VDD.n1400 VDD.n1180 4.5005
R78594 VDD.n1280 VDD.n1180 4.5005
R78595 VDD.n1401 VDD.n1180 4.5005
R78596 VDD.n1279 VDD.n1180 4.5005
R78597 VDD.n1402 VDD.n1180 4.5005
R78598 VDD.n1277 VDD.n1180 4.5005
R78599 VDD.n1403 VDD.n1180 4.5005
R78600 VDD.n1276 VDD.n1180 4.5005
R78601 VDD.n1404 VDD.n1180 4.5005
R78602 VDD.n1274 VDD.n1180 4.5005
R78603 VDD.n1405 VDD.n1180 4.5005
R78604 VDD.n1273 VDD.n1180 4.5005
R78605 VDD.n1406 VDD.n1180 4.5005
R78606 VDD.n1271 VDD.n1180 4.5005
R78607 VDD.n1407 VDD.n1180 4.5005
R78608 VDD.n1270 VDD.n1180 4.5005
R78609 VDD.n1408 VDD.n1180 4.5005
R78610 VDD.n1268 VDD.n1180 4.5005
R78611 VDD.n1409 VDD.n1180 4.5005
R78612 VDD.n1267 VDD.n1180 4.5005
R78613 VDD.n1410 VDD.n1180 4.5005
R78614 VDD.n1265 VDD.n1180 4.5005
R78615 VDD.n1411 VDD.n1180 4.5005
R78616 VDD.n1264 VDD.n1180 4.5005
R78617 VDD.n1412 VDD.n1180 4.5005
R78618 VDD.n1262 VDD.n1180 4.5005
R78619 VDD.n1413 VDD.n1180 4.5005
R78620 VDD.n1261 VDD.n1180 4.5005
R78621 VDD.n1414 VDD.n1180 4.5005
R78622 VDD.n1415 VDD.n1180 4.5005
R78623 VDD.n1674 VDD.n1180 4.5005
R78624 VDD.n1676 VDD.n1210 4.5005
R78625 VDD.n1341 VDD.n1210 4.5005
R78626 VDD.n1342 VDD.n1210 4.5005
R78627 VDD.n1340 VDD.n1210 4.5005
R78628 VDD.n1344 VDD.n1210 4.5005
R78629 VDD.n1339 VDD.n1210 4.5005
R78630 VDD.n1345 VDD.n1210 4.5005
R78631 VDD.n1338 VDD.n1210 4.5005
R78632 VDD.n1347 VDD.n1210 4.5005
R78633 VDD.n1337 VDD.n1210 4.5005
R78634 VDD.n1348 VDD.n1210 4.5005
R78635 VDD.n1336 VDD.n1210 4.5005
R78636 VDD.n1350 VDD.n1210 4.5005
R78637 VDD.n1335 VDD.n1210 4.5005
R78638 VDD.n1351 VDD.n1210 4.5005
R78639 VDD.n1334 VDD.n1210 4.5005
R78640 VDD.n1353 VDD.n1210 4.5005
R78641 VDD.n1333 VDD.n1210 4.5005
R78642 VDD.n1354 VDD.n1210 4.5005
R78643 VDD.n1332 VDD.n1210 4.5005
R78644 VDD.n1356 VDD.n1210 4.5005
R78645 VDD.n1331 VDD.n1210 4.5005
R78646 VDD.n1357 VDD.n1210 4.5005
R78647 VDD.n1330 VDD.n1210 4.5005
R78648 VDD.n1359 VDD.n1210 4.5005
R78649 VDD.n1329 VDD.n1210 4.5005
R78650 VDD.n1360 VDD.n1210 4.5005
R78651 VDD.n1328 VDD.n1210 4.5005
R78652 VDD.n1362 VDD.n1210 4.5005
R78653 VDD.n1327 VDD.n1210 4.5005
R78654 VDD.n1363 VDD.n1210 4.5005
R78655 VDD.n1326 VDD.n1210 4.5005
R78656 VDD.n1365 VDD.n1210 4.5005
R78657 VDD.n1325 VDD.n1210 4.5005
R78658 VDD.n1366 VDD.n1210 4.5005
R78659 VDD.n1324 VDD.n1210 4.5005
R78660 VDD.n1368 VDD.n1210 4.5005
R78661 VDD.n1323 VDD.n1210 4.5005
R78662 VDD.n1369 VDD.n1210 4.5005
R78663 VDD.n1322 VDD.n1210 4.5005
R78664 VDD.n1371 VDD.n1210 4.5005
R78665 VDD.n1321 VDD.n1210 4.5005
R78666 VDD.n1372 VDD.n1210 4.5005
R78667 VDD.n1320 VDD.n1210 4.5005
R78668 VDD.n1374 VDD.n1210 4.5005
R78669 VDD.n1319 VDD.n1210 4.5005
R78670 VDD.n1375 VDD.n1210 4.5005
R78671 VDD.n1318 VDD.n1210 4.5005
R78672 VDD.n1376 VDD.n1210 4.5005
R78673 VDD.n1316 VDD.n1210 4.5005
R78674 VDD.n1377 VDD.n1210 4.5005
R78675 VDD.n1315 VDD.n1210 4.5005
R78676 VDD.n1378 VDD.n1210 4.5005
R78677 VDD.n1313 VDD.n1210 4.5005
R78678 VDD.n1379 VDD.n1210 4.5005
R78679 VDD.n1312 VDD.n1210 4.5005
R78680 VDD.n1380 VDD.n1210 4.5005
R78681 VDD.n1310 VDD.n1210 4.5005
R78682 VDD.n1381 VDD.n1210 4.5005
R78683 VDD.n1309 VDD.n1210 4.5005
R78684 VDD.n1382 VDD.n1210 4.5005
R78685 VDD.n1307 VDD.n1210 4.5005
R78686 VDD.n1383 VDD.n1210 4.5005
R78687 VDD.n1306 VDD.n1210 4.5005
R78688 VDD.n1384 VDD.n1210 4.5005
R78689 VDD.n1304 VDD.n1210 4.5005
R78690 VDD.n1385 VDD.n1210 4.5005
R78691 VDD.n1303 VDD.n1210 4.5005
R78692 VDD.n1386 VDD.n1210 4.5005
R78693 VDD.n1301 VDD.n1210 4.5005
R78694 VDD.n1387 VDD.n1210 4.5005
R78695 VDD.n1300 VDD.n1210 4.5005
R78696 VDD.n1388 VDD.n1210 4.5005
R78697 VDD.n1298 VDD.n1210 4.5005
R78698 VDD.n1389 VDD.n1210 4.5005
R78699 VDD.n1297 VDD.n1210 4.5005
R78700 VDD.n1390 VDD.n1210 4.5005
R78701 VDD.n1295 VDD.n1210 4.5005
R78702 VDD.n1391 VDD.n1210 4.5005
R78703 VDD.n1294 VDD.n1210 4.5005
R78704 VDD.n1392 VDD.n1210 4.5005
R78705 VDD.n1292 VDD.n1210 4.5005
R78706 VDD.n1393 VDD.n1210 4.5005
R78707 VDD.n1291 VDD.n1210 4.5005
R78708 VDD.n1394 VDD.n1210 4.5005
R78709 VDD.n1289 VDD.n1210 4.5005
R78710 VDD.n1395 VDD.n1210 4.5005
R78711 VDD.n1288 VDD.n1210 4.5005
R78712 VDD.n1396 VDD.n1210 4.5005
R78713 VDD.n1286 VDD.n1210 4.5005
R78714 VDD.n1397 VDD.n1210 4.5005
R78715 VDD.n1285 VDD.n1210 4.5005
R78716 VDD.n1398 VDD.n1210 4.5005
R78717 VDD.n1283 VDD.n1210 4.5005
R78718 VDD.n1399 VDD.n1210 4.5005
R78719 VDD.n1282 VDD.n1210 4.5005
R78720 VDD.n1400 VDD.n1210 4.5005
R78721 VDD.n1280 VDD.n1210 4.5005
R78722 VDD.n1401 VDD.n1210 4.5005
R78723 VDD.n1279 VDD.n1210 4.5005
R78724 VDD.n1402 VDD.n1210 4.5005
R78725 VDD.n1277 VDD.n1210 4.5005
R78726 VDD.n1403 VDD.n1210 4.5005
R78727 VDD.n1276 VDD.n1210 4.5005
R78728 VDD.n1404 VDD.n1210 4.5005
R78729 VDD.n1274 VDD.n1210 4.5005
R78730 VDD.n1405 VDD.n1210 4.5005
R78731 VDD.n1273 VDD.n1210 4.5005
R78732 VDD.n1406 VDD.n1210 4.5005
R78733 VDD.n1271 VDD.n1210 4.5005
R78734 VDD.n1407 VDD.n1210 4.5005
R78735 VDD.n1270 VDD.n1210 4.5005
R78736 VDD.n1408 VDD.n1210 4.5005
R78737 VDD.n1268 VDD.n1210 4.5005
R78738 VDD.n1409 VDD.n1210 4.5005
R78739 VDD.n1267 VDD.n1210 4.5005
R78740 VDD.n1410 VDD.n1210 4.5005
R78741 VDD.n1265 VDD.n1210 4.5005
R78742 VDD.n1411 VDD.n1210 4.5005
R78743 VDD.n1264 VDD.n1210 4.5005
R78744 VDD.n1412 VDD.n1210 4.5005
R78745 VDD.n1262 VDD.n1210 4.5005
R78746 VDD.n1413 VDD.n1210 4.5005
R78747 VDD.n1261 VDD.n1210 4.5005
R78748 VDD.n1414 VDD.n1210 4.5005
R78749 VDD.n1415 VDD.n1210 4.5005
R78750 VDD.n1674 VDD.n1210 4.5005
R78751 VDD.n1676 VDD.n1179 4.5005
R78752 VDD.n1341 VDD.n1179 4.5005
R78753 VDD.n1342 VDD.n1179 4.5005
R78754 VDD.n1340 VDD.n1179 4.5005
R78755 VDD.n1344 VDD.n1179 4.5005
R78756 VDD.n1339 VDD.n1179 4.5005
R78757 VDD.n1345 VDD.n1179 4.5005
R78758 VDD.n1338 VDD.n1179 4.5005
R78759 VDD.n1347 VDD.n1179 4.5005
R78760 VDD.n1337 VDD.n1179 4.5005
R78761 VDD.n1348 VDD.n1179 4.5005
R78762 VDD.n1336 VDD.n1179 4.5005
R78763 VDD.n1350 VDD.n1179 4.5005
R78764 VDD.n1335 VDD.n1179 4.5005
R78765 VDD.n1351 VDD.n1179 4.5005
R78766 VDD.n1334 VDD.n1179 4.5005
R78767 VDD.n1353 VDD.n1179 4.5005
R78768 VDD.n1333 VDD.n1179 4.5005
R78769 VDD.n1354 VDD.n1179 4.5005
R78770 VDD.n1332 VDD.n1179 4.5005
R78771 VDD.n1356 VDD.n1179 4.5005
R78772 VDD.n1331 VDD.n1179 4.5005
R78773 VDD.n1357 VDD.n1179 4.5005
R78774 VDD.n1330 VDD.n1179 4.5005
R78775 VDD.n1359 VDD.n1179 4.5005
R78776 VDD.n1329 VDD.n1179 4.5005
R78777 VDD.n1360 VDD.n1179 4.5005
R78778 VDD.n1328 VDD.n1179 4.5005
R78779 VDD.n1362 VDD.n1179 4.5005
R78780 VDD.n1327 VDD.n1179 4.5005
R78781 VDD.n1363 VDD.n1179 4.5005
R78782 VDD.n1326 VDD.n1179 4.5005
R78783 VDD.n1365 VDD.n1179 4.5005
R78784 VDD.n1325 VDD.n1179 4.5005
R78785 VDD.n1366 VDD.n1179 4.5005
R78786 VDD.n1324 VDD.n1179 4.5005
R78787 VDD.n1368 VDD.n1179 4.5005
R78788 VDD.n1323 VDD.n1179 4.5005
R78789 VDD.n1369 VDD.n1179 4.5005
R78790 VDD.n1322 VDD.n1179 4.5005
R78791 VDD.n1371 VDD.n1179 4.5005
R78792 VDD.n1321 VDD.n1179 4.5005
R78793 VDD.n1372 VDD.n1179 4.5005
R78794 VDD.n1320 VDD.n1179 4.5005
R78795 VDD.n1374 VDD.n1179 4.5005
R78796 VDD.n1319 VDD.n1179 4.5005
R78797 VDD.n1375 VDD.n1179 4.5005
R78798 VDD.n1318 VDD.n1179 4.5005
R78799 VDD.n1376 VDD.n1179 4.5005
R78800 VDD.n1316 VDD.n1179 4.5005
R78801 VDD.n1377 VDD.n1179 4.5005
R78802 VDD.n1315 VDD.n1179 4.5005
R78803 VDD.n1378 VDD.n1179 4.5005
R78804 VDD.n1313 VDD.n1179 4.5005
R78805 VDD.n1379 VDD.n1179 4.5005
R78806 VDD.n1312 VDD.n1179 4.5005
R78807 VDD.n1380 VDD.n1179 4.5005
R78808 VDD.n1310 VDD.n1179 4.5005
R78809 VDD.n1381 VDD.n1179 4.5005
R78810 VDD.n1309 VDD.n1179 4.5005
R78811 VDD.n1382 VDD.n1179 4.5005
R78812 VDD.n1307 VDD.n1179 4.5005
R78813 VDD.n1383 VDD.n1179 4.5005
R78814 VDD.n1306 VDD.n1179 4.5005
R78815 VDD.n1384 VDD.n1179 4.5005
R78816 VDD.n1304 VDD.n1179 4.5005
R78817 VDD.n1385 VDD.n1179 4.5005
R78818 VDD.n1303 VDD.n1179 4.5005
R78819 VDD.n1386 VDD.n1179 4.5005
R78820 VDD.n1301 VDD.n1179 4.5005
R78821 VDD.n1387 VDD.n1179 4.5005
R78822 VDD.n1300 VDD.n1179 4.5005
R78823 VDD.n1388 VDD.n1179 4.5005
R78824 VDD.n1298 VDD.n1179 4.5005
R78825 VDD.n1389 VDD.n1179 4.5005
R78826 VDD.n1297 VDD.n1179 4.5005
R78827 VDD.n1390 VDD.n1179 4.5005
R78828 VDD.n1295 VDD.n1179 4.5005
R78829 VDD.n1391 VDD.n1179 4.5005
R78830 VDD.n1294 VDD.n1179 4.5005
R78831 VDD.n1392 VDD.n1179 4.5005
R78832 VDD.n1292 VDD.n1179 4.5005
R78833 VDD.n1393 VDD.n1179 4.5005
R78834 VDD.n1291 VDD.n1179 4.5005
R78835 VDD.n1394 VDD.n1179 4.5005
R78836 VDD.n1289 VDD.n1179 4.5005
R78837 VDD.n1395 VDD.n1179 4.5005
R78838 VDD.n1288 VDD.n1179 4.5005
R78839 VDD.n1396 VDD.n1179 4.5005
R78840 VDD.n1286 VDD.n1179 4.5005
R78841 VDD.n1397 VDD.n1179 4.5005
R78842 VDD.n1285 VDD.n1179 4.5005
R78843 VDD.n1398 VDD.n1179 4.5005
R78844 VDD.n1283 VDD.n1179 4.5005
R78845 VDD.n1399 VDD.n1179 4.5005
R78846 VDD.n1282 VDD.n1179 4.5005
R78847 VDD.n1400 VDD.n1179 4.5005
R78848 VDD.n1280 VDD.n1179 4.5005
R78849 VDD.n1401 VDD.n1179 4.5005
R78850 VDD.n1279 VDD.n1179 4.5005
R78851 VDD.n1402 VDD.n1179 4.5005
R78852 VDD.n1277 VDD.n1179 4.5005
R78853 VDD.n1403 VDD.n1179 4.5005
R78854 VDD.n1276 VDD.n1179 4.5005
R78855 VDD.n1404 VDD.n1179 4.5005
R78856 VDD.n1274 VDD.n1179 4.5005
R78857 VDD.n1405 VDD.n1179 4.5005
R78858 VDD.n1273 VDD.n1179 4.5005
R78859 VDD.n1406 VDD.n1179 4.5005
R78860 VDD.n1271 VDD.n1179 4.5005
R78861 VDD.n1407 VDD.n1179 4.5005
R78862 VDD.n1270 VDD.n1179 4.5005
R78863 VDD.n1408 VDD.n1179 4.5005
R78864 VDD.n1268 VDD.n1179 4.5005
R78865 VDD.n1409 VDD.n1179 4.5005
R78866 VDD.n1267 VDD.n1179 4.5005
R78867 VDD.n1410 VDD.n1179 4.5005
R78868 VDD.n1265 VDD.n1179 4.5005
R78869 VDD.n1411 VDD.n1179 4.5005
R78870 VDD.n1264 VDD.n1179 4.5005
R78871 VDD.n1412 VDD.n1179 4.5005
R78872 VDD.n1262 VDD.n1179 4.5005
R78873 VDD.n1413 VDD.n1179 4.5005
R78874 VDD.n1261 VDD.n1179 4.5005
R78875 VDD.n1414 VDD.n1179 4.5005
R78876 VDD.n1415 VDD.n1179 4.5005
R78877 VDD.n1674 VDD.n1179 4.5005
R78878 VDD.n1676 VDD.n1211 4.5005
R78879 VDD.n1341 VDD.n1211 4.5005
R78880 VDD.n1342 VDD.n1211 4.5005
R78881 VDD.n1340 VDD.n1211 4.5005
R78882 VDD.n1344 VDD.n1211 4.5005
R78883 VDD.n1339 VDD.n1211 4.5005
R78884 VDD.n1345 VDD.n1211 4.5005
R78885 VDD.n1338 VDD.n1211 4.5005
R78886 VDD.n1347 VDD.n1211 4.5005
R78887 VDD.n1337 VDD.n1211 4.5005
R78888 VDD.n1348 VDD.n1211 4.5005
R78889 VDD.n1336 VDD.n1211 4.5005
R78890 VDD.n1350 VDD.n1211 4.5005
R78891 VDD.n1335 VDD.n1211 4.5005
R78892 VDD.n1351 VDD.n1211 4.5005
R78893 VDD.n1334 VDD.n1211 4.5005
R78894 VDD.n1353 VDD.n1211 4.5005
R78895 VDD.n1333 VDD.n1211 4.5005
R78896 VDD.n1354 VDD.n1211 4.5005
R78897 VDD.n1332 VDD.n1211 4.5005
R78898 VDD.n1356 VDD.n1211 4.5005
R78899 VDD.n1331 VDD.n1211 4.5005
R78900 VDD.n1357 VDD.n1211 4.5005
R78901 VDD.n1330 VDD.n1211 4.5005
R78902 VDD.n1359 VDD.n1211 4.5005
R78903 VDD.n1329 VDD.n1211 4.5005
R78904 VDD.n1360 VDD.n1211 4.5005
R78905 VDD.n1328 VDD.n1211 4.5005
R78906 VDD.n1362 VDD.n1211 4.5005
R78907 VDD.n1327 VDD.n1211 4.5005
R78908 VDD.n1363 VDD.n1211 4.5005
R78909 VDD.n1326 VDD.n1211 4.5005
R78910 VDD.n1365 VDD.n1211 4.5005
R78911 VDD.n1325 VDD.n1211 4.5005
R78912 VDD.n1366 VDD.n1211 4.5005
R78913 VDD.n1324 VDD.n1211 4.5005
R78914 VDD.n1368 VDD.n1211 4.5005
R78915 VDD.n1323 VDD.n1211 4.5005
R78916 VDD.n1369 VDD.n1211 4.5005
R78917 VDD.n1322 VDD.n1211 4.5005
R78918 VDD.n1371 VDD.n1211 4.5005
R78919 VDD.n1321 VDD.n1211 4.5005
R78920 VDD.n1372 VDD.n1211 4.5005
R78921 VDD.n1320 VDD.n1211 4.5005
R78922 VDD.n1374 VDD.n1211 4.5005
R78923 VDD.n1319 VDD.n1211 4.5005
R78924 VDD.n1375 VDD.n1211 4.5005
R78925 VDD.n1318 VDD.n1211 4.5005
R78926 VDD.n1376 VDD.n1211 4.5005
R78927 VDD.n1316 VDD.n1211 4.5005
R78928 VDD.n1377 VDD.n1211 4.5005
R78929 VDD.n1315 VDD.n1211 4.5005
R78930 VDD.n1378 VDD.n1211 4.5005
R78931 VDD.n1313 VDD.n1211 4.5005
R78932 VDD.n1379 VDD.n1211 4.5005
R78933 VDD.n1312 VDD.n1211 4.5005
R78934 VDD.n1380 VDD.n1211 4.5005
R78935 VDD.n1310 VDD.n1211 4.5005
R78936 VDD.n1381 VDD.n1211 4.5005
R78937 VDD.n1309 VDD.n1211 4.5005
R78938 VDD.n1382 VDD.n1211 4.5005
R78939 VDD.n1307 VDD.n1211 4.5005
R78940 VDD.n1383 VDD.n1211 4.5005
R78941 VDD.n1306 VDD.n1211 4.5005
R78942 VDD.n1384 VDD.n1211 4.5005
R78943 VDD.n1304 VDD.n1211 4.5005
R78944 VDD.n1385 VDD.n1211 4.5005
R78945 VDD.n1303 VDD.n1211 4.5005
R78946 VDD.n1386 VDD.n1211 4.5005
R78947 VDD.n1301 VDD.n1211 4.5005
R78948 VDD.n1387 VDD.n1211 4.5005
R78949 VDD.n1300 VDD.n1211 4.5005
R78950 VDD.n1388 VDD.n1211 4.5005
R78951 VDD.n1298 VDD.n1211 4.5005
R78952 VDD.n1389 VDD.n1211 4.5005
R78953 VDD.n1297 VDD.n1211 4.5005
R78954 VDD.n1390 VDD.n1211 4.5005
R78955 VDD.n1295 VDD.n1211 4.5005
R78956 VDD.n1391 VDD.n1211 4.5005
R78957 VDD.n1294 VDD.n1211 4.5005
R78958 VDD.n1392 VDD.n1211 4.5005
R78959 VDD.n1292 VDD.n1211 4.5005
R78960 VDD.n1393 VDD.n1211 4.5005
R78961 VDD.n1291 VDD.n1211 4.5005
R78962 VDD.n1394 VDD.n1211 4.5005
R78963 VDD.n1289 VDD.n1211 4.5005
R78964 VDD.n1395 VDD.n1211 4.5005
R78965 VDD.n1288 VDD.n1211 4.5005
R78966 VDD.n1396 VDD.n1211 4.5005
R78967 VDD.n1286 VDD.n1211 4.5005
R78968 VDD.n1397 VDD.n1211 4.5005
R78969 VDD.n1285 VDD.n1211 4.5005
R78970 VDD.n1398 VDD.n1211 4.5005
R78971 VDD.n1283 VDD.n1211 4.5005
R78972 VDD.n1399 VDD.n1211 4.5005
R78973 VDD.n1282 VDD.n1211 4.5005
R78974 VDD.n1400 VDD.n1211 4.5005
R78975 VDD.n1280 VDD.n1211 4.5005
R78976 VDD.n1401 VDD.n1211 4.5005
R78977 VDD.n1279 VDD.n1211 4.5005
R78978 VDD.n1402 VDD.n1211 4.5005
R78979 VDD.n1277 VDD.n1211 4.5005
R78980 VDD.n1403 VDD.n1211 4.5005
R78981 VDD.n1276 VDD.n1211 4.5005
R78982 VDD.n1404 VDD.n1211 4.5005
R78983 VDD.n1274 VDD.n1211 4.5005
R78984 VDD.n1405 VDD.n1211 4.5005
R78985 VDD.n1273 VDD.n1211 4.5005
R78986 VDD.n1406 VDD.n1211 4.5005
R78987 VDD.n1271 VDD.n1211 4.5005
R78988 VDD.n1407 VDD.n1211 4.5005
R78989 VDD.n1270 VDD.n1211 4.5005
R78990 VDD.n1408 VDD.n1211 4.5005
R78991 VDD.n1268 VDD.n1211 4.5005
R78992 VDD.n1409 VDD.n1211 4.5005
R78993 VDD.n1267 VDD.n1211 4.5005
R78994 VDD.n1410 VDD.n1211 4.5005
R78995 VDD.n1265 VDD.n1211 4.5005
R78996 VDD.n1411 VDD.n1211 4.5005
R78997 VDD.n1264 VDD.n1211 4.5005
R78998 VDD.n1412 VDD.n1211 4.5005
R78999 VDD.n1262 VDD.n1211 4.5005
R79000 VDD.n1413 VDD.n1211 4.5005
R79001 VDD.n1261 VDD.n1211 4.5005
R79002 VDD.n1414 VDD.n1211 4.5005
R79003 VDD.n1415 VDD.n1211 4.5005
R79004 VDD.n1674 VDD.n1211 4.5005
R79005 VDD.n1676 VDD.n1178 4.5005
R79006 VDD.n1341 VDD.n1178 4.5005
R79007 VDD.n1342 VDD.n1178 4.5005
R79008 VDD.n1340 VDD.n1178 4.5005
R79009 VDD.n1344 VDD.n1178 4.5005
R79010 VDD.n1339 VDD.n1178 4.5005
R79011 VDD.n1345 VDD.n1178 4.5005
R79012 VDD.n1338 VDD.n1178 4.5005
R79013 VDD.n1347 VDD.n1178 4.5005
R79014 VDD.n1337 VDD.n1178 4.5005
R79015 VDD.n1348 VDD.n1178 4.5005
R79016 VDD.n1336 VDD.n1178 4.5005
R79017 VDD.n1350 VDD.n1178 4.5005
R79018 VDD.n1335 VDD.n1178 4.5005
R79019 VDD.n1351 VDD.n1178 4.5005
R79020 VDD.n1334 VDD.n1178 4.5005
R79021 VDD.n1353 VDD.n1178 4.5005
R79022 VDD.n1333 VDD.n1178 4.5005
R79023 VDD.n1354 VDD.n1178 4.5005
R79024 VDD.n1332 VDD.n1178 4.5005
R79025 VDD.n1356 VDD.n1178 4.5005
R79026 VDD.n1331 VDD.n1178 4.5005
R79027 VDD.n1357 VDD.n1178 4.5005
R79028 VDD.n1330 VDD.n1178 4.5005
R79029 VDD.n1359 VDD.n1178 4.5005
R79030 VDD.n1329 VDD.n1178 4.5005
R79031 VDD.n1360 VDD.n1178 4.5005
R79032 VDD.n1328 VDD.n1178 4.5005
R79033 VDD.n1362 VDD.n1178 4.5005
R79034 VDD.n1327 VDD.n1178 4.5005
R79035 VDD.n1363 VDD.n1178 4.5005
R79036 VDD.n1326 VDD.n1178 4.5005
R79037 VDD.n1365 VDD.n1178 4.5005
R79038 VDD.n1325 VDD.n1178 4.5005
R79039 VDD.n1366 VDD.n1178 4.5005
R79040 VDD.n1324 VDD.n1178 4.5005
R79041 VDD.n1368 VDD.n1178 4.5005
R79042 VDD.n1323 VDD.n1178 4.5005
R79043 VDD.n1369 VDD.n1178 4.5005
R79044 VDD.n1322 VDD.n1178 4.5005
R79045 VDD.n1371 VDD.n1178 4.5005
R79046 VDD.n1321 VDD.n1178 4.5005
R79047 VDD.n1372 VDD.n1178 4.5005
R79048 VDD.n1320 VDD.n1178 4.5005
R79049 VDD.n1374 VDD.n1178 4.5005
R79050 VDD.n1319 VDD.n1178 4.5005
R79051 VDD.n1375 VDD.n1178 4.5005
R79052 VDD.n1318 VDD.n1178 4.5005
R79053 VDD.n1376 VDD.n1178 4.5005
R79054 VDD.n1316 VDD.n1178 4.5005
R79055 VDD.n1377 VDD.n1178 4.5005
R79056 VDD.n1315 VDD.n1178 4.5005
R79057 VDD.n1378 VDD.n1178 4.5005
R79058 VDD.n1313 VDD.n1178 4.5005
R79059 VDD.n1379 VDD.n1178 4.5005
R79060 VDD.n1312 VDD.n1178 4.5005
R79061 VDD.n1380 VDD.n1178 4.5005
R79062 VDD.n1310 VDD.n1178 4.5005
R79063 VDD.n1381 VDD.n1178 4.5005
R79064 VDD.n1309 VDD.n1178 4.5005
R79065 VDD.n1382 VDD.n1178 4.5005
R79066 VDD.n1307 VDD.n1178 4.5005
R79067 VDD.n1383 VDD.n1178 4.5005
R79068 VDD.n1306 VDD.n1178 4.5005
R79069 VDD.n1384 VDD.n1178 4.5005
R79070 VDD.n1304 VDD.n1178 4.5005
R79071 VDD.n1385 VDD.n1178 4.5005
R79072 VDD.n1303 VDD.n1178 4.5005
R79073 VDD.n1386 VDD.n1178 4.5005
R79074 VDD.n1301 VDD.n1178 4.5005
R79075 VDD.n1387 VDD.n1178 4.5005
R79076 VDD.n1300 VDD.n1178 4.5005
R79077 VDD.n1388 VDD.n1178 4.5005
R79078 VDD.n1298 VDD.n1178 4.5005
R79079 VDD.n1389 VDD.n1178 4.5005
R79080 VDD.n1297 VDD.n1178 4.5005
R79081 VDD.n1390 VDD.n1178 4.5005
R79082 VDD.n1295 VDD.n1178 4.5005
R79083 VDD.n1391 VDD.n1178 4.5005
R79084 VDD.n1294 VDD.n1178 4.5005
R79085 VDD.n1392 VDD.n1178 4.5005
R79086 VDD.n1292 VDD.n1178 4.5005
R79087 VDD.n1393 VDD.n1178 4.5005
R79088 VDD.n1291 VDD.n1178 4.5005
R79089 VDD.n1394 VDD.n1178 4.5005
R79090 VDD.n1289 VDD.n1178 4.5005
R79091 VDD.n1395 VDD.n1178 4.5005
R79092 VDD.n1288 VDD.n1178 4.5005
R79093 VDD.n1396 VDD.n1178 4.5005
R79094 VDD.n1286 VDD.n1178 4.5005
R79095 VDD.n1397 VDD.n1178 4.5005
R79096 VDD.n1285 VDD.n1178 4.5005
R79097 VDD.n1398 VDD.n1178 4.5005
R79098 VDD.n1283 VDD.n1178 4.5005
R79099 VDD.n1399 VDD.n1178 4.5005
R79100 VDD.n1282 VDD.n1178 4.5005
R79101 VDD.n1400 VDD.n1178 4.5005
R79102 VDD.n1280 VDD.n1178 4.5005
R79103 VDD.n1401 VDD.n1178 4.5005
R79104 VDD.n1279 VDD.n1178 4.5005
R79105 VDD.n1402 VDD.n1178 4.5005
R79106 VDD.n1277 VDD.n1178 4.5005
R79107 VDD.n1403 VDD.n1178 4.5005
R79108 VDD.n1276 VDD.n1178 4.5005
R79109 VDD.n1404 VDD.n1178 4.5005
R79110 VDD.n1274 VDD.n1178 4.5005
R79111 VDD.n1405 VDD.n1178 4.5005
R79112 VDD.n1273 VDD.n1178 4.5005
R79113 VDD.n1406 VDD.n1178 4.5005
R79114 VDD.n1271 VDD.n1178 4.5005
R79115 VDD.n1407 VDD.n1178 4.5005
R79116 VDD.n1270 VDD.n1178 4.5005
R79117 VDD.n1408 VDD.n1178 4.5005
R79118 VDD.n1268 VDD.n1178 4.5005
R79119 VDD.n1409 VDD.n1178 4.5005
R79120 VDD.n1267 VDD.n1178 4.5005
R79121 VDD.n1410 VDD.n1178 4.5005
R79122 VDD.n1265 VDD.n1178 4.5005
R79123 VDD.n1411 VDD.n1178 4.5005
R79124 VDD.n1264 VDD.n1178 4.5005
R79125 VDD.n1412 VDD.n1178 4.5005
R79126 VDD.n1262 VDD.n1178 4.5005
R79127 VDD.n1413 VDD.n1178 4.5005
R79128 VDD.n1261 VDD.n1178 4.5005
R79129 VDD.n1414 VDD.n1178 4.5005
R79130 VDD.n1415 VDD.n1178 4.5005
R79131 VDD.n1674 VDD.n1178 4.5005
R79132 VDD.n1676 VDD.n1212 4.5005
R79133 VDD.n1341 VDD.n1212 4.5005
R79134 VDD.n1342 VDD.n1212 4.5005
R79135 VDD.n1340 VDD.n1212 4.5005
R79136 VDD.n1344 VDD.n1212 4.5005
R79137 VDD.n1339 VDD.n1212 4.5005
R79138 VDD.n1345 VDD.n1212 4.5005
R79139 VDD.n1338 VDD.n1212 4.5005
R79140 VDD.n1347 VDD.n1212 4.5005
R79141 VDD.n1337 VDD.n1212 4.5005
R79142 VDD.n1348 VDD.n1212 4.5005
R79143 VDD.n1336 VDD.n1212 4.5005
R79144 VDD.n1350 VDD.n1212 4.5005
R79145 VDD.n1335 VDD.n1212 4.5005
R79146 VDD.n1351 VDD.n1212 4.5005
R79147 VDD.n1334 VDD.n1212 4.5005
R79148 VDD.n1353 VDD.n1212 4.5005
R79149 VDD.n1333 VDD.n1212 4.5005
R79150 VDD.n1354 VDD.n1212 4.5005
R79151 VDD.n1332 VDD.n1212 4.5005
R79152 VDD.n1356 VDD.n1212 4.5005
R79153 VDD.n1331 VDD.n1212 4.5005
R79154 VDD.n1357 VDD.n1212 4.5005
R79155 VDD.n1330 VDD.n1212 4.5005
R79156 VDD.n1359 VDD.n1212 4.5005
R79157 VDD.n1329 VDD.n1212 4.5005
R79158 VDD.n1360 VDD.n1212 4.5005
R79159 VDD.n1328 VDD.n1212 4.5005
R79160 VDD.n1362 VDD.n1212 4.5005
R79161 VDD.n1327 VDD.n1212 4.5005
R79162 VDD.n1363 VDD.n1212 4.5005
R79163 VDD.n1326 VDD.n1212 4.5005
R79164 VDD.n1365 VDD.n1212 4.5005
R79165 VDD.n1325 VDD.n1212 4.5005
R79166 VDD.n1366 VDD.n1212 4.5005
R79167 VDD.n1324 VDD.n1212 4.5005
R79168 VDD.n1368 VDD.n1212 4.5005
R79169 VDD.n1323 VDD.n1212 4.5005
R79170 VDD.n1369 VDD.n1212 4.5005
R79171 VDD.n1322 VDD.n1212 4.5005
R79172 VDD.n1371 VDD.n1212 4.5005
R79173 VDD.n1321 VDD.n1212 4.5005
R79174 VDD.n1372 VDD.n1212 4.5005
R79175 VDD.n1320 VDD.n1212 4.5005
R79176 VDD.n1374 VDD.n1212 4.5005
R79177 VDD.n1319 VDD.n1212 4.5005
R79178 VDD.n1375 VDD.n1212 4.5005
R79179 VDD.n1318 VDD.n1212 4.5005
R79180 VDD.n1376 VDD.n1212 4.5005
R79181 VDD.n1316 VDD.n1212 4.5005
R79182 VDD.n1377 VDD.n1212 4.5005
R79183 VDD.n1315 VDD.n1212 4.5005
R79184 VDD.n1378 VDD.n1212 4.5005
R79185 VDD.n1313 VDD.n1212 4.5005
R79186 VDD.n1379 VDD.n1212 4.5005
R79187 VDD.n1312 VDD.n1212 4.5005
R79188 VDD.n1380 VDD.n1212 4.5005
R79189 VDD.n1310 VDD.n1212 4.5005
R79190 VDD.n1381 VDD.n1212 4.5005
R79191 VDD.n1309 VDD.n1212 4.5005
R79192 VDD.n1382 VDD.n1212 4.5005
R79193 VDD.n1307 VDD.n1212 4.5005
R79194 VDD.n1383 VDD.n1212 4.5005
R79195 VDD.n1306 VDD.n1212 4.5005
R79196 VDD.n1384 VDD.n1212 4.5005
R79197 VDD.n1304 VDD.n1212 4.5005
R79198 VDD.n1385 VDD.n1212 4.5005
R79199 VDD.n1303 VDD.n1212 4.5005
R79200 VDD.n1386 VDD.n1212 4.5005
R79201 VDD.n1301 VDD.n1212 4.5005
R79202 VDD.n1387 VDD.n1212 4.5005
R79203 VDD.n1300 VDD.n1212 4.5005
R79204 VDD.n1388 VDD.n1212 4.5005
R79205 VDD.n1298 VDD.n1212 4.5005
R79206 VDD.n1389 VDD.n1212 4.5005
R79207 VDD.n1297 VDD.n1212 4.5005
R79208 VDD.n1390 VDD.n1212 4.5005
R79209 VDD.n1295 VDD.n1212 4.5005
R79210 VDD.n1391 VDD.n1212 4.5005
R79211 VDD.n1294 VDD.n1212 4.5005
R79212 VDD.n1392 VDD.n1212 4.5005
R79213 VDD.n1292 VDD.n1212 4.5005
R79214 VDD.n1393 VDD.n1212 4.5005
R79215 VDD.n1291 VDD.n1212 4.5005
R79216 VDD.n1394 VDD.n1212 4.5005
R79217 VDD.n1289 VDD.n1212 4.5005
R79218 VDD.n1395 VDD.n1212 4.5005
R79219 VDD.n1288 VDD.n1212 4.5005
R79220 VDD.n1396 VDD.n1212 4.5005
R79221 VDD.n1286 VDD.n1212 4.5005
R79222 VDD.n1397 VDD.n1212 4.5005
R79223 VDD.n1285 VDD.n1212 4.5005
R79224 VDD.n1398 VDD.n1212 4.5005
R79225 VDD.n1283 VDD.n1212 4.5005
R79226 VDD.n1399 VDD.n1212 4.5005
R79227 VDD.n1282 VDD.n1212 4.5005
R79228 VDD.n1400 VDD.n1212 4.5005
R79229 VDD.n1280 VDD.n1212 4.5005
R79230 VDD.n1401 VDD.n1212 4.5005
R79231 VDD.n1279 VDD.n1212 4.5005
R79232 VDD.n1402 VDD.n1212 4.5005
R79233 VDD.n1277 VDD.n1212 4.5005
R79234 VDD.n1403 VDD.n1212 4.5005
R79235 VDD.n1276 VDD.n1212 4.5005
R79236 VDD.n1404 VDD.n1212 4.5005
R79237 VDD.n1274 VDD.n1212 4.5005
R79238 VDD.n1405 VDD.n1212 4.5005
R79239 VDD.n1273 VDD.n1212 4.5005
R79240 VDD.n1406 VDD.n1212 4.5005
R79241 VDD.n1271 VDD.n1212 4.5005
R79242 VDD.n1407 VDD.n1212 4.5005
R79243 VDD.n1270 VDD.n1212 4.5005
R79244 VDD.n1408 VDD.n1212 4.5005
R79245 VDD.n1268 VDD.n1212 4.5005
R79246 VDD.n1409 VDD.n1212 4.5005
R79247 VDD.n1267 VDD.n1212 4.5005
R79248 VDD.n1410 VDD.n1212 4.5005
R79249 VDD.n1265 VDD.n1212 4.5005
R79250 VDD.n1411 VDD.n1212 4.5005
R79251 VDD.n1264 VDD.n1212 4.5005
R79252 VDD.n1412 VDD.n1212 4.5005
R79253 VDD.n1262 VDD.n1212 4.5005
R79254 VDD.n1413 VDD.n1212 4.5005
R79255 VDD.n1261 VDD.n1212 4.5005
R79256 VDD.n1414 VDD.n1212 4.5005
R79257 VDD.n1415 VDD.n1212 4.5005
R79258 VDD.n1674 VDD.n1212 4.5005
R79259 VDD.n1676 VDD.n1177 4.5005
R79260 VDD.n1341 VDD.n1177 4.5005
R79261 VDD.n1342 VDD.n1177 4.5005
R79262 VDD.n1340 VDD.n1177 4.5005
R79263 VDD.n1344 VDD.n1177 4.5005
R79264 VDD.n1339 VDD.n1177 4.5005
R79265 VDD.n1345 VDD.n1177 4.5005
R79266 VDD.n1338 VDD.n1177 4.5005
R79267 VDD.n1347 VDD.n1177 4.5005
R79268 VDD.n1337 VDD.n1177 4.5005
R79269 VDD.n1348 VDD.n1177 4.5005
R79270 VDD.n1336 VDD.n1177 4.5005
R79271 VDD.n1350 VDD.n1177 4.5005
R79272 VDD.n1335 VDD.n1177 4.5005
R79273 VDD.n1351 VDD.n1177 4.5005
R79274 VDD.n1334 VDD.n1177 4.5005
R79275 VDD.n1353 VDD.n1177 4.5005
R79276 VDD.n1333 VDD.n1177 4.5005
R79277 VDD.n1354 VDD.n1177 4.5005
R79278 VDD.n1332 VDD.n1177 4.5005
R79279 VDD.n1356 VDD.n1177 4.5005
R79280 VDD.n1331 VDD.n1177 4.5005
R79281 VDD.n1357 VDD.n1177 4.5005
R79282 VDD.n1330 VDD.n1177 4.5005
R79283 VDD.n1359 VDD.n1177 4.5005
R79284 VDD.n1329 VDD.n1177 4.5005
R79285 VDD.n1360 VDD.n1177 4.5005
R79286 VDD.n1328 VDD.n1177 4.5005
R79287 VDD.n1362 VDD.n1177 4.5005
R79288 VDD.n1327 VDD.n1177 4.5005
R79289 VDD.n1363 VDD.n1177 4.5005
R79290 VDD.n1326 VDD.n1177 4.5005
R79291 VDD.n1365 VDD.n1177 4.5005
R79292 VDD.n1325 VDD.n1177 4.5005
R79293 VDD.n1366 VDD.n1177 4.5005
R79294 VDD.n1324 VDD.n1177 4.5005
R79295 VDD.n1368 VDD.n1177 4.5005
R79296 VDD.n1323 VDD.n1177 4.5005
R79297 VDD.n1369 VDD.n1177 4.5005
R79298 VDD.n1322 VDD.n1177 4.5005
R79299 VDD.n1371 VDD.n1177 4.5005
R79300 VDD.n1321 VDD.n1177 4.5005
R79301 VDD.n1372 VDD.n1177 4.5005
R79302 VDD.n1320 VDD.n1177 4.5005
R79303 VDD.n1374 VDD.n1177 4.5005
R79304 VDD.n1319 VDD.n1177 4.5005
R79305 VDD.n1375 VDD.n1177 4.5005
R79306 VDD.n1318 VDD.n1177 4.5005
R79307 VDD.n1376 VDD.n1177 4.5005
R79308 VDD.n1316 VDD.n1177 4.5005
R79309 VDD.n1377 VDD.n1177 4.5005
R79310 VDD.n1315 VDD.n1177 4.5005
R79311 VDD.n1378 VDD.n1177 4.5005
R79312 VDD.n1313 VDD.n1177 4.5005
R79313 VDD.n1379 VDD.n1177 4.5005
R79314 VDD.n1312 VDD.n1177 4.5005
R79315 VDD.n1380 VDD.n1177 4.5005
R79316 VDD.n1310 VDD.n1177 4.5005
R79317 VDD.n1381 VDD.n1177 4.5005
R79318 VDD.n1309 VDD.n1177 4.5005
R79319 VDD.n1382 VDD.n1177 4.5005
R79320 VDD.n1307 VDD.n1177 4.5005
R79321 VDD.n1383 VDD.n1177 4.5005
R79322 VDD.n1306 VDD.n1177 4.5005
R79323 VDD.n1384 VDD.n1177 4.5005
R79324 VDD.n1304 VDD.n1177 4.5005
R79325 VDD.n1385 VDD.n1177 4.5005
R79326 VDD.n1303 VDD.n1177 4.5005
R79327 VDD.n1386 VDD.n1177 4.5005
R79328 VDD.n1301 VDD.n1177 4.5005
R79329 VDD.n1387 VDD.n1177 4.5005
R79330 VDD.n1300 VDD.n1177 4.5005
R79331 VDD.n1388 VDD.n1177 4.5005
R79332 VDD.n1298 VDD.n1177 4.5005
R79333 VDD.n1389 VDD.n1177 4.5005
R79334 VDD.n1297 VDD.n1177 4.5005
R79335 VDD.n1390 VDD.n1177 4.5005
R79336 VDD.n1295 VDD.n1177 4.5005
R79337 VDD.n1391 VDD.n1177 4.5005
R79338 VDD.n1294 VDD.n1177 4.5005
R79339 VDD.n1392 VDD.n1177 4.5005
R79340 VDD.n1292 VDD.n1177 4.5005
R79341 VDD.n1393 VDD.n1177 4.5005
R79342 VDD.n1291 VDD.n1177 4.5005
R79343 VDD.n1394 VDD.n1177 4.5005
R79344 VDD.n1289 VDD.n1177 4.5005
R79345 VDD.n1395 VDD.n1177 4.5005
R79346 VDD.n1288 VDD.n1177 4.5005
R79347 VDD.n1396 VDD.n1177 4.5005
R79348 VDD.n1286 VDD.n1177 4.5005
R79349 VDD.n1397 VDD.n1177 4.5005
R79350 VDD.n1285 VDD.n1177 4.5005
R79351 VDD.n1398 VDD.n1177 4.5005
R79352 VDD.n1283 VDD.n1177 4.5005
R79353 VDD.n1399 VDD.n1177 4.5005
R79354 VDD.n1282 VDD.n1177 4.5005
R79355 VDD.n1400 VDD.n1177 4.5005
R79356 VDD.n1280 VDD.n1177 4.5005
R79357 VDD.n1401 VDD.n1177 4.5005
R79358 VDD.n1279 VDD.n1177 4.5005
R79359 VDD.n1402 VDD.n1177 4.5005
R79360 VDD.n1277 VDD.n1177 4.5005
R79361 VDD.n1403 VDD.n1177 4.5005
R79362 VDD.n1276 VDD.n1177 4.5005
R79363 VDD.n1404 VDD.n1177 4.5005
R79364 VDD.n1274 VDD.n1177 4.5005
R79365 VDD.n1405 VDD.n1177 4.5005
R79366 VDD.n1273 VDD.n1177 4.5005
R79367 VDD.n1406 VDD.n1177 4.5005
R79368 VDD.n1271 VDD.n1177 4.5005
R79369 VDD.n1407 VDD.n1177 4.5005
R79370 VDD.n1270 VDD.n1177 4.5005
R79371 VDD.n1408 VDD.n1177 4.5005
R79372 VDD.n1268 VDD.n1177 4.5005
R79373 VDD.n1409 VDD.n1177 4.5005
R79374 VDD.n1267 VDD.n1177 4.5005
R79375 VDD.n1410 VDD.n1177 4.5005
R79376 VDD.n1265 VDD.n1177 4.5005
R79377 VDD.n1411 VDD.n1177 4.5005
R79378 VDD.n1264 VDD.n1177 4.5005
R79379 VDD.n1412 VDD.n1177 4.5005
R79380 VDD.n1262 VDD.n1177 4.5005
R79381 VDD.n1413 VDD.n1177 4.5005
R79382 VDD.n1261 VDD.n1177 4.5005
R79383 VDD.n1414 VDD.n1177 4.5005
R79384 VDD.n1415 VDD.n1177 4.5005
R79385 VDD.n1674 VDD.n1177 4.5005
R79386 VDD.n1676 VDD.n1213 4.5005
R79387 VDD.n1341 VDD.n1213 4.5005
R79388 VDD.n1342 VDD.n1213 4.5005
R79389 VDD.n1340 VDD.n1213 4.5005
R79390 VDD.n1344 VDD.n1213 4.5005
R79391 VDD.n1339 VDD.n1213 4.5005
R79392 VDD.n1345 VDD.n1213 4.5005
R79393 VDD.n1338 VDD.n1213 4.5005
R79394 VDD.n1347 VDD.n1213 4.5005
R79395 VDD.n1337 VDD.n1213 4.5005
R79396 VDD.n1348 VDD.n1213 4.5005
R79397 VDD.n1336 VDD.n1213 4.5005
R79398 VDD.n1350 VDD.n1213 4.5005
R79399 VDD.n1335 VDD.n1213 4.5005
R79400 VDD.n1351 VDD.n1213 4.5005
R79401 VDD.n1334 VDD.n1213 4.5005
R79402 VDD.n1353 VDD.n1213 4.5005
R79403 VDD.n1333 VDD.n1213 4.5005
R79404 VDD.n1354 VDD.n1213 4.5005
R79405 VDD.n1332 VDD.n1213 4.5005
R79406 VDD.n1356 VDD.n1213 4.5005
R79407 VDD.n1331 VDD.n1213 4.5005
R79408 VDD.n1357 VDD.n1213 4.5005
R79409 VDD.n1330 VDD.n1213 4.5005
R79410 VDD.n1359 VDD.n1213 4.5005
R79411 VDD.n1329 VDD.n1213 4.5005
R79412 VDD.n1360 VDD.n1213 4.5005
R79413 VDD.n1328 VDD.n1213 4.5005
R79414 VDD.n1362 VDD.n1213 4.5005
R79415 VDD.n1327 VDD.n1213 4.5005
R79416 VDD.n1363 VDD.n1213 4.5005
R79417 VDD.n1326 VDD.n1213 4.5005
R79418 VDD.n1365 VDD.n1213 4.5005
R79419 VDD.n1325 VDD.n1213 4.5005
R79420 VDD.n1366 VDD.n1213 4.5005
R79421 VDD.n1324 VDD.n1213 4.5005
R79422 VDD.n1368 VDD.n1213 4.5005
R79423 VDD.n1323 VDD.n1213 4.5005
R79424 VDD.n1369 VDD.n1213 4.5005
R79425 VDD.n1322 VDD.n1213 4.5005
R79426 VDD.n1371 VDD.n1213 4.5005
R79427 VDD.n1321 VDD.n1213 4.5005
R79428 VDD.n1372 VDD.n1213 4.5005
R79429 VDD.n1320 VDD.n1213 4.5005
R79430 VDD.n1374 VDD.n1213 4.5005
R79431 VDD.n1319 VDD.n1213 4.5005
R79432 VDD.n1375 VDD.n1213 4.5005
R79433 VDD.n1318 VDD.n1213 4.5005
R79434 VDD.n1376 VDD.n1213 4.5005
R79435 VDD.n1316 VDD.n1213 4.5005
R79436 VDD.n1377 VDD.n1213 4.5005
R79437 VDD.n1315 VDD.n1213 4.5005
R79438 VDD.n1378 VDD.n1213 4.5005
R79439 VDD.n1313 VDD.n1213 4.5005
R79440 VDD.n1379 VDD.n1213 4.5005
R79441 VDD.n1312 VDD.n1213 4.5005
R79442 VDD.n1380 VDD.n1213 4.5005
R79443 VDD.n1310 VDD.n1213 4.5005
R79444 VDD.n1381 VDD.n1213 4.5005
R79445 VDD.n1309 VDD.n1213 4.5005
R79446 VDD.n1382 VDD.n1213 4.5005
R79447 VDD.n1307 VDD.n1213 4.5005
R79448 VDD.n1383 VDD.n1213 4.5005
R79449 VDD.n1306 VDD.n1213 4.5005
R79450 VDD.n1384 VDD.n1213 4.5005
R79451 VDD.n1304 VDD.n1213 4.5005
R79452 VDD.n1385 VDD.n1213 4.5005
R79453 VDD.n1303 VDD.n1213 4.5005
R79454 VDD.n1386 VDD.n1213 4.5005
R79455 VDD.n1301 VDD.n1213 4.5005
R79456 VDD.n1387 VDD.n1213 4.5005
R79457 VDD.n1300 VDD.n1213 4.5005
R79458 VDD.n1388 VDD.n1213 4.5005
R79459 VDD.n1298 VDD.n1213 4.5005
R79460 VDD.n1389 VDD.n1213 4.5005
R79461 VDD.n1297 VDD.n1213 4.5005
R79462 VDD.n1390 VDD.n1213 4.5005
R79463 VDD.n1295 VDD.n1213 4.5005
R79464 VDD.n1391 VDD.n1213 4.5005
R79465 VDD.n1294 VDD.n1213 4.5005
R79466 VDD.n1392 VDD.n1213 4.5005
R79467 VDD.n1292 VDD.n1213 4.5005
R79468 VDD.n1393 VDD.n1213 4.5005
R79469 VDD.n1291 VDD.n1213 4.5005
R79470 VDD.n1394 VDD.n1213 4.5005
R79471 VDD.n1289 VDD.n1213 4.5005
R79472 VDD.n1395 VDD.n1213 4.5005
R79473 VDD.n1288 VDD.n1213 4.5005
R79474 VDD.n1396 VDD.n1213 4.5005
R79475 VDD.n1286 VDD.n1213 4.5005
R79476 VDD.n1397 VDD.n1213 4.5005
R79477 VDD.n1285 VDD.n1213 4.5005
R79478 VDD.n1398 VDD.n1213 4.5005
R79479 VDD.n1283 VDD.n1213 4.5005
R79480 VDD.n1399 VDD.n1213 4.5005
R79481 VDD.n1282 VDD.n1213 4.5005
R79482 VDD.n1400 VDD.n1213 4.5005
R79483 VDD.n1280 VDD.n1213 4.5005
R79484 VDD.n1401 VDD.n1213 4.5005
R79485 VDD.n1279 VDD.n1213 4.5005
R79486 VDD.n1402 VDD.n1213 4.5005
R79487 VDD.n1277 VDD.n1213 4.5005
R79488 VDD.n1403 VDD.n1213 4.5005
R79489 VDD.n1276 VDD.n1213 4.5005
R79490 VDD.n1404 VDD.n1213 4.5005
R79491 VDD.n1274 VDD.n1213 4.5005
R79492 VDD.n1405 VDD.n1213 4.5005
R79493 VDD.n1273 VDD.n1213 4.5005
R79494 VDD.n1406 VDD.n1213 4.5005
R79495 VDD.n1271 VDD.n1213 4.5005
R79496 VDD.n1407 VDD.n1213 4.5005
R79497 VDD.n1270 VDD.n1213 4.5005
R79498 VDD.n1408 VDD.n1213 4.5005
R79499 VDD.n1268 VDD.n1213 4.5005
R79500 VDD.n1409 VDD.n1213 4.5005
R79501 VDD.n1267 VDD.n1213 4.5005
R79502 VDD.n1410 VDD.n1213 4.5005
R79503 VDD.n1265 VDD.n1213 4.5005
R79504 VDD.n1411 VDD.n1213 4.5005
R79505 VDD.n1264 VDD.n1213 4.5005
R79506 VDD.n1412 VDD.n1213 4.5005
R79507 VDD.n1262 VDD.n1213 4.5005
R79508 VDD.n1413 VDD.n1213 4.5005
R79509 VDD.n1261 VDD.n1213 4.5005
R79510 VDD.n1414 VDD.n1213 4.5005
R79511 VDD.n1415 VDD.n1213 4.5005
R79512 VDD.n1674 VDD.n1213 4.5005
R79513 VDD.n1676 VDD.n1176 4.5005
R79514 VDD.n1341 VDD.n1176 4.5005
R79515 VDD.n1342 VDD.n1176 4.5005
R79516 VDD.n1340 VDD.n1176 4.5005
R79517 VDD.n1344 VDD.n1176 4.5005
R79518 VDD.n1339 VDD.n1176 4.5005
R79519 VDD.n1345 VDD.n1176 4.5005
R79520 VDD.n1338 VDD.n1176 4.5005
R79521 VDD.n1347 VDD.n1176 4.5005
R79522 VDD.n1337 VDD.n1176 4.5005
R79523 VDD.n1348 VDD.n1176 4.5005
R79524 VDD.n1336 VDD.n1176 4.5005
R79525 VDD.n1350 VDD.n1176 4.5005
R79526 VDD.n1335 VDD.n1176 4.5005
R79527 VDD.n1351 VDD.n1176 4.5005
R79528 VDD.n1334 VDD.n1176 4.5005
R79529 VDD.n1353 VDD.n1176 4.5005
R79530 VDD.n1333 VDD.n1176 4.5005
R79531 VDD.n1354 VDD.n1176 4.5005
R79532 VDD.n1332 VDD.n1176 4.5005
R79533 VDD.n1356 VDD.n1176 4.5005
R79534 VDD.n1331 VDD.n1176 4.5005
R79535 VDD.n1357 VDD.n1176 4.5005
R79536 VDD.n1330 VDD.n1176 4.5005
R79537 VDD.n1359 VDD.n1176 4.5005
R79538 VDD.n1329 VDD.n1176 4.5005
R79539 VDD.n1360 VDD.n1176 4.5005
R79540 VDD.n1328 VDD.n1176 4.5005
R79541 VDD.n1362 VDD.n1176 4.5005
R79542 VDD.n1327 VDD.n1176 4.5005
R79543 VDD.n1363 VDD.n1176 4.5005
R79544 VDD.n1326 VDD.n1176 4.5005
R79545 VDD.n1365 VDD.n1176 4.5005
R79546 VDD.n1325 VDD.n1176 4.5005
R79547 VDD.n1366 VDD.n1176 4.5005
R79548 VDD.n1324 VDD.n1176 4.5005
R79549 VDD.n1368 VDD.n1176 4.5005
R79550 VDD.n1323 VDD.n1176 4.5005
R79551 VDD.n1369 VDD.n1176 4.5005
R79552 VDD.n1322 VDD.n1176 4.5005
R79553 VDD.n1371 VDD.n1176 4.5005
R79554 VDD.n1321 VDD.n1176 4.5005
R79555 VDD.n1372 VDD.n1176 4.5005
R79556 VDD.n1320 VDD.n1176 4.5005
R79557 VDD.n1374 VDD.n1176 4.5005
R79558 VDD.n1319 VDD.n1176 4.5005
R79559 VDD.n1375 VDD.n1176 4.5005
R79560 VDD.n1318 VDD.n1176 4.5005
R79561 VDD.n1376 VDD.n1176 4.5005
R79562 VDD.n1316 VDD.n1176 4.5005
R79563 VDD.n1377 VDD.n1176 4.5005
R79564 VDD.n1315 VDD.n1176 4.5005
R79565 VDD.n1378 VDD.n1176 4.5005
R79566 VDD.n1313 VDD.n1176 4.5005
R79567 VDD.n1379 VDD.n1176 4.5005
R79568 VDD.n1312 VDD.n1176 4.5005
R79569 VDD.n1380 VDD.n1176 4.5005
R79570 VDD.n1310 VDD.n1176 4.5005
R79571 VDD.n1381 VDD.n1176 4.5005
R79572 VDD.n1309 VDD.n1176 4.5005
R79573 VDD.n1382 VDD.n1176 4.5005
R79574 VDD.n1307 VDD.n1176 4.5005
R79575 VDD.n1383 VDD.n1176 4.5005
R79576 VDD.n1306 VDD.n1176 4.5005
R79577 VDD.n1384 VDD.n1176 4.5005
R79578 VDD.n1304 VDD.n1176 4.5005
R79579 VDD.n1385 VDD.n1176 4.5005
R79580 VDD.n1303 VDD.n1176 4.5005
R79581 VDD.n1386 VDD.n1176 4.5005
R79582 VDD.n1301 VDD.n1176 4.5005
R79583 VDD.n1387 VDD.n1176 4.5005
R79584 VDD.n1300 VDD.n1176 4.5005
R79585 VDD.n1388 VDD.n1176 4.5005
R79586 VDD.n1298 VDD.n1176 4.5005
R79587 VDD.n1389 VDD.n1176 4.5005
R79588 VDD.n1297 VDD.n1176 4.5005
R79589 VDD.n1390 VDD.n1176 4.5005
R79590 VDD.n1295 VDD.n1176 4.5005
R79591 VDD.n1391 VDD.n1176 4.5005
R79592 VDD.n1294 VDD.n1176 4.5005
R79593 VDD.n1392 VDD.n1176 4.5005
R79594 VDD.n1292 VDD.n1176 4.5005
R79595 VDD.n1393 VDD.n1176 4.5005
R79596 VDD.n1291 VDD.n1176 4.5005
R79597 VDD.n1394 VDD.n1176 4.5005
R79598 VDD.n1289 VDD.n1176 4.5005
R79599 VDD.n1395 VDD.n1176 4.5005
R79600 VDD.n1288 VDD.n1176 4.5005
R79601 VDD.n1396 VDD.n1176 4.5005
R79602 VDD.n1286 VDD.n1176 4.5005
R79603 VDD.n1397 VDD.n1176 4.5005
R79604 VDD.n1285 VDD.n1176 4.5005
R79605 VDD.n1398 VDD.n1176 4.5005
R79606 VDD.n1283 VDD.n1176 4.5005
R79607 VDD.n1399 VDD.n1176 4.5005
R79608 VDD.n1282 VDD.n1176 4.5005
R79609 VDD.n1400 VDD.n1176 4.5005
R79610 VDD.n1280 VDD.n1176 4.5005
R79611 VDD.n1401 VDD.n1176 4.5005
R79612 VDD.n1279 VDD.n1176 4.5005
R79613 VDD.n1402 VDD.n1176 4.5005
R79614 VDD.n1277 VDD.n1176 4.5005
R79615 VDD.n1403 VDD.n1176 4.5005
R79616 VDD.n1276 VDD.n1176 4.5005
R79617 VDD.n1404 VDD.n1176 4.5005
R79618 VDD.n1274 VDD.n1176 4.5005
R79619 VDD.n1405 VDD.n1176 4.5005
R79620 VDD.n1273 VDD.n1176 4.5005
R79621 VDD.n1406 VDD.n1176 4.5005
R79622 VDD.n1271 VDD.n1176 4.5005
R79623 VDD.n1407 VDD.n1176 4.5005
R79624 VDD.n1270 VDD.n1176 4.5005
R79625 VDD.n1408 VDD.n1176 4.5005
R79626 VDD.n1268 VDD.n1176 4.5005
R79627 VDD.n1409 VDD.n1176 4.5005
R79628 VDD.n1267 VDD.n1176 4.5005
R79629 VDD.n1410 VDD.n1176 4.5005
R79630 VDD.n1265 VDD.n1176 4.5005
R79631 VDD.n1411 VDD.n1176 4.5005
R79632 VDD.n1264 VDD.n1176 4.5005
R79633 VDD.n1412 VDD.n1176 4.5005
R79634 VDD.n1262 VDD.n1176 4.5005
R79635 VDD.n1413 VDD.n1176 4.5005
R79636 VDD.n1261 VDD.n1176 4.5005
R79637 VDD.n1414 VDD.n1176 4.5005
R79638 VDD.n1415 VDD.n1176 4.5005
R79639 VDD.n1674 VDD.n1176 4.5005
R79640 VDD.n1676 VDD.n1214 4.5005
R79641 VDD.n1341 VDD.n1214 4.5005
R79642 VDD.n1342 VDD.n1214 4.5005
R79643 VDD.n1340 VDD.n1214 4.5005
R79644 VDD.n1344 VDD.n1214 4.5005
R79645 VDD.n1339 VDD.n1214 4.5005
R79646 VDD.n1345 VDD.n1214 4.5005
R79647 VDD.n1338 VDD.n1214 4.5005
R79648 VDD.n1347 VDD.n1214 4.5005
R79649 VDD.n1337 VDD.n1214 4.5005
R79650 VDD.n1348 VDD.n1214 4.5005
R79651 VDD.n1336 VDD.n1214 4.5005
R79652 VDD.n1350 VDD.n1214 4.5005
R79653 VDD.n1335 VDD.n1214 4.5005
R79654 VDD.n1351 VDD.n1214 4.5005
R79655 VDD.n1334 VDD.n1214 4.5005
R79656 VDD.n1353 VDD.n1214 4.5005
R79657 VDD.n1333 VDD.n1214 4.5005
R79658 VDD.n1354 VDD.n1214 4.5005
R79659 VDD.n1332 VDD.n1214 4.5005
R79660 VDD.n1356 VDD.n1214 4.5005
R79661 VDD.n1331 VDD.n1214 4.5005
R79662 VDD.n1357 VDD.n1214 4.5005
R79663 VDD.n1330 VDD.n1214 4.5005
R79664 VDD.n1359 VDD.n1214 4.5005
R79665 VDD.n1329 VDD.n1214 4.5005
R79666 VDD.n1360 VDD.n1214 4.5005
R79667 VDD.n1328 VDD.n1214 4.5005
R79668 VDD.n1362 VDD.n1214 4.5005
R79669 VDD.n1327 VDD.n1214 4.5005
R79670 VDD.n1363 VDD.n1214 4.5005
R79671 VDD.n1326 VDD.n1214 4.5005
R79672 VDD.n1365 VDD.n1214 4.5005
R79673 VDD.n1325 VDD.n1214 4.5005
R79674 VDD.n1366 VDD.n1214 4.5005
R79675 VDD.n1324 VDD.n1214 4.5005
R79676 VDD.n1368 VDD.n1214 4.5005
R79677 VDD.n1323 VDD.n1214 4.5005
R79678 VDD.n1369 VDD.n1214 4.5005
R79679 VDD.n1322 VDD.n1214 4.5005
R79680 VDD.n1371 VDD.n1214 4.5005
R79681 VDD.n1321 VDD.n1214 4.5005
R79682 VDD.n1372 VDD.n1214 4.5005
R79683 VDD.n1320 VDD.n1214 4.5005
R79684 VDD.n1374 VDD.n1214 4.5005
R79685 VDD.n1319 VDD.n1214 4.5005
R79686 VDD.n1375 VDD.n1214 4.5005
R79687 VDD.n1318 VDD.n1214 4.5005
R79688 VDD.n1376 VDD.n1214 4.5005
R79689 VDD.n1316 VDD.n1214 4.5005
R79690 VDD.n1377 VDD.n1214 4.5005
R79691 VDD.n1315 VDD.n1214 4.5005
R79692 VDD.n1378 VDD.n1214 4.5005
R79693 VDD.n1313 VDD.n1214 4.5005
R79694 VDD.n1379 VDD.n1214 4.5005
R79695 VDD.n1312 VDD.n1214 4.5005
R79696 VDD.n1380 VDD.n1214 4.5005
R79697 VDD.n1310 VDD.n1214 4.5005
R79698 VDD.n1381 VDD.n1214 4.5005
R79699 VDD.n1309 VDD.n1214 4.5005
R79700 VDD.n1382 VDD.n1214 4.5005
R79701 VDD.n1307 VDD.n1214 4.5005
R79702 VDD.n1383 VDD.n1214 4.5005
R79703 VDD.n1306 VDD.n1214 4.5005
R79704 VDD.n1384 VDD.n1214 4.5005
R79705 VDD.n1304 VDD.n1214 4.5005
R79706 VDD.n1385 VDD.n1214 4.5005
R79707 VDD.n1303 VDD.n1214 4.5005
R79708 VDD.n1386 VDD.n1214 4.5005
R79709 VDD.n1301 VDD.n1214 4.5005
R79710 VDD.n1387 VDD.n1214 4.5005
R79711 VDD.n1300 VDD.n1214 4.5005
R79712 VDD.n1388 VDD.n1214 4.5005
R79713 VDD.n1298 VDD.n1214 4.5005
R79714 VDD.n1389 VDD.n1214 4.5005
R79715 VDD.n1297 VDD.n1214 4.5005
R79716 VDD.n1390 VDD.n1214 4.5005
R79717 VDD.n1295 VDD.n1214 4.5005
R79718 VDD.n1391 VDD.n1214 4.5005
R79719 VDD.n1294 VDD.n1214 4.5005
R79720 VDD.n1392 VDD.n1214 4.5005
R79721 VDD.n1292 VDD.n1214 4.5005
R79722 VDD.n1393 VDD.n1214 4.5005
R79723 VDD.n1291 VDD.n1214 4.5005
R79724 VDD.n1394 VDD.n1214 4.5005
R79725 VDD.n1289 VDD.n1214 4.5005
R79726 VDD.n1395 VDD.n1214 4.5005
R79727 VDD.n1288 VDD.n1214 4.5005
R79728 VDD.n1396 VDD.n1214 4.5005
R79729 VDD.n1286 VDD.n1214 4.5005
R79730 VDD.n1397 VDD.n1214 4.5005
R79731 VDD.n1285 VDD.n1214 4.5005
R79732 VDD.n1398 VDD.n1214 4.5005
R79733 VDD.n1283 VDD.n1214 4.5005
R79734 VDD.n1399 VDD.n1214 4.5005
R79735 VDD.n1282 VDD.n1214 4.5005
R79736 VDD.n1400 VDD.n1214 4.5005
R79737 VDD.n1280 VDD.n1214 4.5005
R79738 VDD.n1401 VDD.n1214 4.5005
R79739 VDD.n1279 VDD.n1214 4.5005
R79740 VDD.n1402 VDD.n1214 4.5005
R79741 VDD.n1277 VDD.n1214 4.5005
R79742 VDD.n1403 VDD.n1214 4.5005
R79743 VDD.n1276 VDD.n1214 4.5005
R79744 VDD.n1404 VDD.n1214 4.5005
R79745 VDD.n1274 VDD.n1214 4.5005
R79746 VDD.n1405 VDD.n1214 4.5005
R79747 VDD.n1273 VDD.n1214 4.5005
R79748 VDD.n1406 VDD.n1214 4.5005
R79749 VDD.n1271 VDD.n1214 4.5005
R79750 VDD.n1407 VDD.n1214 4.5005
R79751 VDD.n1270 VDD.n1214 4.5005
R79752 VDD.n1408 VDD.n1214 4.5005
R79753 VDD.n1268 VDD.n1214 4.5005
R79754 VDD.n1409 VDD.n1214 4.5005
R79755 VDD.n1267 VDD.n1214 4.5005
R79756 VDD.n1410 VDD.n1214 4.5005
R79757 VDD.n1265 VDD.n1214 4.5005
R79758 VDD.n1411 VDD.n1214 4.5005
R79759 VDD.n1264 VDD.n1214 4.5005
R79760 VDD.n1412 VDD.n1214 4.5005
R79761 VDD.n1262 VDD.n1214 4.5005
R79762 VDD.n1413 VDD.n1214 4.5005
R79763 VDD.n1261 VDD.n1214 4.5005
R79764 VDD.n1414 VDD.n1214 4.5005
R79765 VDD.n1415 VDD.n1214 4.5005
R79766 VDD.n1674 VDD.n1214 4.5005
R79767 VDD.n1676 VDD.n1175 4.5005
R79768 VDD.n1341 VDD.n1175 4.5005
R79769 VDD.n1342 VDD.n1175 4.5005
R79770 VDD.n1340 VDD.n1175 4.5005
R79771 VDD.n1344 VDD.n1175 4.5005
R79772 VDD.n1339 VDD.n1175 4.5005
R79773 VDD.n1345 VDD.n1175 4.5005
R79774 VDD.n1338 VDD.n1175 4.5005
R79775 VDD.n1347 VDD.n1175 4.5005
R79776 VDD.n1337 VDD.n1175 4.5005
R79777 VDD.n1348 VDD.n1175 4.5005
R79778 VDD.n1336 VDD.n1175 4.5005
R79779 VDD.n1350 VDD.n1175 4.5005
R79780 VDD.n1335 VDD.n1175 4.5005
R79781 VDD.n1351 VDD.n1175 4.5005
R79782 VDD.n1334 VDD.n1175 4.5005
R79783 VDD.n1353 VDD.n1175 4.5005
R79784 VDD.n1333 VDD.n1175 4.5005
R79785 VDD.n1354 VDD.n1175 4.5005
R79786 VDD.n1332 VDD.n1175 4.5005
R79787 VDD.n1356 VDD.n1175 4.5005
R79788 VDD.n1331 VDD.n1175 4.5005
R79789 VDD.n1357 VDD.n1175 4.5005
R79790 VDD.n1330 VDD.n1175 4.5005
R79791 VDD.n1359 VDD.n1175 4.5005
R79792 VDD.n1329 VDD.n1175 4.5005
R79793 VDD.n1360 VDD.n1175 4.5005
R79794 VDD.n1328 VDD.n1175 4.5005
R79795 VDD.n1362 VDD.n1175 4.5005
R79796 VDD.n1327 VDD.n1175 4.5005
R79797 VDD.n1363 VDD.n1175 4.5005
R79798 VDD.n1326 VDD.n1175 4.5005
R79799 VDD.n1365 VDD.n1175 4.5005
R79800 VDD.n1325 VDD.n1175 4.5005
R79801 VDD.n1366 VDD.n1175 4.5005
R79802 VDD.n1324 VDD.n1175 4.5005
R79803 VDD.n1368 VDD.n1175 4.5005
R79804 VDD.n1323 VDD.n1175 4.5005
R79805 VDD.n1369 VDD.n1175 4.5005
R79806 VDD.n1322 VDD.n1175 4.5005
R79807 VDD.n1371 VDD.n1175 4.5005
R79808 VDD.n1321 VDD.n1175 4.5005
R79809 VDD.n1372 VDD.n1175 4.5005
R79810 VDD.n1320 VDD.n1175 4.5005
R79811 VDD.n1374 VDD.n1175 4.5005
R79812 VDD.n1319 VDD.n1175 4.5005
R79813 VDD.n1375 VDD.n1175 4.5005
R79814 VDD.n1318 VDD.n1175 4.5005
R79815 VDD.n1376 VDD.n1175 4.5005
R79816 VDD.n1316 VDD.n1175 4.5005
R79817 VDD.n1377 VDD.n1175 4.5005
R79818 VDD.n1315 VDD.n1175 4.5005
R79819 VDD.n1378 VDD.n1175 4.5005
R79820 VDD.n1313 VDD.n1175 4.5005
R79821 VDD.n1379 VDD.n1175 4.5005
R79822 VDD.n1312 VDD.n1175 4.5005
R79823 VDD.n1380 VDD.n1175 4.5005
R79824 VDD.n1310 VDD.n1175 4.5005
R79825 VDD.n1381 VDD.n1175 4.5005
R79826 VDD.n1309 VDD.n1175 4.5005
R79827 VDD.n1382 VDD.n1175 4.5005
R79828 VDD.n1307 VDD.n1175 4.5005
R79829 VDD.n1383 VDD.n1175 4.5005
R79830 VDD.n1306 VDD.n1175 4.5005
R79831 VDD.n1384 VDD.n1175 4.5005
R79832 VDD.n1304 VDD.n1175 4.5005
R79833 VDD.n1385 VDD.n1175 4.5005
R79834 VDD.n1303 VDD.n1175 4.5005
R79835 VDD.n1386 VDD.n1175 4.5005
R79836 VDD.n1301 VDD.n1175 4.5005
R79837 VDD.n1387 VDD.n1175 4.5005
R79838 VDD.n1300 VDD.n1175 4.5005
R79839 VDD.n1388 VDD.n1175 4.5005
R79840 VDD.n1298 VDD.n1175 4.5005
R79841 VDD.n1389 VDD.n1175 4.5005
R79842 VDD.n1297 VDD.n1175 4.5005
R79843 VDD.n1390 VDD.n1175 4.5005
R79844 VDD.n1295 VDD.n1175 4.5005
R79845 VDD.n1391 VDD.n1175 4.5005
R79846 VDD.n1294 VDD.n1175 4.5005
R79847 VDD.n1392 VDD.n1175 4.5005
R79848 VDD.n1292 VDD.n1175 4.5005
R79849 VDD.n1393 VDD.n1175 4.5005
R79850 VDD.n1291 VDD.n1175 4.5005
R79851 VDD.n1394 VDD.n1175 4.5005
R79852 VDD.n1289 VDD.n1175 4.5005
R79853 VDD.n1395 VDD.n1175 4.5005
R79854 VDD.n1288 VDD.n1175 4.5005
R79855 VDD.n1396 VDD.n1175 4.5005
R79856 VDD.n1286 VDD.n1175 4.5005
R79857 VDD.n1397 VDD.n1175 4.5005
R79858 VDD.n1285 VDD.n1175 4.5005
R79859 VDD.n1398 VDD.n1175 4.5005
R79860 VDD.n1283 VDD.n1175 4.5005
R79861 VDD.n1399 VDD.n1175 4.5005
R79862 VDD.n1282 VDD.n1175 4.5005
R79863 VDD.n1400 VDD.n1175 4.5005
R79864 VDD.n1280 VDD.n1175 4.5005
R79865 VDD.n1401 VDD.n1175 4.5005
R79866 VDD.n1279 VDD.n1175 4.5005
R79867 VDD.n1402 VDD.n1175 4.5005
R79868 VDD.n1277 VDD.n1175 4.5005
R79869 VDD.n1403 VDD.n1175 4.5005
R79870 VDD.n1276 VDD.n1175 4.5005
R79871 VDD.n1404 VDD.n1175 4.5005
R79872 VDD.n1274 VDD.n1175 4.5005
R79873 VDD.n1405 VDD.n1175 4.5005
R79874 VDD.n1273 VDD.n1175 4.5005
R79875 VDD.n1406 VDD.n1175 4.5005
R79876 VDD.n1271 VDD.n1175 4.5005
R79877 VDD.n1407 VDD.n1175 4.5005
R79878 VDD.n1270 VDD.n1175 4.5005
R79879 VDD.n1408 VDD.n1175 4.5005
R79880 VDD.n1268 VDD.n1175 4.5005
R79881 VDD.n1409 VDD.n1175 4.5005
R79882 VDD.n1267 VDD.n1175 4.5005
R79883 VDD.n1410 VDD.n1175 4.5005
R79884 VDD.n1265 VDD.n1175 4.5005
R79885 VDD.n1411 VDD.n1175 4.5005
R79886 VDD.n1264 VDD.n1175 4.5005
R79887 VDD.n1412 VDD.n1175 4.5005
R79888 VDD.n1262 VDD.n1175 4.5005
R79889 VDD.n1413 VDD.n1175 4.5005
R79890 VDD.n1261 VDD.n1175 4.5005
R79891 VDD.n1414 VDD.n1175 4.5005
R79892 VDD.n1415 VDD.n1175 4.5005
R79893 VDD.n1674 VDD.n1175 4.5005
R79894 VDD.n1676 VDD.n1215 4.5005
R79895 VDD.n1341 VDD.n1215 4.5005
R79896 VDD.n1342 VDD.n1215 4.5005
R79897 VDD.n1340 VDD.n1215 4.5005
R79898 VDD.n1344 VDD.n1215 4.5005
R79899 VDD.n1339 VDD.n1215 4.5005
R79900 VDD.n1345 VDD.n1215 4.5005
R79901 VDD.n1338 VDD.n1215 4.5005
R79902 VDD.n1347 VDD.n1215 4.5005
R79903 VDD.n1337 VDD.n1215 4.5005
R79904 VDD.n1348 VDD.n1215 4.5005
R79905 VDD.n1336 VDD.n1215 4.5005
R79906 VDD.n1350 VDD.n1215 4.5005
R79907 VDD.n1335 VDD.n1215 4.5005
R79908 VDD.n1351 VDD.n1215 4.5005
R79909 VDD.n1334 VDD.n1215 4.5005
R79910 VDD.n1353 VDD.n1215 4.5005
R79911 VDD.n1333 VDD.n1215 4.5005
R79912 VDD.n1354 VDD.n1215 4.5005
R79913 VDD.n1332 VDD.n1215 4.5005
R79914 VDD.n1356 VDD.n1215 4.5005
R79915 VDD.n1331 VDD.n1215 4.5005
R79916 VDD.n1357 VDD.n1215 4.5005
R79917 VDD.n1330 VDD.n1215 4.5005
R79918 VDD.n1359 VDD.n1215 4.5005
R79919 VDD.n1329 VDD.n1215 4.5005
R79920 VDD.n1360 VDD.n1215 4.5005
R79921 VDD.n1328 VDD.n1215 4.5005
R79922 VDD.n1362 VDD.n1215 4.5005
R79923 VDD.n1327 VDD.n1215 4.5005
R79924 VDD.n1363 VDD.n1215 4.5005
R79925 VDD.n1326 VDD.n1215 4.5005
R79926 VDD.n1365 VDD.n1215 4.5005
R79927 VDD.n1325 VDD.n1215 4.5005
R79928 VDD.n1366 VDD.n1215 4.5005
R79929 VDD.n1324 VDD.n1215 4.5005
R79930 VDD.n1368 VDD.n1215 4.5005
R79931 VDD.n1323 VDD.n1215 4.5005
R79932 VDD.n1369 VDD.n1215 4.5005
R79933 VDD.n1322 VDD.n1215 4.5005
R79934 VDD.n1371 VDD.n1215 4.5005
R79935 VDD.n1321 VDD.n1215 4.5005
R79936 VDD.n1372 VDD.n1215 4.5005
R79937 VDD.n1320 VDD.n1215 4.5005
R79938 VDD.n1374 VDD.n1215 4.5005
R79939 VDD.n1319 VDD.n1215 4.5005
R79940 VDD.n1375 VDD.n1215 4.5005
R79941 VDD.n1318 VDD.n1215 4.5005
R79942 VDD.n1376 VDD.n1215 4.5005
R79943 VDD.n1316 VDD.n1215 4.5005
R79944 VDD.n1377 VDD.n1215 4.5005
R79945 VDD.n1315 VDD.n1215 4.5005
R79946 VDD.n1378 VDD.n1215 4.5005
R79947 VDD.n1313 VDD.n1215 4.5005
R79948 VDD.n1379 VDD.n1215 4.5005
R79949 VDD.n1312 VDD.n1215 4.5005
R79950 VDD.n1380 VDD.n1215 4.5005
R79951 VDD.n1310 VDD.n1215 4.5005
R79952 VDD.n1381 VDD.n1215 4.5005
R79953 VDD.n1309 VDD.n1215 4.5005
R79954 VDD.n1382 VDD.n1215 4.5005
R79955 VDD.n1307 VDD.n1215 4.5005
R79956 VDD.n1383 VDD.n1215 4.5005
R79957 VDD.n1306 VDD.n1215 4.5005
R79958 VDD.n1384 VDD.n1215 4.5005
R79959 VDD.n1304 VDD.n1215 4.5005
R79960 VDD.n1385 VDD.n1215 4.5005
R79961 VDD.n1303 VDD.n1215 4.5005
R79962 VDD.n1386 VDD.n1215 4.5005
R79963 VDD.n1301 VDD.n1215 4.5005
R79964 VDD.n1387 VDD.n1215 4.5005
R79965 VDD.n1300 VDD.n1215 4.5005
R79966 VDD.n1388 VDD.n1215 4.5005
R79967 VDD.n1298 VDD.n1215 4.5005
R79968 VDD.n1389 VDD.n1215 4.5005
R79969 VDD.n1297 VDD.n1215 4.5005
R79970 VDD.n1390 VDD.n1215 4.5005
R79971 VDD.n1295 VDD.n1215 4.5005
R79972 VDD.n1391 VDD.n1215 4.5005
R79973 VDD.n1294 VDD.n1215 4.5005
R79974 VDD.n1392 VDD.n1215 4.5005
R79975 VDD.n1292 VDD.n1215 4.5005
R79976 VDD.n1393 VDD.n1215 4.5005
R79977 VDD.n1291 VDD.n1215 4.5005
R79978 VDD.n1394 VDD.n1215 4.5005
R79979 VDD.n1289 VDD.n1215 4.5005
R79980 VDD.n1395 VDD.n1215 4.5005
R79981 VDD.n1288 VDD.n1215 4.5005
R79982 VDD.n1396 VDD.n1215 4.5005
R79983 VDD.n1286 VDD.n1215 4.5005
R79984 VDD.n1397 VDD.n1215 4.5005
R79985 VDD.n1285 VDD.n1215 4.5005
R79986 VDD.n1398 VDD.n1215 4.5005
R79987 VDD.n1283 VDD.n1215 4.5005
R79988 VDD.n1399 VDD.n1215 4.5005
R79989 VDD.n1282 VDD.n1215 4.5005
R79990 VDD.n1400 VDD.n1215 4.5005
R79991 VDD.n1280 VDD.n1215 4.5005
R79992 VDD.n1401 VDD.n1215 4.5005
R79993 VDD.n1279 VDD.n1215 4.5005
R79994 VDD.n1402 VDD.n1215 4.5005
R79995 VDD.n1277 VDD.n1215 4.5005
R79996 VDD.n1403 VDD.n1215 4.5005
R79997 VDD.n1276 VDD.n1215 4.5005
R79998 VDD.n1404 VDD.n1215 4.5005
R79999 VDD.n1274 VDD.n1215 4.5005
R80000 VDD.n1405 VDD.n1215 4.5005
R80001 VDD.n1273 VDD.n1215 4.5005
R80002 VDD.n1406 VDD.n1215 4.5005
R80003 VDD.n1271 VDD.n1215 4.5005
R80004 VDD.n1407 VDD.n1215 4.5005
R80005 VDD.n1270 VDD.n1215 4.5005
R80006 VDD.n1408 VDD.n1215 4.5005
R80007 VDD.n1268 VDD.n1215 4.5005
R80008 VDD.n1409 VDD.n1215 4.5005
R80009 VDD.n1267 VDD.n1215 4.5005
R80010 VDD.n1410 VDD.n1215 4.5005
R80011 VDD.n1265 VDD.n1215 4.5005
R80012 VDD.n1411 VDD.n1215 4.5005
R80013 VDD.n1264 VDD.n1215 4.5005
R80014 VDD.n1412 VDD.n1215 4.5005
R80015 VDD.n1262 VDD.n1215 4.5005
R80016 VDD.n1413 VDD.n1215 4.5005
R80017 VDD.n1261 VDD.n1215 4.5005
R80018 VDD.n1414 VDD.n1215 4.5005
R80019 VDD.n1415 VDD.n1215 4.5005
R80020 VDD.n1674 VDD.n1215 4.5005
R80021 VDD.n1676 VDD.n1174 4.5005
R80022 VDD.n1341 VDD.n1174 4.5005
R80023 VDD.n1342 VDD.n1174 4.5005
R80024 VDD.n1340 VDD.n1174 4.5005
R80025 VDD.n1344 VDD.n1174 4.5005
R80026 VDD.n1339 VDD.n1174 4.5005
R80027 VDD.n1345 VDD.n1174 4.5005
R80028 VDD.n1338 VDD.n1174 4.5005
R80029 VDD.n1347 VDD.n1174 4.5005
R80030 VDD.n1337 VDD.n1174 4.5005
R80031 VDD.n1348 VDD.n1174 4.5005
R80032 VDD.n1336 VDD.n1174 4.5005
R80033 VDD.n1350 VDD.n1174 4.5005
R80034 VDD.n1335 VDD.n1174 4.5005
R80035 VDD.n1351 VDD.n1174 4.5005
R80036 VDD.n1334 VDD.n1174 4.5005
R80037 VDD.n1353 VDD.n1174 4.5005
R80038 VDD.n1333 VDD.n1174 4.5005
R80039 VDD.n1354 VDD.n1174 4.5005
R80040 VDD.n1332 VDD.n1174 4.5005
R80041 VDD.n1356 VDD.n1174 4.5005
R80042 VDD.n1331 VDD.n1174 4.5005
R80043 VDD.n1357 VDD.n1174 4.5005
R80044 VDD.n1330 VDD.n1174 4.5005
R80045 VDD.n1359 VDD.n1174 4.5005
R80046 VDD.n1329 VDD.n1174 4.5005
R80047 VDD.n1360 VDD.n1174 4.5005
R80048 VDD.n1328 VDD.n1174 4.5005
R80049 VDD.n1362 VDD.n1174 4.5005
R80050 VDD.n1327 VDD.n1174 4.5005
R80051 VDD.n1363 VDD.n1174 4.5005
R80052 VDD.n1326 VDD.n1174 4.5005
R80053 VDD.n1365 VDD.n1174 4.5005
R80054 VDD.n1325 VDD.n1174 4.5005
R80055 VDD.n1366 VDD.n1174 4.5005
R80056 VDD.n1324 VDD.n1174 4.5005
R80057 VDD.n1368 VDD.n1174 4.5005
R80058 VDD.n1323 VDD.n1174 4.5005
R80059 VDD.n1369 VDD.n1174 4.5005
R80060 VDD.n1322 VDD.n1174 4.5005
R80061 VDD.n1371 VDD.n1174 4.5005
R80062 VDD.n1321 VDD.n1174 4.5005
R80063 VDD.n1372 VDD.n1174 4.5005
R80064 VDD.n1320 VDD.n1174 4.5005
R80065 VDD.n1374 VDD.n1174 4.5005
R80066 VDD.n1319 VDD.n1174 4.5005
R80067 VDD.n1375 VDD.n1174 4.5005
R80068 VDD.n1318 VDD.n1174 4.5005
R80069 VDD.n1376 VDD.n1174 4.5005
R80070 VDD.n1316 VDD.n1174 4.5005
R80071 VDD.n1377 VDD.n1174 4.5005
R80072 VDD.n1315 VDD.n1174 4.5005
R80073 VDD.n1378 VDD.n1174 4.5005
R80074 VDD.n1313 VDD.n1174 4.5005
R80075 VDD.n1379 VDD.n1174 4.5005
R80076 VDD.n1312 VDD.n1174 4.5005
R80077 VDD.n1380 VDD.n1174 4.5005
R80078 VDD.n1310 VDD.n1174 4.5005
R80079 VDD.n1381 VDD.n1174 4.5005
R80080 VDD.n1309 VDD.n1174 4.5005
R80081 VDD.n1382 VDD.n1174 4.5005
R80082 VDD.n1307 VDD.n1174 4.5005
R80083 VDD.n1383 VDD.n1174 4.5005
R80084 VDD.n1306 VDD.n1174 4.5005
R80085 VDD.n1384 VDD.n1174 4.5005
R80086 VDD.n1304 VDD.n1174 4.5005
R80087 VDD.n1385 VDD.n1174 4.5005
R80088 VDD.n1303 VDD.n1174 4.5005
R80089 VDD.n1386 VDD.n1174 4.5005
R80090 VDD.n1301 VDD.n1174 4.5005
R80091 VDD.n1387 VDD.n1174 4.5005
R80092 VDD.n1300 VDD.n1174 4.5005
R80093 VDD.n1388 VDD.n1174 4.5005
R80094 VDD.n1298 VDD.n1174 4.5005
R80095 VDD.n1389 VDD.n1174 4.5005
R80096 VDD.n1297 VDD.n1174 4.5005
R80097 VDD.n1390 VDD.n1174 4.5005
R80098 VDD.n1295 VDD.n1174 4.5005
R80099 VDD.n1391 VDD.n1174 4.5005
R80100 VDD.n1294 VDD.n1174 4.5005
R80101 VDD.n1392 VDD.n1174 4.5005
R80102 VDD.n1292 VDD.n1174 4.5005
R80103 VDD.n1393 VDD.n1174 4.5005
R80104 VDD.n1291 VDD.n1174 4.5005
R80105 VDD.n1394 VDD.n1174 4.5005
R80106 VDD.n1289 VDD.n1174 4.5005
R80107 VDD.n1395 VDD.n1174 4.5005
R80108 VDD.n1288 VDD.n1174 4.5005
R80109 VDD.n1396 VDD.n1174 4.5005
R80110 VDD.n1286 VDD.n1174 4.5005
R80111 VDD.n1397 VDD.n1174 4.5005
R80112 VDD.n1285 VDD.n1174 4.5005
R80113 VDD.n1398 VDD.n1174 4.5005
R80114 VDD.n1283 VDD.n1174 4.5005
R80115 VDD.n1399 VDD.n1174 4.5005
R80116 VDD.n1282 VDD.n1174 4.5005
R80117 VDD.n1400 VDD.n1174 4.5005
R80118 VDD.n1280 VDD.n1174 4.5005
R80119 VDD.n1401 VDD.n1174 4.5005
R80120 VDD.n1279 VDD.n1174 4.5005
R80121 VDD.n1402 VDD.n1174 4.5005
R80122 VDD.n1277 VDD.n1174 4.5005
R80123 VDD.n1403 VDD.n1174 4.5005
R80124 VDD.n1276 VDD.n1174 4.5005
R80125 VDD.n1404 VDD.n1174 4.5005
R80126 VDD.n1274 VDD.n1174 4.5005
R80127 VDD.n1405 VDD.n1174 4.5005
R80128 VDD.n1273 VDD.n1174 4.5005
R80129 VDD.n1406 VDD.n1174 4.5005
R80130 VDD.n1271 VDD.n1174 4.5005
R80131 VDD.n1407 VDD.n1174 4.5005
R80132 VDD.n1270 VDD.n1174 4.5005
R80133 VDD.n1408 VDD.n1174 4.5005
R80134 VDD.n1268 VDD.n1174 4.5005
R80135 VDD.n1409 VDD.n1174 4.5005
R80136 VDD.n1267 VDD.n1174 4.5005
R80137 VDD.n1410 VDD.n1174 4.5005
R80138 VDD.n1265 VDD.n1174 4.5005
R80139 VDD.n1411 VDD.n1174 4.5005
R80140 VDD.n1264 VDD.n1174 4.5005
R80141 VDD.n1412 VDD.n1174 4.5005
R80142 VDD.n1262 VDD.n1174 4.5005
R80143 VDD.n1413 VDD.n1174 4.5005
R80144 VDD.n1261 VDD.n1174 4.5005
R80145 VDD.n1414 VDD.n1174 4.5005
R80146 VDD.n1415 VDD.n1174 4.5005
R80147 VDD.n1674 VDD.n1174 4.5005
R80148 VDD.n1676 VDD.n1216 4.5005
R80149 VDD.n1341 VDD.n1216 4.5005
R80150 VDD.n1342 VDD.n1216 4.5005
R80151 VDD.n1340 VDD.n1216 4.5005
R80152 VDD.n1344 VDD.n1216 4.5005
R80153 VDD.n1339 VDD.n1216 4.5005
R80154 VDD.n1345 VDD.n1216 4.5005
R80155 VDD.n1338 VDD.n1216 4.5005
R80156 VDD.n1347 VDD.n1216 4.5005
R80157 VDD.n1337 VDD.n1216 4.5005
R80158 VDD.n1348 VDD.n1216 4.5005
R80159 VDD.n1336 VDD.n1216 4.5005
R80160 VDD.n1350 VDD.n1216 4.5005
R80161 VDD.n1335 VDD.n1216 4.5005
R80162 VDD.n1351 VDD.n1216 4.5005
R80163 VDD.n1334 VDD.n1216 4.5005
R80164 VDD.n1353 VDD.n1216 4.5005
R80165 VDD.n1333 VDD.n1216 4.5005
R80166 VDD.n1354 VDD.n1216 4.5005
R80167 VDD.n1332 VDD.n1216 4.5005
R80168 VDD.n1356 VDD.n1216 4.5005
R80169 VDD.n1331 VDD.n1216 4.5005
R80170 VDD.n1357 VDD.n1216 4.5005
R80171 VDD.n1330 VDD.n1216 4.5005
R80172 VDD.n1359 VDD.n1216 4.5005
R80173 VDD.n1329 VDD.n1216 4.5005
R80174 VDD.n1360 VDD.n1216 4.5005
R80175 VDD.n1328 VDD.n1216 4.5005
R80176 VDD.n1362 VDD.n1216 4.5005
R80177 VDD.n1327 VDD.n1216 4.5005
R80178 VDD.n1363 VDD.n1216 4.5005
R80179 VDD.n1326 VDD.n1216 4.5005
R80180 VDD.n1365 VDD.n1216 4.5005
R80181 VDD.n1325 VDD.n1216 4.5005
R80182 VDD.n1366 VDD.n1216 4.5005
R80183 VDD.n1324 VDD.n1216 4.5005
R80184 VDD.n1368 VDD.n1216 4.5005
R80185 VDD.n1323 VDD.n1216 4.5005
R80186 VDD.n1369 VDD.n1216 4.5005
R80187 VDD.n1322 VDD.n1216 4.5005
R80188 VDD.n1371 VDD.n1216 4.5005
R80189 VDD.n1321 VDD.n1216 4.5005
R80190 VDD.n1372 VDD.n1216 4.5005
R80191 VDD.n1320 VDD.n1216 4.5005
R80192 VDD.n1374 VDD.n1216 4.5005
R80193 VDD.n1319 VDD.n1216 4.5005
R80194 VDD.n1375 VDD.n1216 4.5005
R80195 VDD.n1318 VDD.n1216 4.5005
R80196 VDD.n1376 VDD.n1216 4.5005
R80197 VDD.n1316 VDD.n1216 4.5005
R80198 VDD.n1377 VDD.n1216 4.5005
R80199 VDD.n1315 VDD.n1216 4.5005
R80200 VDD.n1378 VDD.n1216 4.5005
R80201 VDD.n1313 VDD.n1216 4.5005
R80202 VDD.n1379 VDD.n1216 4.5005
R80203 VDD.n1312 VDD.n1216 4.5005
R80204 VDD.n1380 VDD.n1216 4.5005
R80205 VDD.n1310 VDD.n1216 4.5005
R80206 VDD.n1381 VDD.n1216 4.5005
R80207 VDD.n1309 VDD.n1216 4.5005
R80208 VDD.n1382 VDD.n1216 4.5005
R80209 VDD.n1307 VDD.n1216 4.5005
R80210 VDD.n1383 VDD.n1216 4.5005
R80211 VDD.n1306 VDD.n1216 4.5005
R80212 VDD.n1384 VDD.n1216 4.5005
R80213 VDD.n1304 VDD.n1216 4.5005
R80214 VDD.n1385 VDD.n1216 4.5005
R80215 VDD.n1303 VDD.n1216 4.5005
R80216 VDD.n1386 VDD.n1216 4.5005
R80217 VDD.n1301 VDD.n1216 4.5005
R80218 VDD.n1387 VDD.n1216 4.5005
R80219 VDD.n1300 VDD.n1216 4.5005
R80220 VDD.n1388 VDD.n1216 4.5005
R80221 VDD.n1298 VDD.n1216 4.5005
R80222 VDD.n1389 VDD.n1216 4.5005
R80223 VDD.n1297 VDD.n1216 4.5005
R80224 VDD.n1390 VDD.n1216 4.5005
R80225 VDD.n1295 VDD.n1216 4.5005
R80226 VDD.n1391 VDD.n1216 4.5005
R80227 VDD.n1294 VDD.n1216 4.5005
R80228 VDD.n1392 VDD.n1216 4.5005
R80229 VDD.n1292 VDD.n1216 4.5005
R80230 VDD.n1393 VDD.n1216 4.5005
R80231 VDD.n1291 VDD.n1216 4.5005
R80232 VDD.n1394 VDD.n1216 4.5005
R80233 VDD.n1289 VDD.n1216 4.5005
R80234 VDD.n1395 VDD.n1216 4.5005
R80235 VDD.n1288 VDD.n1216 4.5005
R80236 VDD.n1396 VDD.n1216 4.5005
R80237 VDD.n1286 VDD.n1216 4.5005
R80238 VDD.n1397 VDD.n1216 4.5005
R80239 VDD.n1285 VDD.n1216 4.5005
R80240 VDD.n1398 VDD.n1216 4.5005
R80241 VDD.n1283 VDD.n1216 4.5005
R80242 VDD.n1399 VDD.n1216 4.5005
R80243 VDD.n1282 VDD.n1216 4.5005
R80244 VDD.n1400 VDD.n1216 4.5005
R80245 VDD.n1280 VDD.n1216 4.5005
R80246 VDD.n1401 VDD.n1216 4.5005
R80247 VDD.n1279 VDD.n1216 4.5005
R80248 VDD.n1402 VDD.n1216 4.5005
R80249 VDD.n1277 VDD.n1216 4.5005
R80250 VDD.n1403 VDD.n1216 4.5005
R80251 VDD.n1276 VDD.n1216 4.5005
R80252 VDD.n1404 VDD.n1216 4.5005
R80253 VDD.n1274 VDD.n1216 4.5005
R80254 VDD.n1405 VDD.n1216 4.5005
R80255 VDD.n1273 VDD.n1216 4.5005
R80256 VDD.n1406 VDD.n1216 4.5005
R80257 VDD.n1271 VDD.n1216 4.5005
R80258 VDD.n1407 VDD.n1216 4.5005
R80259 VDD.n1270 VDD.n1216 4.5005
R80260 VDD.n1408 VDD.n1216 4.5005
R80261 VDD.n1268 VDD.n1216 4.5005
R80262 VDD.n1409 VDD.n1216 4.5005
R80263 VDD.n1267 VDD.n1216 4.5005
R80264 VDD.n1410 VDD.n1216 4.5005
R80265 VDD.n1265 VDD.n1216 4.5005
R80266 VDD.n1411 VDD.n1216 4.5005
R80267 VDD.n1264 VDD.n1216 4.5005
R80268 VDD.n1412 VDD.n1216 4.5005
R80269 VDD.n1262 VDD.n1216 4.5005
R80270 VDD.n1413 VDD.n1216 4.5005
R80271 VDD.n1261 VDD.n1216 4.5005
R80272 VDD.n1414 VDD.n1216 4.5005
R80273 VDD.n1415 VDD.n1216 4.5005
R80274 VDD.n1674 VDD.n1216 4.5005
R80275 VDD.n1676 VDD.n1173 4.5005
R80276 VDD.n1341 VDD.n1173 4.5005
R80277 VDD.n1342 VDD.n1173 4.5005
R80278 VDD.n1340 VDD.n1173 4.5005
R80279 VDD.n1344 VDD.n1173 4.5005
R80280 VDD.n1339 VDD.n1173 4.5005
R80281 VDD.n1345 VDD.n1173 4.5005
R80282 VDD.n1338 VDD.n1173 4.5005
R80283 VDD.n1347 VDD.n1173 4.5005
R80284 VDD.n1337 VDD.n1173 4.5005
R80285 VDD.n1348 VDD.n1173 4.5005
R80286 VDD.n1336 VDD.n1173 4.5005
R80287 VDD.n1350 VDD.n1173 4.5005
R80288 VDD.n1335 VDD.n1173 4.5005
R80289 VDD.n1351 VDD.n1173 4.5005
R80290 VDD.n1334 VDD.n1173 4.5005
R80291 VDD.n1353 VDD.n1173 4.5005
R80292 VDD.n1333 VDD.n1173 4.5005
R80293 VDD.n1354 VDD.n1173 4.5005
R80294 VDD.n1332 VDD.n1173 4.5005
R80295 VDD.n1356 VDD.n1173 4.5005
R80296 VDD.n1331 VDD.n1173 4.5005
R80297 VDD.n1357 VDD.n1173 4.5005
R80298 VDD.n1330 VDD.n1173 4.5005
R80299 VDD.n1359 VDD.n1173 4.5005
R80300 VDD.n1329 VDD.n1173 4.5005
R80301 VDD.n1360 VDD.n1173 4.5005
R80302 VDD.n1328 VDD.n1173 4.5005
R80303 VDD.n1362 VDD.n1173 4.5005
R80304 VDD.n1327 VDD.n1173 4.5005
R80305 VDD.n1363 VDD.n1173 4.5005
R80306 VDD.n1326 VDD.n1173 4.5005
R80307 VDD.n1365 VDD.n1173 4.5005
R80308 VDD.n1325 VDD.n1173 4.5005
R80309 VDD.n1366 VDD.n1173 4.5005
R80310 VDD.n1324 VDD.n1173 4.5005
R80311 VDD.n1368 VDD.n1173 4.5005
R80312 VDD.n1323 VDD.n1173 4.5005
R80313 VDD.n1369 VDD.n1173 4.5005
R80314 VDD.n1322 VDD.n1173 4.5005
R80315 VDD.n1371 VDD.n1173 4.5005
R80316 VDD.n1321 VDD.n1173 4.5005
R80317 VDD.n1372 VDD.n1173 4.5005
R80318 VDD.n1320 VDD.n1173 4.5005
R80319 VDD.n1374 VDD.n1173 4.5005
R80320 VDD.n1319 VDD.n1173 4.5005
R80321 VDD.n1375 VDD.n1173 4.5005
R80322 VDD.n1318 VDD.n1173 4.5005
R80323 VDD.n1376 VDD.n1173 4.5005
R80324 VDD.n1316 VDD.n1173 4.5005
R80325 VDD.n1377 VDD.n1173 4.5005
R80326 VDD.n1315 VDD.n1173 4.5005
R80327 VDD.n1378 VDD.n1173 4.5005
R80328 VDD.n1313 VDD.n1173 4.5005
R80329 VDD.n1379 VDD.n1173 4.5005
R80330 VDD.n1312 VDD.n1173 4.5005
R80331 VDD.n1380 VDD.n1173 4.5005
R80332 VDD.n1310 VDD.n1173 4.5005
R80333 VDD.n1381 VDD.n1173 4.5005
R80334 VDD.n1309 VDD.n1173 4.5005
R80335 VDD.n1382 VDD.n1173 4.5005
R80336 VDD.n1307 VDD.n1173 4.5005
R80337 VDD.n1383 VDD.n1173 4.5005
R80338 VDD.n1306 VDD.n1173 4.5005
R80339 VDD.n1384 VDD.n1173 4.5005
R80340 VDD.n1304 VDD.n1173 4.5005
R80341 VDD.n1385 VDD.n1173 4.5005
R80342 VDD.n1303 VDD.n1173 4.5005
R80343 VDD.n1386 VDD.n1173 4.5005
R80344 VDD.n1301 VDD.n1173 4.5005
R80345 VDD.n1387 VDD.n1173 4.5005
R80346 VDD.n1300 VDD.n1173 4.5005
R80347 VDD.n1388 VDD.n1173 4.5005
R80348 VDD.n1298 VDD.n1173 4.5005
R80349 VDD.n1389 VDD.n1173 4.5005
R80350 VDD.n1297 VDD.n1173 4.5005
R80351 VDD.n1390 VDD.n1173 4.5005
R80352 VDD.n1295 VDD.n1173 4.5005
R80353 VDD.n1391 VDD.n1173 4.5005
R80354 VDD.n1294 VDD.n1173 4.5005
R80355 VDD.n1392 VDD.n1173 4.5005
R80356 VDD.n1292 VDD.n1173 4.5005
R80357 VDD.n1393 VDD.n1173 4.5005
R80358 VDD.n1291 VDD.n1173 4.5005
R80359 VDD.n1394 VDD.n1173 4.5005
R80360 VDD.n1289 VDD.n1173 4.5005
R80361 VDD.n1395 VDD.n1173 4.5005
R80362 VDD.n1288 VDD.n1173 4.5005
R80363 VDD.n1396 VDD.n1173 4.5005
R80364 VDD.n1286 VDD.n1173 4.5005
R80365 VDD.n1397 VDD.n1173 4.5005
R80366 VDD.n1285 VDD.n1173 4.5005
R80367 VDD.n1398 VDD.n1173 4.5005
R80368 VDD.n1283 VDD.n1173 4.5005
R80369 VDD.n1399 VDD.n1173 4.5005
R80370 VDD.n1282 VDD.n1173 4.5005
R80371 VDD.n1400 VDD.n1173 4.5005
R80372 VDD.n1280 VDD.n1173 4.5005
R80373 VDD.n1401 VDD.n1173 4.5005
R80374 VDD.n1279 VDD.n1173 4.5005
R80375 VDD.n1402 VDD.n1173 4.5005
R80376 VDD.n1277 VDD.n1173 4.5005
R80377 VDD.n1403 VDD.n1173 4.5005
R80378 VDD.n1276 VDD.n1173 4.5005
R80379 VDD.n1404 VDD.n1173 4.5005
R80380 VDD.n1274 VDD.n1173 4.5005
R80381 VDD.n1405 VDD.n1173 4.5005
R80382 VDD.n1273 VDD.n1173 4.5005
R80383 VDD.n1406 VDD.n1173 4.5005
R80384 VDD.n1271 VDD.n1173 4.5005
R80385 VDD.n1407 VDD.n1173 4.5005
R80386 VDD.n1270 VDD.n1173 4.5005
R80387 VDD.n1408 VDD.n1173 4.5005
R80388 VDD.n1268 VDD.n1173 4.5005
R80389 VDD.n1409 VDD.n1173 4.5005
R80390 VDD.n1267 VDD.n1173 4.5005
R80391 VDD.n1410 VDD.n1173 4.5005
R80392 VDD.n1265 VDD.n1173 4.5005
R80393 VDD.n1411 VDD.n1173 4.5005
R80394 VDD.n1264 VDD.n1173 4.5005
R80395 VDD.n1412 VDD.n1173 4.5005
R80396 VDD.n1262 VDD.n1173 4.5005
R80397 VDD.n1413 VDD.n1173 4.5005
R80398 VDD.n1261 VDD.n1173 4.5005
R80399 VDD.n1414 VDD.n1173 4.5005
R80400 VDD.n1415 VDD.n1173 4.5005
R80401 VDD.n1674 VDD.n1173 4.5005
R80402 VDD.n1676 VDD.n1217 4.5005
R80403 VDD.n1341 VDD.n1217 4.5005
R80404 VDD.n1342 VDD.n1217 4.5005
R80405 VDD.n1340 VDD.n1217 4.5005
R80406 VDD.n1344 VDD.n1217 4.5005
R80407 VDD.n1339 VDD.n1217 4.5005
R80408 VDD.n1345 VDD.n1217 4.5005
R80409 VDD.n1338 VDD.n1217 4.5005
R80410 VDD.n1347 VDD.n1217 4.5005
R80411 VDD.n1337 VDD.n1217 4.5005
R80412 VDD.n1348 VDD.n1217 4.5005
R80413 VDD.n1336 VDD.n1217 4.5005
R80414 VDD.n1350 VDD.n1217 4.5005
R80415 VDD.n1335 VDD.n1217 4.5005
R80416 VDD.n1351 VDD.n1217 4.5005
R80417 VDD.n1334 VDD.n1217 4.5005
R80418 VDD.n1353 VDD.n1217 4.5005
R80419 VDD.n1333 VDD.n1217 4.5005
R80420 VDD.n1354 VDD.n1217 4.5005
R80421 VDD.n1332 VDD.n1217 4.5005
R80422 VDD.n1356 VDD.n1217 4.5005
R80423 VDD.n1331 VDD.n1217 4.5005
R80424 VDD.n1357 VDD.n1217 4.5005
R80425 VDD.n1330 VDD.n1217 4.5005
R80426 VDD.n1359 VDD.n1217 4.5005
R80427 VDD.n1329 VDD.n1217 4.5005
R80428 VDD.n1360 VDD.n1217 4.5005
R80429 VDD.n1328 VDD.n1217 4.5005
R80430 VDD.n1362 VDD.n1217 4.5005
R80431 VDD.n1327 VDD.n1217 4.5005
R80432 VDD.n1363 VDD.n1217 4.5005
R80433 VDD.n1326 VDD.n1217 4.5005
R80434 VDD.n1365 VDD.n1217 4.5005
R80435 VDD.n1325 VDD.n1217 4.5005
R80436 VDD.n1366 VDD.n1217 4.5005
R80437 VDD.n1324 VDD.n1217 4.5005
R80438 VDD.n1368 VDD.n1217 4.5005
R80439 VDD.n1323 VDD.n1217 4.5005
R80440 VDD.n1369 VDD.n1217 4.5005
R80441 VDD.n1322 VDD.n1217 4.5005
R80442 VDD.n1371 VDD.n1217 4.5005
R80443 VDD.n1321 VDD.n1217 4.5005
R80444 VDD.n1372 VDD.n1217 4.5005
R80445 VDD.n1320 VDD.n1217 4.5005
R80446 VDD.n1374 VDD.n1217 4.5005
R80447 VDD.n1319 VDD.n1217 4.5005
R80448 VDD.n1375 VDD.n1217 4.5005
R80449 VDD.n1318 VDD.n1217 4.5005
R80450 VDD.n1376 VDD.n1217 4.5005
R80451 VDD.n1316 VDD.n1217 4.5005
R80452 VDD.n1377 VDD.n1217 4.5005
R80453 VDD.n1315 VDD.n1217 4.5005
R80454 VDD.n1378 VDD.n1217 4.5005
R80455 VDD.n1313 VDD.n1217 4.5005
R80456 VDD.n1379 VDD.n1217 4.5005
R80457 VDD.n1312 VDD.n1217 4.5005
R80458 VDD.n1380 VDD.n1217 4.5005
R80459 VDD.n1310 VDD.n1217 4.5005
R80460 VDD.n1381 VDD.n1217 4.5005
R80461 VDD.n1309 VDD.n1217 4.5005
R80462 VDD.n1382 VDD.n1217 4.5005
R80463 VDD.n1307 VDD.n1217 4.5005
R80464 VDD.n1383 VDD.n1217 4.5005
R80465 VDD.n1306 VDD.n1217 4.5005
R80466 VDD.n1384 VDD.n1217 4.5005
R80467 VDD.n1304 VDD.n1217 4.5005
R80468 VDD.n1385 VDD.n1217 4.5005
R80469 VDD.n1303 VDD.n1217 4.5005
R80470 VDD.n1386 VDD.n1217 4.5005
R80471 VDD.n1301 VDD.n1217 4.5005
R80472 VDD.n1387 VDD.n1217 4.5005
R80473 VDD.n1300 VDD.n1217 4.5005
R80474 VDD.n1388 VDD.n1217 4.5005
R80475 VDD.n1298 VDD.n1217 4.5005
R80476 VDD.n1389 VDD.n1217 4.5005
R80477 VDD.n1297 VDD.n1217 4.5005
R80478 VDD.n1390 VDD.n1217 4.5005
R80479 VDD.n1295 VDD.n1217 4.5005
R80480 VDD.n1391 VDD.n1217 4.5005
R80481 VDD.n1294 VDD.n1217 4.5005
R80482 VDD.n1392 VDD.n1217 4.5005
R80483 VDD.n1292 VDD.n1217 4.5005
R80484 VDD.n1393 VDD.n1217 4.5005
R80485 VDD.n1291 VDD.n1217 4.5005
R80486 VDD.n1394 VDD.n1217 4.5005
R80487 VDD.n1289 VDD.n1217 4.5005
R80488 VDD.n1395 VDD.n1217 4.5005
R80489 VDD.n1288 VDD.n1217 4.5005
R80490 VDD.n1396 VDD.n1217 4.5005
R80491 VDD.n1286 VDD.n1217 4.5005
R80492 VDD.n1397 VDD.n1217 4.5005
R80493 VDD.n1285 VDD.n1217 4.5005
R80494 VDD.n1398 VDD.n1217 4.5005
R80495 VDD.n1283 VDD.n1217 4.5005
R80496 VDD.n1399 VDD.n1217 4.5005
R80497 VDD.n1282 VDD.n1217 4.5005
R80498 VDD.n1400 VDD.n1217 4.5005
R80499 VDD.n1280 VDD.n1217 4.5005
R80500 VDD.n1401 VDD.n1217 4.5005
R80501 VDD.n1279 VDD.n1217 4.5005
R80502 VDD.n1402 VDD.n1217 4.5005
R80503 VDD.n1277 VDD.n1217 4.5005
R80504 VDD.n1403 VDD.n1217 4.5005
R80505 VDD.n1276 VDD.n1217 4.5005
R80506 VDD.n1404 VDD.n1217 4.5005
R80507 VDD.n1274 VDD.n1217 4.5005
R80508 VDD.n1405 VDD.n1217 4.5005
R80509 VDD.n1273 VDD.n1217 4.5005
R80510 VDD.n1406 VDD.n1217 4.5005
R80511 VDD.n1271 VDD.n1217 4.5005
R80512 VDD.n1407 VDD.n1217 4.5005
R80513 VDD.n1270 VDD.n1217 4.5005
R80514 VDD.n1408 VDD.n1217 4.5005
R80515 VDD.n1268 VDD.n1217 4.5005
R80516 VDD.n1409 VDD.n1217 4.5005
R80517 VDD.n1267 VDD.n1217 4.5005
R80518 VDD.n1410 VDD.n1217 4.5005
R80519 VDD.n1265 VDD.n1217 4.5005
R80520 VDD.n1411 VDD.n1217 4.5005
R80521 VDD.n1264 VDD.n1217 4.5005
R80522 VDD.n1412 VDD.n1217 4.5005
R80523 VDD.n1262 VDD.n1217 4.5005
R80524 VDD.n1413 VDD.n1217 4.5005
R80525 VDD.n1261 VDD.n1217 4.5005
R80526 VDD.n1414 VDD.n1217 4.5005
R80527 VDD.n1415 VDD.n1217 4.5005
R80528 VDD.n1674 VDD.n1217 4.5005
R80529 VDD.n1676 VDD.n1172 4.5005
R80530 VDD.n1341 VDD.n1172 4.5005
R80531 VDD.n1342 VDD.n1172 4.5005
R80532 VDD.n1340 VDD.n1172 4.5005
R80533 VDD.n1344 VDD.n1172 4.5005
R80534 VDD.n1339 VDD.n1172 4.5005
R80535 VDD.n1345 VDD.n1172 4.5005
R80536 VDD.n1338 VDD.n1172 4.5005
R80537 VDD.n1347 VDD.n1172 4.5005
R80538 VDD.n1337 VDD.n1172 4.5005
R80539 VDD.n1348 VDD.n1172 4.5005
R80540 VDD.n1336 VDD.n1172 4.5005
R80541 VDD.n1350 VDD.n1172 4.5005
R80542 VDD.n1335 VDD.n1172 4.5005
R80543 VDD.n1351 VDD.n1172 4.5005
R80544 VDD.n1334 VDD.n1172 4.5005
R80545 VDD.n1353 VDD.n1172 4.5005
R80546 VDD.n1333 VDD.n1172 4.5005
R80547 VDD.n1354 VDD.n1172 4.5005
R80548 VDD.n1332 VDD.n1172 4.5005
R80549 VDD.n1356 VDD.n1172 4.5005
R80550 VDD.n1331 VDD.n1172 4.5005
R80551 VDD.n1357 VDD.n1172 4.5005
R80552 VDD.n1330 VDD.n1172 4.5005
R80553 VDD.n1359 VDD.n1172 4.5005
R80554 VDD.n1329 VDD.n1172 4.5005
R80555 VDD.n1360 VDD.n1172 4.5005
R80556 VDD.n1328 VDD.n1172 4.5005
R80557 VDD.n1362 VDD.n1172 4.5005
R80558 VDD.n1327 VDD.n1172 4.5005
R80559 VDD.n1363 VDD.n1172 4.5005
R80560 VDD.n1326 VDD.n1172 4.5005
R80561 VDD.n1365 VDD.n1172 4.5005
R80562 VDD.n1325 VDD.n1172 4.5005
R80563 VDD.n1366 VDD.n1172 4.5005
R80564 VDD.n1324 VDD.n1172 4.5005
R80565 VDD.n1368 VDD.n1172 4.5005
R80566 VDD.n1323 VDD.n1172 4.5005
R80567 VDD.n1369 VDD.n1172 4.5005
R80568 VDD.n1322 VDD.n1172 4.5005
R80569 VDD.n1371 VDD.n1172 4.5005
R80570 VDD.n1321 VDD.n1172 4.5005
R80571 VDD.n1372 VDD.n1172 4.5005
R80572 VDD.n1320 VDD.n1172 4.5005
R80573 VDD.n1374 VDD.n1172 4.5005
R80574 VDD.n1319 VDD.n1172 4.5005
R80575 VDD.n1375 VDD.n1172 4.5005
R80576 VDD.n1318 VDD.n1172 4.5005
R80577 VDD.n1376 VDD.n1172 4.5005
R80578 VDD.n1316 VDD.n1172 4.5005
R80579 VDD.n1377 VDD.n1172 4.5005
R80580 VDD.n1315 VDD.n1172 4.5005
R80581 VDD.n1378 VDD.n1172 4.5005
R80582 VDD.n1313 VDD.n1172 4.5005
R80583 VDD.n1379 VDD.n1172 4.5005
R80584 VDD.n1312 VDD.n1172 4.5005
R80585 VDD.n1380 VDD.n1172 4.5005
R80586 VDD.n1310 VDD.n1172 4.5005
R80587 VDD.n1381 VDD.n1172 4.5005
R80588 VDD.n1309 VDD.n1172 4.5005
R80589 VDD.n1382 VDD.n1172 4.5005
R80590 VDD.n1307 VDD.n1172 4.5005
R80591 VDD.n1383 VDD.n1172 4.5005
R80592 VDD.n1306 VDD.n1172 4.5005
R80593 VDD.n1384 VDD.n1172 4.5005
R80594 VDD.n1304 VDD.n1172 4.5005
R80595 VDD.n1385 VDD.n1172 4.5005
R80596 VDD.n1303 VDD.n1172 4.5005
R80597 VDD.n1386 VDD.n1172 4.5005
R80598 VDD.n1301 VDD.n1172 4.5005
R80599 VDD.n1387 VDD.n1172 4.5005
R80600 VDD.n1300 VDD.n1172 4.5005
R80601 VDD.n1388 VDD.n1172 4.5005
R80602 VDD.n1298 VDD.n1172 4.5005
R80603 VDD.n1389 VDD.n1172 4.5005
R80604 VDD.n1297 VDD.n1172 4.5005
R80605 VDD.n1390 VDD.n1172 4.5005
R80606 VDD.n1295 VDD.n1172 4.5005
R80607 VDD.n1391 VDD.n1172 4.5005
R80608 VDD.n1294 VDD.n1172 4.5005
R80609 VDD.n1392 VDD.n1172 4.5005
R80610 VDD.n1292 VDD.n1172 4.5005
R80611 VDD.n1393 VDD.n1172 4.5005
R80612 VDD.n1291 VDD.n1172 4.5005
R80613 VDD.n1394 VDD.n1172 4.5005
R80614 VDD.n1289 VDD.n1172 4.5005
R80615 VDD.n1395 VDD.n1172 4.5005
R80616 VDD.n1288 VDD.n1172 4.5005
R80617 VDD.n1396 VDD.n1172 4.5005
R80618 VDD.n1286 VDD.n1172 4.5005
R80619 VDD.n1397 VDD.n1172 4.5005
R80620 VDD.n1285 VDD.n1172 4.5005
R80621 VDD.n1398 VDD.n1172 4.5005
R80622 VDD.n1283 VDD.n1172 4.5005
R80623 VDD.n1399 VDD.n1172 4.5005
R80624 VDD.n1282 VDD.n1172 4.5005
R80625 VDD.n1400 VDD.n1172 4.5005
R80626 VDD.n1280 VDD.n1172 4.5005
R80627 VDD.n1401 VDD.n1172 4.5005
R80628 VDD.n1279 VDD.n1172 4.5005
R80629 VDD.n1402 VDD.n1172 4.5005
R80630 VDD.n1277 VDD.n1172 4.5005
R80631 VDD.n1403 VDD.n1172 4.5005
R80632 VDD.n1276 VDD.n1172 4.5005
R80633 VDD.n1404 VDD.n1172 4.5005
R80634 VDD.n1274 VDD.n1172 4.5005
R80635 VDD.n1405 VDD.n1172 4.5005
R80636 VDD.n1273 VDD.n1172 4.5005
R80637 VDD.n1406 VDD.n1172 4.5005
R80638 VDD.n1271 VDD.n1172 4.5005
R80639 VDD.n1407 VDD.n1172 4.5005
R80640 VDD.n1270 VDD.n1172 4.5005
R80641 VDD.n1408 VDD.n1172 4.5005
R80642 VDD.n1268 VDD.n1172 4.5005
R80643 VDD.n1409 VDD.n1172 4.5005
R80644 VDD.n1267 VDD.n1172 4.5005
R80645 VDD.n1410 VDD.n1172 4.5005
R80646 VDD.n1265 VDD.n1172 4.5005
R80647 VDD.n1411 VDD.n1172 4.5005
R80648 VDD.n1264 VDD.n1172 4.5005
R80649 VDD.n1412 VDD.n1172 4.5005
R80650 VDD.n1262 VDD.n1172 4.5005
R80651 VDD.n1413 VDD.n1172 4.5005
R80652 VDD.n1261 VDD.n1172 4.5005
R80653 VDD.n1414 VDD.n1172 4.5005
R80654 VDD.n1415 VDD.n1172 4.5005
R80655 VDD.n1674 VDD.n1172 4.5005
R80656 VDD.n1676 VDD.n1218 4.5005
R80657 VDD.n1341 VDD.n1218 4.5005
R80658 VDD.n1342 VDD.n1218 4.5005
R80659 VDD.n1340 VDD.n1218 4.5005
R80660 VDD.n1344 VDD.n1218 4.5005
R80661 VDD.n1339 VDD.n1218 4.5005
R80662 VDD.n1345 VDD.n1218 4.5005
R80663 VDD.n1338 VDD.n1218 4.5005
R80664 VDD.n1347 VDD.n1218 4.5005
R80665 VDD.n1337 VDD.n1218 4.5005
R80666 VDD.n1348 VDD.n1218 4.5005
R80667 VDD.n1336 VDD.n1218 4.5005
R80668 VDD.n1350 VDD.n1218 4.5005
R80669 VDD.n1335 VDD.n1218 4.5005
R80670 VDD.n1351 VDD.n1218 4.5005
R80671 VDD.n1334 VDD.n1218 4.5005
R80672 VDD.n1353 VDD.n1218 4.5005
R80673 VDD.n1333 VDD.n1218 4.5005
R80674 VDD.n1354 VDD.n1218 4.5005
R80675 VDD.n1332 VDD.n1218 4.5005
R80676 VDD.n1356 VDD.n1218 4.5005
R80677 VDD.n1331 VDD.n1218 4.5005
R80678 VDD.n1357 VDD.n1218 4.5005
R80679 VDD.n1330 VDD.n1218 4.5005
R80680 VDD.n1359 VDD.n1218 4.5005
R80681 VDD.n1329 VDD.n1218 4.5005
R80682 VDD.n1360 VDD.n1218 4.5005
R80683 VDD.n1328 VDD.n1218 4.5005
R80684 VDD.n1362 VDD.n1218 4.5005
R80685 VDD.n1327 VDD.n1218 4.5005
R80686 VDD.n1363 VDD.n1218 4.5005
R80687 VDD.n1326 VDD.n1218 4.5005
R80688 VDD.n1365 VDD.n1218 4.5005
R80689 VDD.n1325 VDD.n1218 4.5005
R80690 VDD.n1366 VDD.n1218 4.5005
R80691 VDD.n1324 VDD.n1218 4.5005
R80692 VDD.n1368 VDD.n1218 4.5005
R80693 VDD.n1323 VDD.n1218 4.5005
R80694 VDD.n1369 VDD.n1218 4.5005
R80695 VDD.n1322 VDD.n1218 4.5005
R80696 VDD.n1371 VDD.n1218 4.5005
R80697 VDD.n1321 VDD.n1218 4.5005
R80698 VDD.n1372 VDD.n1218 4.5005
R80699 VDD.n1320 VDD.n1218 4.5005
R80700 VDD.n1374 VDD.n1218 4.5005
R80701 VDD.n1319 VDD.n1218 4.5005
R80702 VDD.n1375 VDD.n1218 4.5005
R80703 VDD.n1318 VDD.n1218 4.5005
R80704 VDD.n1376 VDD.n1218 4.5005
R80705 VDD.n1316 VDD.n1218 4.5005
R80706 VDD.n1377 VDD.n1218 4.5005
R80707 VDD.n1315 VDD.n1218 4.5005
R80708 VDD.n1378 VDD.n1218 4.5005
R80709 VDD.n1313 VDD.n1218 4.5005
R80710 VDD.n1379 VDD.n1218 4.5005
R80711 VDD.n1312 VDD.n1218 4.5005
R80712 VDD.n1380 VDD.n1218 4.5005
R80713 VDD.n1310 VDD.n1218 4.5005
R80714 VDD.n1381 VDD.n1218 4.5005
R80715 VDD.n1309 VDD.n1218 4.5005
R80716 VDD.n1382 VDD.n1218 4.5005
R80717 VDD.n1307 VDD.n1218 4.5005
R80718 VDD.n1383 VDD.n1218 4.5005
R80719 VDD.n1306 VDD.n1218 4.5005
R80720 VDD.n1384 VDD.n1218 4.5005
R80721 VDD.n1304 VDD.n1218 4.5005
R80722 VDD.n1385 VDD.n1218 4.5005
R80723 VDD.n1303 VDD.n1218 4.5005
R80724 VDD.n1386 VDD.n1218 4.5005
R80725 VDD.n1301 VDD.n1218 4.5005
R80726 VDD.n1387 VDD.n1218 4.5005
R80727 VDD.n1300 VDD.n1218 4.5005
R80728 VDD.n1388 VDD.n1218 4.5005
R80729 VDD.n1298 VDD.n1218 4.5005
R80730 VDD.n1389 VDD.n1218 4.5005
R80731 VDD.n1297 VDD.n1218 4.5005
R80732 VDD.n1390 VDD.n1218 4.5005
R80733 VDD.n1295 VDD.n1218 4.5005
R80734 VDD.n1391 VDD.n1218 4.5005
R80735 VDD.n1294 VDD.n1218 4.5005
R80736 VDD.n1392 VDD.n1218 4.5005
R80737 VDD.n1292 VDD.n1218 4.5005
R80738 VDD.n1393 VDD.n1218 4.5005
R80739 VDD.n1291 VDD.n1218 4.5005
R80740 VDD.n1394 VDD.n1218 4.5005
R80741 VDD.n1289 VDD.n1218 4.5005
R80742 VDD.n1395 VDD.n1218 4.5005
R80743 VDD.n1288 VDD.n1218 4.5005
R80744 VDD.n1396 VDD.n1218 4.5005
R80745 VDD.n1286 VDD.n1218 4.5005
R80746 VDD.n1397 VDD.n1218 4.5005
R80747 VDD.n1285 VDD.n1218 4.5005
R80748 VDD.n1398 VDD.n1218 4.5005
R80749 VDD.n1283 VDD.n1218 4.5005
R80750 VDD.n1399 VDD.n1218 4.5005
R80751 VDD.n1282 VDD.n1218 4.5005
R80752 VDD.n1400 VDD.n1218 4.5005
R80753 VDD.n1280 VDD.n1218 4.5005
R80754 VDD.n1401 VDD.n1218 4.5005
R80755 VDD.n1279 VDD.n1218 4.5005
R80756 VDD.n1402 VDD.n1218 4.5005
R80757 VDD.n1277 VDD.n1218 4.5005
R80758 VDD.n1403 VDD.n1218 4.5005
R80759 VDD.n1276 VDD.n1218 4.5005
R80760 VDD.n1404 VDD.n1218 4.5005
R80761 VDD.n1274 VDD.n1218 4.5005
R80762 VDD.n1405 VDD.n1218 4.5005
R80763 VDD.n1273 VDD.n1218 4.5005
R80764 VDD.n1406 VDD.n1218 4.5005
R80765 VDD.n1271 VDD.n1218 4.5005
R80766 VDD.n1407 VDD.n1218 4.5005
R80767 VDD.n1270 VDD.n1218 4.5005
R80768 VDD.n1408 VDD.n1218 4.5005
R80769 VDD.n1268 VDD.n1218 4.5005
R80770 VDD.n1409 VDD.n1218 4.5005
R80771 VDD.n1267 VDD.n1218 4.5005
R80772 VDD.n1410 VDD.n1218 4.5005
R80773 VDD.n1265 VDD.n1218 4.5005
R80774 VDD.n1411 VDD.n1218 4.5005
R80775 VDD.n1264 VDD.n1218 4.5005
R80776 VDD.n1412 VDD.n1218 4.5005
R80777 VDD.n1262 VDD.n1218 4.5005
R80778 VDD.n1413 VDD.n1218 4.5005
R80779 VDD.n1261 VDD.n1218 4.5005
R80780 VDD.n1414 VDD.n1218 4.5005
R80781 VDD.n1415 VDD.n1218 4.5005
R80782 VDD.n1674 VDD.n1218 4.5005
R80783 VDD.n1676 VDD.n1171 4.5005
R80784 VDD.n1341 VDD.n1171 4.5005
R80785 VDD.n1342 VDD.n1171 4.5005
R80786 VDD.n1340 VDD.n1171 4.5005
R80787 VDD.n1344 VDD.n1171 4.5005
R80788 VDD.n1339 VDD.n1171 4.5005
R80789 VDD.n1345 VDD.n1171 4.5005
R80790 VDD.n1338 VDD.n1171 4.5005
R80791 VDD.n1347 VDD.n1171 4.5005
R80792 VDD.n1337 VDD.n1171 4.5005
R80793 VDD.n1348 VDD.n1171 4.5005
R80794 VDD.n1336 VDD.n1171 4.5005
R80795 VDD.n1350 VDD.n1171 4.5005
R80796 VDD.n1335 VDD.n1171 4.5005
R80797 VDD.n1351 VDD.n1171 4.5005
R80798 VDD.n1334 VDD.n1171 4.5005
R80799 VDD.n1353 VDD.n1171 4.5005
R80800 VDD.n1333 VDD.n1171 4.5005
R80801 VDD.n1354 VDD.n1171 4.5005
R80802 VDD.n1332 VDD.n1171 4.5005
R80803 VDD.n1356 VDD.n1171 4.5005
R80804 VDD.n1331 VDD.n1171 4.5005
R80805 VDD.n1357 VDD.n1171 4.5005
R80806 VDD.n1330 VDD.n1171 4.5005
R80807 VDD.n1359 VDD.n1171 4.5005
R80808 VDD.n1329 VDD.n1171 4.5005
R80809 VDD.n1360 VDD.n1171 4.5005
R80810 VDD.n1328 VDD.n1171 4.5005
R80811 VDD.n1362 VDD.n1171 4.5005
R80812 VDD.n1327 VDD.n1171 4.5005
R80813 VDD.n1363 VDD.n1171 4.5005
R80814 VDD.n1326 VDD.n1171 4.5005
R80815 VDD.n1365 VDD.n1171 4.5005
R80816 VDD.n1325 VDD.n1171 4.5005
R80817 VDD.n1366 VDD.n1171 4.5005
R80818 VDD.n1324 VDD.n1171 4.5005
R80819 VDD.n1368 VDD.n1171 4.5005
R80820 VDD.n1323 VDD.n1171 4.5005
R80821 VDD.n1369 VDD.n1171 4.5005
R80822 VDD.n1322 VDD.n1171 4.5005
R80823 VDD.n1371 VDD.n1171 4.5005
R80824 VDD.n1321 VDD.n1171 4.5005
R80825 VDD.n1372 VDD.n1171 4.5005
R80826 VDD.n1320 VDD.n1171 4.5005
R80827 VDD.n1374 VDD.n1171 4.5005
R80828 VDD.n1319 VDD.n1171 4.5005
R80829 VDD.n1375 VDD.n1171 4.5005
R80830 VDD.n1318 VDD.n1171 4.5005
R80831 VDD.n1376 VDD.n1171 4.5005
R80832 VDD.n1316 VDD.n1171 4.5005
R80833 VDD.n1377 VDD.n1171 4.5005
R80834 VDD.n1315 VDD.n1171 4.5005
R80835 VDD.n1378 VDD.n1171 4.5005
R80836 VDD.n1313 VDD.n1171 4.5005
R80837 VDD.n1379 VDD.n1171 4.5005
R80838 VDD.n1312 VDD.n1171 4.5005
R80839 VDD.n1380 VDD.n1171 4.5005
R80840 VDD.n1310 VDD.n1171 4.5005
R80841 VDD.n1381 VDD.n1171 4.5005
R80842 VDD.n1309 VDD.n1171 4.5005
R80843 VDD.n1382 VDD.n1171 4.5005
R80844 VDD.n1307 VDD.n1171 4.5005
R80845 VDD.n1383 VDD.n1171 4.5005
R80846 VDD.n1306 VDD.n1171 4.5005
R80847 VDD.n1384 VDD.n1171 4.5005
R80848 VDD.n1304 VDD.n1171 4.5005
R80849 VDD.n1385 VDD.n1171 4.5005
R80850 VDD.n1303 VDD.n1171 4.5005
R80851 VDD.n1386 VDD.n1171 4.5005
R80852 VDD.n1301 VDD.n1171 4.5005
R80853 VDD.n1387 VDD.n1171 4.5005
R80854 VDD.n1300 VDD.n1171 4.5005
R80855 VDD.n1388 VDD.n1171 4.5005
R80856 VDD.n1298 VDD.n1171 4.5005
R80857 VDD.n1389 VDD.n1171 4.5005
R80858 VDD.n1297 VDD.n1171 4.5005
R80859 VDD.n1390 VDD.n1171 4.5005
R80860 VDD.n1295 VDD.n1171 4.5005
R80861 VDD.n1391 VDD.n1171 4.5005
R80862 VDD.n1294 VDD.n1171 4.5005
R80863 VDD.n1392 VDD.n1171 4.5005
R80864 VDD.n1292 VDD.n1171 4.5005
R80865 VDD.n1393 VDD.n1171 4.5005
R80866 VDD.n1291 VDD.n1171 4.5005
R80867 VDD.n1394 VDD.n1171 4.5005
R80868 VDD.n1289 VDD.n1171 4.5005
R80869 VDD.n1395 VDD.n1171 4.5005
R80870 VDD.n1288 VDD.n1171 4.5005
R80871 VDD.n1396 VDD.n1171 4.5005
R80872 VDD.n1286 VDD.n1171 4.5005
R80873 VDD.n1397 VDD.n1171 4.5005
R80874 VDD.n1285 VDD.n1171 4.5005
R80875 VDD.n1398 VDD.n1171 4.5005
R80876 VDD.n1283 VDD.n1171 4.5005
R80877 VDD.n1399 VDD.n1171 4.5005
R80878 VDD.n1282 VDD.n1171 4.5005
R80879 VDD.n1400 VDD.n1171 4.5005
R80880 VDD.n1280 VDD.n1171 4.5005
R80881 VDD.n1401 VDD.n1171 4.5005
R80882 VDD.n1279 VDD.n1171 4.5005
R80883 VDD.n1402 VDD.n1171 4.5005
R80884 VDD.n1277 VDD.n1171 4.5005
R80885 VDD.n1403 VDD.n1171 4.5005
R80886 VDD.n1276 VDD.n1171 4.5005
R80887 VDD.n1404 VDD.n1171 4.5005
R80888 VDD.n1274 VDD.n1171 4.5005
R80889 VDD.n1405 VDD.n1171 4.5005
R80890 VDD.n1273 VDD.n1171 4.5005
R80891 VDD.n1406 VDD.n1171 4.5005
R80892 VDD.n1271 VDD.n1171 4.5005
R80893 VDD.n1407 VDD.n1171 4.5005
R80894 VDD.n1270 VDD.n1171 4.5005
R80895 VDD.n1408 VDD.n1171 4.5005
R80896 VDD.n1268 VDD.n1171 4.5005
R80897 VDD.n1409 VDD.n1171 4.5005
R80898 VDD.n1267 VDD.n1171 4.5005
R80899 VDD.n1410 VDD.n1171 4.5005
R80900 VDD.n1265 VDD.n1171 4.5005
R80901 VDD.n1411 VDD.n1171 4.5005
R80902 VDD.n1264 VDD.n1171 4.5005
R80903 VDD.n1412 VDD.n1171 4.5005
R80904 VDD.n1262 VDD.n1171 4.5005
R80905 VDD.n1413 VDD.n1171 4.5005
R80906 VDD.n1261 VDD.n1171 4.5005
R80907 VDD.n1414 VDD.n1171 4.5005
R80908 VDD.n1415 VDD.n1171 4.5005
R80909 VDD.n1674 VDD.n1171 4.5005
R80910 VDD.n1676 VDD.n1219 4.5005
R80911 VDD.n1341 VDD.n1219 4.5005
R80912 VDD.n1342 VDD.n1219 4.5005
R80913 VDD.n1340 VDD.n1219 4.5005
R80914 VDD.n1344 VDD.n1219 4.5005
R80915 VDD.n1339 VDD.n1219 4.5005
R80916 VDD.n1345 VDD.n1219 4.5005
R80917 VDD.n1338 VDD.n1219 4.5005
R80918 VDD.n1347 VDD.n1219 4.5005
R80919 VDD.n1337 VDD.n1219 4.5005
R80920 VDD.n1348 VDD.n1219 4.5005
R80921 VDD.n1336 VDD.n1219 4.5005
R80922 VDD.n1350 VDD.n1219 4.5005
R80923 VDD.n1335 VDD.n1219 4.5005
R80924 VDD.n1351 VDD.n1219 4.5005
R80925 VDD.n1334 VDD.n1219 4.5005
R80926 VDD.n1353 VDD.n1219 4.5005
R80927 VDD.n1333 VDD.n1219 4.5005
R80928 VDD.n1354 VDD.n1219 4.5005
R80929 VDD.n1332 VDD.n1219 4.5005
R80930 VDD.n1356 VDD.n1219 4.5005
R80931 VDD.n1331 VDD.n1219 4.5005
R80932 VDD.n1357 VDD.n1219 4.5005
R80933 VDD.n1330 VDD.n1219 4.5005
R80934 VDD.n1359 VDD.n1219 4.5005
R80935 VDD.n1329 VDD.n1219 4.5005
R80936 VDD.n1360 VDD.n1219 4.5005
R80937 VDD.n1328 VDD.n1219 4.5005
R80938 VDD.n1362 VDD.n1219 4.5005
R80939 VDD.n1327 VDD.n1219 4.5005
R80940 VDD.n1363 VDD.n1219 4.5005
R80941 VDD.n1326 VDD.n1219 4.5005
R80942 VDD.n1365 VDD.n1219 4.5005
R80943 VDD.n1325 VDD.n1219 4.5005
R80944 VDD.n1366 VDD.n1219 4.5005
R80945 VDD.n1324 VDD.n1219 4.5005
R80946 VDD.n1368 VDD.n1219 4.5005
R80947 VDD.n1323 VDD.n1219 4.5005
R80948 VDD.n1369 VDD.n1219 4.5005
R80949 VDD.n1322 VDD.n1219 4.5005
R80950 VDD.n1371 VDD.n1219 4.5005
R80951 VDD.n1321 VDD.n1219 4.5005
R80952 VDD.n1372 VDD.n1219 4.5005
R80953 VDD.n1320 VDD.n1219 4.5005
R80954 VDD.n1374 VDD.n1219 4.5005
R80955 VDD.n1319 VDD.n1219 4.5005
R80956 VDD.n1375 VDD.n1219 4.5005
R80957 VDD.n1318 VDD.n1219 4.5005
R80958 VDD.n1376 VDD.n1219 4.5005
R80959 VDD.n1316 VDD.n1219 4.5005
R80960 VDD.n1377 VDD.n1219 4.5005
R80961 VDD.n1315 VDD.n1219 4.5005
R80962 VDD.n1378 VDD.n1219 4.5005
R80963 VDD.n1313 VDD.n1219 4.5005
R80964 VDD.n1379 VDD.n1219 4.5005
R80965 VDD.n1312 VDD.n1219 4.5005
R80966 VDD.n1380 VDD.n1219 4.5005
R80967 VDD.n1310 VDD.n1219 4.5005
R80968 VDD.n1381 VDD.n1219 4.5005
R80969 VDD.n1309 VDD.n1219 4.5005
R80970 VDD.n1382 VDD.n1219 4.5005
R80971 VDD.n1307 VDD.n1219 4.5005
R80972 VDD.n1383 VDD.n1219 4.5005
R80973 VDD.n1306 VDD.n1219 4.5005
R80974 VDD.n1384 VDD.n1219 4.5005
R80975 VDD.n1304 VDD.n1219 4.5005
R80976 VDD.n1385 VDD.n1219 4.5005
R80977 VDD.n1303 VDD.n1219 4.5005
R80978 VDD.n1386 VDD.n1219 4.5005
R80979 VDD.n1301 VDD.n1219 4.5005
R80980 VDD.n1387 VDD.n1219 4.5005
R80981 VDD.n1300 VDD.n1219 4.5005
R80982 VDD.n1388 VDD.n1219 4.5005
R80983 VDD.n1298 VDD.n1219 4.5005
R80984 VDD.n1389 VDD.n1219 4.5005
R80985 VDD.n1297 VDD.n1219 4.5005
R80986 VDD.n1390 VDD.n1219 4.5005
R80987 VDD.n1295 VDD.n1219 4.5005
R80988 VDD.n1391 VDD.n1219 4.5005
R80989 VDD.n1294 VDD.n1219 4.5005
R80990 VDD.n1392 VDD.n1219 4.5005
R80991 VDD.n1292 VDD.n1219 4.5005
R80992 VDD.n1393 VDD.n1219 4.5005
R80993 VDD.n1291 VDD.n1219 4.5005
R80994 VDD.n1394 VDD.n1219 4.5005
R80995 VDD.n1289 VDD.n1219 4.5005
R80996 VDD.n1395 VDD.n1219 4.5005
R80997 VDD.n1288 VDD.n1219 4.5005
R80998 VDD.n1396 VDD.n1219 4.5005
R80999 VDD.n1286 VDD.n1219 4.5005
R81000 VDD.n1397 VDD.n1219 4.5005
R81001 VDD.n1285 VDD.n1219 4.5005
R81002 VDD.n1398 VDD.n1219 4.5005
R81003 VDD.n1283 VDD.n1219 4.5005
R81004 VDD.n1399 VDD.n1219 4.5005
R81005 VDD.n1282 VDD.n1219 4.5005
R81006 VDD.n1400 VDD.n1219 4.5005
R81007 VDD.n1280 VDD.n1219 4.5005
R81008 VDD.n1401 VDD.n1219 4.5005
R81009 VDD.n1279 VDD.n1219 4.5005
R81010 VDD.n1402 VDD.n1219 4.5005
R81011 VDD.n1277 VDD.n1219 4.5005
R81012 VDD.n1403 VDD.n1219 4.5005
R81013 VDD.n1276 VDD.n1219 4.5005
R81014 VDD.n1404 VDD.n1219 4.5005
R81015 VDD.n1274 VDD.n1219 4.5005
R81016 VDD.n1405 VDD.n1219 4.5005
R81017 VDD.n1273 VDD.n1219 4.5005
R81018 VDD.n1406 VDD.n1219 4.5005
R81019 VDD.n1271 VDD.n1219 4.5005
R81020 VDD.n1407 VDD.n1219 4.5005
R81021 VDD.n1270 VDD.n1219 4.5005
R81022 VDD.n1408 VDD.n1219 4.5005
R81023 VDD.n1268 VDD.n1219 4.5005
R81024 VDD.n1409 VDD.n1219 4.5005
R81025 VDD.n1267 VDD.n1219 4.5005
R81026 VDD.n1410 VDD.n1219 4.5005
R81027 VDD.n1265 VDD.n1219 4.5005
R81028 VDD.n1411 VDD.n1219 4.5005
R81029 VDD.n1264 VDD.n1219 4.5005
R81030 VDD.n1412 VDD.n1219 4.5005
R81031 VDD.n1262 VDD.n1219 4.5005
R81032 VDD.n1413 VDD.n1219 4.5005
R81033 VDD.n1261 VDD.n1219 4.5005
R81034 VDD.n1414 VDD.n1219 4.5005
R81035 VDD.n1415 VDD.n1219 4.5005
R81036 VDD.n1674 VDD.n1219 4.5005
R81037 VDD.n1676 VDD.n1170 4.5005
R81038 VDD.n1341 VDD.n1170 4.5005
R81039 VDD.n1342 VDD.n1170 4.5005
R81040 VDD.n1340 VDD.n1170 4.5005
R81041 VDD.n1344 VDD.n1170 4.5005
R81042 VDD.n1339 VDD.n1170 4.5005
R81043 VDD.n1345 VDD.n1170 4.5005
R81044 VDD.n1338 VDD.n1170 4.5005
R81045 VDD.n1347 VDD.n1170 4.5005
R81046 VDD.n1337 VDD.n1170 4.5005
R81047 VDD.n1348 VDD.n1170 4.5005
R81048 VDD.n1336 VDD.n1170 4.5005
R81049 VDD.n1350 VDD.n1170 4.5005
R81050 VDD.n1335 VDD.n1170 4.5005
R81051 VDD.n1351 VDD.n1170 4.5005
R81052 VDD.n1334 VDD.n1170 4.5005
R81053 VDD.n1353 VDD.n1170 4.5005
R81054 VDD.n1333 VDD.n1170 4.5005
R81055 VDD.n1354 VDD.n1170 4.5005
R81056 VDD.n1332 VDD.n1170 4.5005
R81057 VDD.n1356 VDD.n1170 4.5005
R81058 VDD.n1331 VDD.n1170 4.5005
R81059 VDD.n1357 VDD.n1170 4.5005
R81060 VDD.n1330 VDD.n1170 4.5005
R81061 VDD.n1359 VDD.n1170 4.5005
R81062 VDD.n1329 VDD.n1170 4.5005
R81063 VDD.n1360 VDD.n1170 4.5005
R81064 VDD.n1328 VDD.n1170 4.5005
R81065 VDD.n1362 VDD.n1170 4.5005
R81066 VDD.n1327 VDD.n1170 4.5005
R81067 VDD.n1363 VDD.n1170 4.5005
R81068 VDD.n1326 VDD.n1170 4.5005
R81069 VDD.n1365 VDD.n1170 4.5005
R81070 VDD.n1325 VDD.n1170 4.5005
R81071 VDD.n1366 VDD.n1170 4.5005
R81072 VDD.n1324 VDD.n1170 4.5005
R81073 VDD.n1368 VDD.n1170 4.5005
R81074 VDD.n1323 VDD.n1170 4.5005
R81075 VDD.n1369 VDD.n1170 4.5005
R81076 VDD.n1322 VDD.n1170 4.5005
R81077 VDD.n1371 VDD.n1170 4.5005
R81078 VDD.n1321 VDD.n1170 4.5005
R81079 VDD.n1372 VDD.n1170 4.5005
R81080 VDD.n1320 VDD.n1170 4.5005
R81081 VDD.n1374 VDD.n1170 4.5005
R81082 VDD.n1319 VDD.n1170 4.5005
R81083 VDD.n1375 VDD.n1170 4.5005
R81084 VDD.n1318 VDD.n1170 4.5005
R81085 VDD.n1376 VDD.n1170 4.5005
R81086 VDD.n1316 VDD.n1170 4.5005
R81087 VDD.n1377 VDD.n1170 4.5005
R81088 VDD.n1315 VDD.n1170 4.5005
R81089 VDD.n1378 VDD.n1170 4.5005
R81090 VDD.n1313 VDD.n1170 4.5005
R81091 VDD.n1379 VDD.n1170 4.5005
R81092 VDD.n1312 VDD.n1170 4.5005
R81093 VDD.n1380 VDD.n1170 4.5005
R81094 VDD.n1310 VDD.n1170 4.5005
R81095 VDD.n1381 VDD.n1170 4.5005
R81096 VDD.n1309 VDD.n1170 4.5005
R81097 VDD.n1382 VDD.n1170 4.5005
R81098 VDD.n1307 VDD.n1170 4.5005
R81099 VDD.n1383 VDD.n1170 4.5005
R81100 VDD.n1306 VDD.n1170 4.5005
R81101 VDD.n1384 VDD.n1170 4.5005
R81102 VDD.n1304 VDD.n1170 4.5005
R81103 VDD.n1385 VDD.n1170 4.5005
R81104 VDD.n1303 VDD.n1170 4.5005
R81105 VDD.n1386 VDD.n1170 4.5005
R81106 VDD.n1301 VDD.n1170 4.5005
R81107 VDD.n1387 VDD.n1170 4.5005
R81108 VDD.n1300 VDD.n1170 4.5005
R81109 VDD.n1388 VDD.n1170 4.5005
R81110 VDD.n1298 VDD.n1170 4.5005
R81111 VDD.n1389 VDD.n1170 4.5005
R81112 VDD.n1297 VDD.n1170 4.5005
R81113 VDD.n1390 VDD.n1170 4.5005
R81114 VDD.n1295 VDD.n1170 4.5005
R81115 VDD.n1391 VDD.n1170 4.5005
R81116 VDD.n1294 VDD.n1170 4.5005
R81117 VDD.n1392 VDD.n1170 4.5005
R81118 VDD.n1292 VDD.n1170 4.5005
R81119 VDD.n1393 VDD.n1170 4.5005
R81120 VDD.n1291 VDD.n1170 4.5005
R81121 VDD.n1394 VDD.n1170 4.5005
R81122 VDD.n1289 VDD.n1170 4.5005
R81123 VDD.n1395 VDD.n1170 4.5005
R81124 VDD.n1288 VDD.n1170 4.5005
R81125 VDD.n1396 VDD.n1170 4.5005
R81126 VDD.n1286 VDD.n1170 4.5005
R81127 VDD.n1397 VDD.n1170 4.5005
R81128 VDD.n1285 VDD.n1170 4.5005
R81129 VDD.n1398 VDD.n1170 4.5005
R81130 VDD.n1283 VDD.n1170 4.5005
R81131 VDD.n1399 VDD.n1170 4.5005
R81132 VDD.n1282 VDD.n1170 4.5005
R81133 VDD.n1400 VDD.n1170 4.5005
R81134 VDD.n1280 VDD.n1170 4.5005
R81135 VDD.n1401 VDD.n1170 4.5005
R81136 VDD.n1279 VDD.n1170 4.5005
R81137 VDD.n1402 VDD.n1170 4.5005
R81138 VDD.n1277 VDD.n1170 4.5005
R81139 VDD.n1403 VDD.n1170 4.5005
R81140 VDD.n1276 VDD.n1170 4.5005
R81141 VDD.n1404 VDD.n1170 4.5005
R81142 VDD.n1274 VDD.n1170 4.5005
R81143 VDD.n1405 VDD.n1170 4.5005
R81144 VDD.n1273 VDD.n1170 4.5005
R81145 VDD.n1406 VDD.n1170 4.5005
R81146 VDD.n1271 VDD.n1170 4.5005
R81147 VDD.n1407 VDD.n1170 4.5005
R81148 VDD.n1270 VDD.n1170 4.5005
R81149 VDD.n1408 VDD.n1170 4.5005
R81150 VDD.n1268 VDD.n1170 4.5005
R81151 VDD.n1409 VDD.n1170 4.5005
R81152 VDD.n1267 VDD.n1170 4.5005
R81153 VDD.n1410 VDD.n1170 4.5005
R81154 VDD.n1265 VDD.n1170 4.5005
R81155 VDD.n1411 VDD.n1170 4.5005
R81156 VDD.n1264 VDD.n1170 4.5005
R81157 VDD.n1412 VDD.n1170 4.5005
R81158 VDD.n1262 VDD.n1170 4.5005
R81159 VDD.n1413 VDD.n1170 4.5005
R81160 VDD.n1261 VDD.n1170 4.5005
R81161 VDD.n1414 VDD.n1170 4.5005
R81162 VDD.n1415 VDD.n1170 4.5005
R81163 VDD.n1674 VDD.n1170 4.5005
R81164 VDD.n1676 VDD.n1220 4.5005
R81165 VDD.n1341 VDD.n1220 4.5005
R81166 VDD.n1342 VDD.n1220 4.5005
R81167 VDD.n1340 VDD.n1220 4.5005
R81168 VDD.n1344 VDD.n1220 4.5005
R81169 VDD.n1339 VDD.n1220 4.5005
R81170 VDD.n1345 VDD.n1220 4.5005
R81171 VDD.n1338 VDD.n1220 4.5005
R81172 VDD.n1347 VDD.n1220 4.5005
R81173 VDD.n1337 VDD.n1220 4.5005
R81174 VDD.n1348 VDD.n1220 4.5005
R81175 VDD.n1336 VDD.n1220 4.5005
R81176 VDD.n1350 VDD.n1220 4.5005
R81177 VDD.n1335 VDD.n1220 4.5005
R81178 VDD.n1351 VDD.n1220 4.5005
R81179 VDD.n1334 VDD.n1220 4.5005
R81180 VDD.n1353 VDD.n1220 4.5005
R81181 VDD.n1333 VDD.n1220 4.5005
R81182 VDD.n1354 VDD.n1220 4.5005
R81183 VDD.n1332 VDD.n1220 4.5005
R81184 VDD.n1356 VDD.n1220 4.5005
R81185 VDD.n1331 VDD.n1220 4.5005
R81186 VDD.n1357 VDD.n1220 4.5005
R81187 VDD.n1330 VDD.n1220 4.5005
R81188 VDD.n1359 VDD.n1220 4.5005
R81189 VDD.n1329 VDD.n1220 4.5005
R81190 VDD.n1360 VDD.n1220 4.5005
R81191 VDD.n1328 VDD.n1220 4.5005
R81192 VDD.n1362 VDD.n1220 4.5005
R81193 VDD.n1327 VDD.n1220 4.5005
R81194 VDD.n1363 VDD.n1220 4.5005
R81195 VDD.n1326 VDD.n1220 4.5005
R81196 VDD.n1365 VDD.n1220 4.5005
R81197 VDD.n1325 VDD.n1220 4.5005
R81198 VDD.n1366 VDD.n1220 4.5005
R81199 VDD.n1324 VDD.n1220 4.5005
R81200 VDD.n1368 VDD.n1220 4.5005
R81201 VDD.n1323 VDD.n1220 4.5005
R81202 VDD.n1369 VDD.n1220 4.5005
R81203 VDD.n1322 VDD.n1220 4.5005
R81204 VDD.n1371 VDD.n1220 4.5005
R81205 VDD.n1321 VDD.n1220 4.5005
R81206 VDD.n1372 VDD.n1220 4.5005
R81207 VDD.n1320 VDD.n1220 4.5005
R81208 VDD.n1374 VDD.n1220 4.5005
R81209 VDD.n1319 VDD.n1220 4.5005
R81210 VDD.n1375 VDD.n1220 4.5005
R81211 VDD.n1318 VDD.n1220 4.5005
R81212 VDD.n1376 VDD.n1220 4.5005
R81213 VDD.n1316 VDD.n1220 4.5005
R81214 VDD.n1377 VDD.n1220 4.5005
R81215 VDD.n1315 VDD.n1220 4.5005
R81216 VDD.n1378 VDD.n1220 4.5005
R81217 VDD.n1313 VDD.n1220 4.5005
R81218 VDD.n1379 VDD.n1220 4.5005
R81219 VDD.n1312 VDD.n1220 4.5005
R81220 VDD.n1380 VDD.n1220 4.5005
R81221 VDD.n1310 VDD.n1220 4.5005
R81222 VDD.n1381 VDD.n1220 4.5005
R81223 VDD.n1309 VDD.n1220 4.5005
R81224 VDD.n1382 VDD.n1220 4.5005
R81225 VDD.n1307 VDD.n1220 4.5005
R81226 VDD.n1383 VDD.n1220 4.5005
R81227 VDD.n1306 VDD.n1220 4.5005
R81228 VDD.n1384 VDD.n1220 4.5005
R81229 VDD.n1304 VDD.n1220 4.5005
R81230 VDD.n1385 VDD.n1220 4.5005
R81231 VDD.n1303 VDD.n1220 4.5005
R81232 VDD.n1386 VDD.n1220 4.5005
R81233 VDD.n1301 VDD.n1220 4.5005
R81234 VDD.n1387 VDD.n1220 4.5005
R81235 VDD.n1300 VDD.n1220 4.5005
R81236 VDD.n1388 VDD.n1220 4.5005
R81237 VDD.n1298 VDD.n1220 4.5005
R81238 VDD.n1389 VDD.n1220 4.5005
R81239 VDD.n1297 VDD.n1220 4.5005
R81240 VDD.n1390 VDD.n1220 4.5005
R81241 VDD.n1295 VDD.n1220 4.5005
R81242 VDD.n1391 VDD.n1220 4.5005
R81243 VDD.n1294 VDD.n1220 4.5005
R81244 VDD.n1392 VDD.n1220 4.5005
R81245 VDD.n1292 VDD.n1220 4.5005
R81246 VDD.n1393 VDD.n1220 4.5005
R81247 VDD.n1291 VDD.n1220 4.5005
R81248 VDD.n1394 VDD.n1220 4.5005
R81249 VDD.n1289 VDD.n1220 4.5005
R81250 VDD.n1395 VDD.n1220 4.5005
R81251 VDD.n1288 VDD.n1220 4.5005
R81252 VDD.n1396 VDD.n1220 4.5005
R81253 VDD.n1286 VDD.n1220 4.5005
R81254 VDD.n1397 VDD.n1220 4.5005
R81255 VDD.n1285 VDD.n1220 4.5005
R81256 VDD.n1398 VDD.n1220 4.5005
R81257 VDD.n1283 VDD.n1220 4.5005
R81258 VDD.n1399 VDD.n1220 4.5005
R81259 VDD.n1282 VDD.n1220 4.5005
R81260 VDD.n1400 VDD.n1220 4.5005
R81261 VDD.n1280 VDD.n1220 4.5005
R81262 VDD.n1401 VDD.n1220 4.5005
R81263 VDD.n1279 VDD.n1220 4.5005
R81264 VDD.n1402 VDD.n1220 4.5005
R81265 VDD.n1277 VDD.n1220 4.5005
R81266 VDD.n1403 VDD.n1220 4.5005
R81267 VDD.n1276 VDD.n1220 4.5005
R81268 VDD.n1404 VDD.n1220 4.5005
R81269 VDD.n1274 VDD.n1220 4.5005
R81270 VDD.n1405 VDD.n1220 4.5005
R81271 VDD.n1273 VDD.n1220 4.5005
R81272 VDD.n1406 VDD.n1220 4.5005
R81273 VDD.n1271 VDD.n1220 4.5005
R81274 VDD.n1407 VDD.n1220 4.5005
R81275 VDD.n1270 VDD.n1220 4.5005
R81276 VDD.n1408 VDD.n1220 4.5005
R81277 VDD.n1268 VDD.n1220 4.5005
R81278 VDD.n1409 VDD.n1220 4.5005
R81279 VDD.n1267 VDD.n1220 4.5005
R81280 VDD.n1410 VDD.n1220 4.5005
R81281 VDD.n1265 VDD.n1220 4.5005
R81282 VDD.n1411 VDD.n1220 4.5005
R81283 VDD.n1264 VDD.n1220 4.5005
R81284 VDD.n1412 VDD.n1220 4.5005
R81285 VDD.n1262 VDD.n1220 4.5005
R81286 VDD.n1413 VDD.n1220 4.5005
R81287 VDD.n1261 VDD.n1220 4.5005
R81288 VDD.n1414 VDD.n1220 4.5005
R81289 VDD.n1415 VDD.n1220 4.5005
R81290 VDD.n1674 VDD.n1220 4.5005
R81291 VDD.n1676 VDD.n1169 4.5005
R81292 VDD.n1341 VDD.n1169 4.5005
R81293 VDD.n1342 VDD.n1169 4.5005
R81294 VDD.n1340 VDD.n1169 4.5005
R81295 VDD.n1344 VDD.n1169 4.5005
R81296 VDD.n1339 VDD.n1169 4.5005
R81297 VDD.n1345 VDD.n1169 4.5005
R81298 VDD.n1338 VDD.n1169 4.5005
R81299 VDD.n1347 VDD.n1169 4.5005
R81300 VDD.n1337 VDD.n1169 4.5005
R81301 VDD.n1348 VDD.n1169 4.5005
R81302 VDD.n1336 VDD.n1169 4.5005
R81303 VDD.n1350 VDD.n1169 4.5005
R81304 VDD.n1335 VDD.n1169 4.5005
R81305 VDD.n1351 VDD.n1169 4.5005
R81306 VDD.n1334 VDD.n1169 4.5005
R81307 VDD.n1353 VDD.n1169 4.5005
R81308 VDD.n1333 VDD.n1169 4.5005
R81309 VDD.n1354 VDD.n1169 4.5005
R81310 VDD.n1332 VDD.n1169 4.5005
R81311 VDD.n1356 VDD.n1169 4.5005
R81312 VDD.n1331 VDD.n1169 4.5005
R81313 VDD.n1357 VDD.n1169 4.5005
R81314 VDD.n1330 VDD.n1169 4.5005
R81315 VDD.n1359 VDD.n1169 4.5005
R81316 VDD.n1329 VDD.n1169 4.5005
R81317 VDD.n1360 VDD.n1169 4.5005
R81318 VDD.n1328 VDD.n1169 4.5005
R81319 VDD.n1362 VDD.n1169 4.5005
R81320 VDD.n1327 VDD.n1169 4.5005
R81321 VDD.n1363 VDD.n1169 4.5005
R81322 VDD.n1326 VDD.n1169 4.5005
R81323 VDD.n1365 VDD.n1169 4.5005
R81324 VDD.n1325 VDD.n1169 4.5005
R81325 VDD.n1366 VDD.n1169 4.5005
R81326 VDD.n1324 VDD.n1169 4.5005
R81327 VDD.n1368 VDD.n1169 4.5005
R81328 VDD.n1323 VDD.n1169 4.5005
R81329 VDD.n1369 VDD.n1169 4.5005
R81330 VDD.n1322 VDD.n1169 4.5005
R81331 VDD.n1371 VDD.n1169 4.5005
R81332 VDD.n1321 VDD.n1169 4.5005
R81333 VDD.n1372 VDD.n1169 4.5005
R81334 VDD.n1320 VDD.n1169 4.5005
R81335 VDD.n1374 VDD.n1169 4.5005
R81336 VDD.n1319 VDD.n1169 4.5005
R81337 VDD.n1375 VDD.n1169 4.5005
R81338 VDD.n1318 VDD.n1169 4.5005
R81339 VDD.n1376 VDD.n1169 4.5005
R81340 VDD.n1316 VDD.n1169 4.5005
R81341 VDD.n1377 VDD.n1169 4.5005
R81342 VDD.n1315 VDD.n1169 4.5005
R81343 VDD.n1378 VDD.n1169 4.5005
R81344 VDD.n1313 VDD.n1169 4.5005
R81345 VDD.n1379 VDD.n1169 4.5005
R81346 VDD.n1312 VDD.n1169 4.5005
R81347 VDD.n1380 VDD.n1169 4.5005
R81348 VDD.n1310 VDD.n1169 4.5005
R81349 VDD.n1381 VDD.n1169 4.5005
R81350 VDD.n1309 VDD.n1169 4.5005
R81351 VDD.n1382 VDD.n1169 4.5005
R81352 VDD.n1307 VDD.n1169 4.5005
R81353 VDD.n1383 VDD.n1169 4.5005
R81354 VDD.n1306 VDD.n1169 4.5005
R81355 VDD.n1384 VDD.n1169 4.5005
R81356 VDD.n1304 VDD.n1169 4.5005
R81357 VDD.n1385 VDD.n1169 4.5005
R81358 VDD.n1303 VDD.n1169 4.5005
R81359 VDD.n1386 VDD.n1169 4.5005
R81360 VDD.n1301 VDD.n1169 4.5005
R81361 VDD.n1387 VDD.n1169 4.5005
R81362 VDD.n1300 VDD.n1169 4.5005
R81363 VDD.n1388 VDD.n1169 4.5005
R81364 VDD.n1298 VDD.n1169 4.5005
R81365 VDD.n1389 VDD.n1169 4.5005
R81366 VDD.n1297 VDD.n1169 4.5005
R81367 VDD.n1390 VDD.n1169 4.5005
R81368 VDD.n1295 VDD.n1169 4.5005
R81369 VDD.n1391 VDD.n1169 4.5005
R81370 VDD.n1294 VDD.n1169 4.5005
R81371 VDD.n1392 VDD.n1169 4.5005
R81372 VDD.n1292 VDD.n1169 4.5005
R81373 VDD.n1393 VDD.n1169 4.5005
R81374 VDD.n1291 VDD.n1169 4.5005
R81375 VDD.n1394 VDD.n1169 4.5005
R81376 VDD.n1289 VDD.n1169 4.5005
R81377 VDD.n1395 VDD.n1169 4.5005
R81378 VDD.n1288 VDD.n1169 4.5005
R81379 VDD.n1396 VDD.n1169 4.5005
R81380 VDD.n1286 VDD.n1169 4.5005
R81381 VDD.n1397 VDD.n1169 4.5005
R81382 VDD.n1285 VDD.n1169 4.5005
R81383 VDD.n1398 VDD.n1169 4.5005
R81384 VDD.n1283 VDD.n1169 4.5005
R81385 VDD.n1399 VDD.n1169 4.5005
R81386 VDD.n1282 VDD.n1169 4.5005
R81387 VDD.n1400 VDD.n1169 4.5005
R81388 VDD.n1280 VDD.n1169 4.5005
R81389 VDD.n1401 VDD.n1169 4.5005
R81390 VDD.n1279 VDD.n1169 4.5005
R81391 VDD.n1402 VDD.n1169 4.5005
R81392 VDD.n1277 VDD.n1169 4.5005
R81393 VDD.n1403 VDD.n1169 4.5005
R81394 VDD.n1276 VDD.n1169 4.5005
R81395 VDD.n1404 VDD.n1169 4.5005
R81396 VDD.n1274 VDD.n1169 4.5005
R81397 VDD.n1405 VDD.n1169 4.5005
R81398 VDD.n1273 VDD.n1169 4.5005
R81399 VDD.n1406 VDD.n1169 4.5005
R81400 VDD.n1271 VDD.n1169 4.5005
R81401 VDD.n1407 VDD.n1169 4.5005
R81402 VDD.n1270 VDD.n1169 4.5005
R81403 VDD.n1408 VDD.n1169 4.5005
R81404 VDD.n1268 VDD.n1169 4.5005
R81405 VDD.n1409 VDD.n1169 4.5005
R81406 VDD.n1267 VDD.n1169 4.5005
R81407 VDD.n1410 VDD.n1169 4.5005
R81408 VDD.n1265 VDD.n1169 4.5005
R81409 VDD.n1411 VDD.n1169 4.5005
R81410 VDD.n1264 VDD.n1169 4.5005
R81411 VDD.n1412 VDD.n1169 4.5005
R81412 VDD.n1262 VDD.n1169 4.5005
R81413 VDD.n1413 VDD.n1169 4.5005
R81414 VDD.n1261 VDD.n1169 4.5005
R81415 VDD.n1414 VDD.n1169 4.5005
R81416 VDD.n1415 VDD.n1169 4.5005
R81417 VDD.n1674 VDD.n1169 4.5005
R81418 VDD.n1676 VDD.n1221 4.5005
R81419 VDD.n1341 VDD.n1221 4.5005
R81420 VDD.n1342 VDD.n1221 4.5005
R81421 VDD.n1340 VDD.n1221 4.5005
R81422 VDD.n1344 VDD.n1221 4.5005
R81423 VDD.n1339 VDD.n1221 4.5005
R81424 VDD.n1345 VDD.n1221 4.5005
R81425 VDD.n1338 VDD.n1221 4.5005
R81426 VDD.n1347 VDD.n1221 4.5005
R81427 VDD.n1337 VDD.n1221 4.5005
R81428 VDD.n1348 VDD.n1221 4.5005
R81429 VDD.n1336 VDD.n1221 4.5005
R81430 VDD.n1350 VDD.n1221 4.5005
R81431 VDD.n1335 VDD.n1221 4.5005
R81432 VDD.n1351 VDD.n1221 4.5005
R81433 VDD.n1334 VDD.n1221 4.5005
R81434 VDD.n1353 VDD.n1221 4.5005
R81435 VDD.n1333 VDD.n1221 4.5005
R81436 VDD.n1354 VDD.n1221 4.5005
R81437 VDD.n1332 VDD.n1221 4.5005
R81438 VDD.n1356 VDD.n1221 4.5005
R81439 VDD.n1331 VDD.n1221 4.5005
R81440 VDD.n1357 VDD.n1221 4.5005
R81441 VDD.n1330 VDD.n1221 4.5005
R81442 VDD.n1359 VDD.n1221 4.5005
R81443 VDD.n1329 VDD.n1221 4.5005
R81444 VDD.n1360 VDD.n1221 4.5005
R81445 VDD.n1328 VDD.n1221 4.5005
R81446 VDD.n1362 VDD.n1221 4.5005
R81447 VDD.n1327 VDD.n1221 4.5005
R81448 VDD.n1363 VDD.n1221 4.5005
R81449 VDD.n1326 VDD.n1221 4.5005
R81450 VDD.n1365 VDD.n1221 4.5005
R81451 VDD.n1325 VDD.n1221 4.5005
R81452 VDD.n1366 VDD.n1221 4.5005
R81453 VDD.n1324 VDD.n1221 4.5005
R81454 VDD.n1368 VDD.n1221 4.5005
R81455 VDD.n1323 VDD.n1221 4.5005
R81456 VDD.n1369 VDD.n1221 4.5005
R81457 VDD.n1322 VDD.n1221 4.5005
R81458 VDD.n1371 VDD.n1221 4.5005
R81459 VDD.n1321 VDD.n1221 4.5005
R81460 VDD.n1372 VDD.n1221 4.5005
R81461 VDD.n1320 VDD.n1221 4.5005
R81462 VDD.n1374 VDD.n1221 4.5005
R81463 VDD.n1319 VDD.n1221 4.5005
R81464 VDD.n1375 VDD.n1221 4.5005
R81465 VDD.n1318 VDD.n1221 4.5005
R81466 VDD.n1376 VDD.n1221 4.5005
R81467 VDD.n1316 VDD.n1221 4.5005
R81468 VDD.n1377 VDD.n1221 4.5005
R81469 VDD.n1315 VDD.n1221 4.5005
R81470 VDD.n1378 VDD.n1221 4.5005
R81471 VDD.n1313 VDD.n1221 4.5005
R81472 VDD.n1379 VDD.n1221 4.5005
R81473 VDD.n1312 VDD.n1221 4.5005
R81474 VDD.n1380 VDD.n1221 4.5005
R81475 VDD.n1310 VDD.n1221 4.5005
R81476 VDD.n1381 VDD.n1221 4.5005
R81477 VDD.n1309 VDD.n1221 4.5005
R81478 VDD.n1382 VDD.n1221 4.5005
R81479 VDD.n1307 VDD.n1221 4.5005
R81480 VDD.n1383 VDD.n1221 4.5005
R81481 VDD.n1306 VDD.n1221 4.5005
R81482 VDD.n1384 VDD.n1221 4.5005
R81483 VDD.n1304 VDD.n1221 4.5005
R81484 VDD.n1385 VDD.n1221 4.5005
R81485 VDD.n1303 VDD.n1221 4.5005
R81486 VDD.n1386 VDD.n1221 4.5005
R81487 VDD.n1301 VDD.n1221 4.5005
R81488 VDD.n1387 VDD.n1221 4.5005
R81489 VDD.n1300 VDD.n1221 4.5005
R81490 VDD.n1388 VDD.n1221 4.5005
R81491 VDD.n1298 VDD.n1221 4.5005
R81492 VDD.n1389 VDD.n1221 4.5005
R81493 VDD.n1297 VDD.n1221 4.5005
R81494 VDD.n1390 VDD.n1221 4.5005
R81495 VDD.n1295 VDD.n1221 4.5005
R81496 VDD.n1391 VDD.n1221 4.5005
R81497 VDD.n1294 VDD.n1221 4.5005
R81498 VDD.n1392 VDD.n1221 4.5005
R81499 VDD.n1292 VDD.n1221 4.5005
R81500 VDD.n1393 VDD.n1221 4.5005
R81501 VDD.n1291 VDD.n1221 4.5005
R81502 VDD.n1394 VDD.n1221 4.5005
R81503 VDD.n1289 VDD.n1221 4.5005
R81504 VDD.n1395 VDD.n1221 4.5005
R81505 VDD.n1288 VDD.n1221 4.5005
R81506 VDD.n1396 VDD.n1221 4.5005
R81507 VDD.n1286 VDD.n1221 4.5005
R81508 VDD.n1397 VDD.n1221 4.5005
R81509 VDD.n1285 VDD.n1221 4.5005
R81510 VDD.n1398 VDD.n1221 4.5005
R81511 VDD.n1283 VDD.n1221 4.5005
R81512 VDD.n1399 VDD.n1221 4.5005
R81513 VDD.n1282 VDD.n1221 4.5005
R81514 VDD.n1400 VDD.n1221 4.5005
R81515 VDD.n1280 VDD.n1221 4.5005
R81516 VDD.n1401 VDD.n1221 4.5005
R81517 VDD.n1279 VDD.n1221 4.5005
R81518 VDD.n1402 VDD.n1221 4.5005
R81519 VDD.n1277 VDD.n1221 4.5005
R81520 VDD.n1403 VDD.n1221 4.5005
R81521 VDD.n1276 VDD.n1221 4.5005
R81522 VDD.n1404 VDD.n1221 4.5005
R81523 VDD.n1274 VDD.n1221 4.5005
R81524 VDD.n1405 VDD.n1221 4.5005
R81525 VDD.n1273 VDD.n1221 4.5005
R81526 VDD.n1406 VDD.n1221 4.5005
R81527 VDD.n1271 VDD.n1221 4.5005
R81528 VDD.n1407 VDD.n1221 4.5005
R81529 VDD.n1270 VDD.n1221 4.5005
R81530 VDD.n1408 VDD.n1221 4.5005
R81531 VDD.n1268 VDD.n1221 4.5005
R81532 VDD.n1409 VDD.n1221 4.5005
R81533 VDD.n1267 VDD.n1221 4.5005
R81534 VDD.n1410 VDD.n1221 4.5005
R81535 VDD.n1265 VDD.n1221 4.5005
R81536 VDD.n1411 VDD.n1221 4.5005
R81537 VDD.n1264 VDD.n1221 4.5005
R81538 VDD.n1412 VDD.n1221 4.5005
R81539 VDD.n1262 VDD.n1221 4.5005
R81540 VDD.n1413 VDD.n1221 4.5005
R81541 VDD.n1261 VDD.n1221 4.5005
R81542 VDD.n1414 VDD.n1221 4.5005
R81543 VDD.n1415 VDD.n1221 4.5005
R81544 VDD.n1674 VDD.n1221 4.5005
R81545 VDD.n1676 VDD.n1168 4.5005
R81546 VDD.n1341 VDD.n1168 4.5005
R81547 VDD.n1342 VDD.n1168 4.5005
R81548 VDD.n1340 VDD.n1168 4.5005
R81549 VDD.n1344 VDD.n1168 4.5005
R81550 VDD.n1339 VDD.n1168 4.5005
R81551 VDD.n1345 VDD.n1168 4.5005
R81552 VDD.n1338 VDD.n1168 4.5005
R81553 VDD.n1347 VDD.n1168 4.5005
R81554 VDD.n1337 VDD.n1168 4.5005
R81555 VDD.n1348 VDD.n1168 4.5005
R81556 VDD.n1336 VDD.n1168 4.5005
R81557 VDD.n1350 VDD.n1168 4.5005
R81558 VDD.n1335 VDD.n1168 4.5005
R81559 VDD.n1351 VDD.n1168 4.5005
R81560 VDD.n1334 VDD.n1168 4.5005
R81561 VDD.n1353 VDD.n1168 4.5005
R81562 VDD.n1333 VDD.n1168 4.5005
R81563 VDD.n1354 VDD.n1168 4.5005
R81564 VDD.n1332 VDD.n1168 4.5005
R81565 VDD.n1356 VDD.n1168 4.5005
R81566 VDD.n1331 VDD.n1168 4.5005
R81567 VDD.n1357 VDD.n1168 4.5005
R81568 VDD.n1330 VDD.n1168 4.5005
R81569 VDD.n1359 VDD.n1168 4.5005
R81570 VDD.n1329 VDD.n1168 4.5005
R81571 VDD.n1360 VDD.n1168 4.5005
R81572 VDD.n1328 VDD.n1168 4.5005
R81573 VDD.n1362 VDD.n1168 4.5005
R81574 VDD.n1327 VDD.n1168 4.5005
R81575 VDD.n1363 VDD.n1168 4.5005
R81576 VDD.n1326 VDD.n1168 4.5005
R81577 VDD.n1365 VDD.n1168 4.5005
R81578 VDD.n1325 VDD.n1168 4.5005
R81579 VDD.n1366 VDD.n1168 4.5005
R81580 VDD.n1324 VDD.n1168 4.5005
R81581 VDD.n1368 VDD.n1168 4.5005
R81582 VDD.n1323 VDD.n1168 4.5005
R81583 VDD.n1369 VDD.n1168 4.5005
R81584 VDD.n1322 VDD.n1168 4.5005
R81585 VDD.n1371 VDD.n1168 4.5005
R81586 VDD.n1321 VDD.n1168 4.5005
R81587 VDD.n1372 VDD.n1168 4.5005
R81588 VDD.n1320 VDD.n1168 4.5005
R81589 VDD.n1374 VDD.n1168 4.5005
R81590 VDD.n1319 VDD.n1168 4.5005
R81591 VDD.n1375 VDD.n1168 4.5005
R81592 VDD.n1318 VDD.n1168 4.5005
R81593 VDD.n1376 VDD.n1168 4.5005
R81594 VDD.n1316 VDD.n1168 4.5005
R81595 VDD.n1377 VDD.n1168 4.5005
R81596 VDD.n1315 VDD.n1168 4.5005
R81597 VDD.n1378 VDD.n1168 4.5005
R81598 VDD.n1313 VDD.n1168 4.5005
R81599 VDD.n1379 VDD.n1168 4.5005
R81600 VDD.n1312 VDD.n1168 4.5005
R81601 VDD.n1380 VDD.n1168 4.5005
R81602 VDD.n1310 VDD.n1168 4.5005
R81603 VDD.n1381 VDD.n1168 4.5005
R81604 VDD.n1309 VDD.n1168 4.5005
R81605 VDD.n1382 VDD.n1168 4.5005
R81606 VDD.n1307 VDD.n1168 4.5005
R81607 VDD.n1383 VDD.n1168 4.5005
R81608 VDD.n1306 VDD.n1168 4.5005
R81609 VDD.n1384 VDD.n1168 4.5005
R81610 VDD.n1304 VDD.n1168 4.5005
R81611 VDD.n1385 VDD.n1168 4.5005
R81612 VDD.n1303 VDD.n1168 4.5005
R81613 VDD.n1386 VDD.n1168 4.5005
R81614 VDD.n1301 VDD.n1168 4.5005
R81615 VDD.n1387 VDD.n1168 4.5005
R81616 VDD.n1300 VDD.n1168 4.5005
R81617 VDD.n1388 VDD.n1168 4.5005
R81618 VDD.n1298 VDD.n1168 4.5005
R81619 VDD.n1389 VDD.n1168 4.5005
R81620 VDD.n1297 VDD.n1168 4.5005
R81621 VDD.n1390 VDD.n1168 4.5005
R81622 VDD.n1295 VDD.n1168 4.5005
R81623 VDD.n1391 VDD.n1168 4.5005
R81624 VDD.n1294 VDD.n1168 4.5005
R81625 VDD.n1392 VDD.n1168 4.5005
R81626 VDD.n1292 VDD.n1168 4.5005
R81627 VDD.n1393 VDD.n1168 4.5005
R81628 VDD.n1291 VDD.n1168 4.5005
R81629 VDD.n1394 VDD.n1168 4.5005
R81630 VDD.n1289 VDD.n1168 4.5005
R81631 VDD.n1395 VDD.n1168 4.5005
R81632 VDD.n1288 VDD.n1168 4.5005
R81633 VDD.n1396 VDD.n1168 4.5005
R81634 VDD.n1286 VDD.n1168 4.5005
R81635 VDD.n1397 VDD.n1168 4.5005
R81636 VDD.n1285 VDD.n1168 4.5005
R81637 VDD.n1398 VDD.n1168 4.5005
R81638 VDD.n1283 VDD.n1168 4.5005
R81639 VDD.n1399 VDD.n1168 4.5005
R81640 VDD.n1282 VDD.n1168 4.5005
R81641 VDD.n1400 VDD.n1168 4.5005
R81642 VDD.n1280 VDD.n1168 4.5005
R81643 VDD.n1401 VDD.n1168 4.5005
R81644 VDD.n1279 VDD.n1168 4.5005
R81645 VDD.n1402 VDD.n1168 4.5005
R81646 VDD.n1277 VDD.n1168 4.5005
R81647 VDD.n1403 VDD.n1168 4.5005
R81648 VDD.n1276 VDD.n1168 4.5005
R81649 VDD.n1404 VDD.n1168 4.5005
R81650 VDD.n1274 VDD.n1168 4.5005
R81651 VDD.n1405 VDD.n1168 4.5005
R81652 VDD.n1273 VDD.n1168 4.5005
R81653 VDD.n1406 VDD.n1168 4.5005
R81654 VDD.n1271 VDD.n1168 4.5005
R81655 VDD.n1407 VDD.n1168 4.5005
R81656 VDD.n1270 VDD.n1168 4.5005
R81657 VDD.n1408 VDD.n1168 4.5005
R81658 VDD.n1268 VDD.n1168 4.5005
R81659 VDD.n1409 VDD.n1168 4.5005
R81660 VDD.n1267 VDD.n1168 4.5005
R81661 VDD.n1410 VDD.n1168 4.5005
R81662 VDD.n1265 VDD.n1168 4.5005
R81663 VDD.n1411 VDD.n1168 4.5005
R81664 VDD.n1264 VDD.n1168 4.5005
R81665 VDD.n1412 VDD.n1168 4.5005
R81666 VDD.n1262 VDD.n1168 4.5005
R81667 VDD.n1413 VDD.n1168 4.5005
R81668 VDD.n1261 VDD.n1168 4.5005
R81669 VDD.n1414 VDD.n1168 4.5005
R81670 VDD.n1415 VDD.n1168 4.5005
R81671 VDD.n1674 VDD.n1168 4.5005
R81672 VDD.n1676 VDD.n1222 4.5005
R81673 VDD.n1341 VDD.n1222 4.5005
R81674 VDD.n1342 VDD.n1222 4.5005
R81675 VDD.n1340 VDD.n1222 4.5005
R81676 VDD.n1344 VDD.n1222 4.5005
R81677 VDD.n1339 VDD.n1222 4.5005
R81678 VDD.n1345 VDD.n1222 4.5005
R81679 VDD.n1338 VDD.n1222 4.5005
R81680 VDD.n1347 VDD.n1222 4.5005
R81681 VDD.n1337 VDD.n1222 4.5005
R81682 VDD.n1348 VDD.n1222 4.5005
R81683 VDD.n1336 VDD.n1222 4.5005
R81684 VDD.n1350 VDD.n1222 4.5005
R81685 VDD.n1335 VDD.n1222 4.5005
R81686 VDD.n1351 VDD.n1222 4.5005
R81687 VDD.n1334 VDD.n1222 4.5005
R81688 VDD.n1353 VDD.n1222 4.5005
R81689 VDD.n1333 VDD.n1222 4.5005
R81690 VDD.n1354 VDD.n1222 4.5005
R81691 VDD.n1332 VDD.n1222 4.5005
R81692 VDD.n1356 VDD.n1222 4.5005
R81693 VDD.n1331 VDD.n1222 4.5005
R81694 VDD.n1357 VDD.n1222 4.5005
R81695 VDD.n1330 VDD.n1222 4.5005
R81696 VDD.n1359 VDD.n1222 4.5005
R81697 VDD.n1329 VDD.n1222 4.5005
R81698 VDD.n1360 VDD.n1222 4.5005
R81699 VDD.n1328 VDD.n1222 4.5005
R81700 VDD.n1362 VDD.n1222 4.5005
R81701 VDD.n1327 VDD.n1222 4.5005
R81702 VDD.n1363 VDD.n1222 4.5005
R81703 VDD.n1326 VDD.n1222 4.5005
R81704 VDD.n1365 VDD.n1222 4.5005
R81705 VDD.n1325 VDD.n1222 4.5005
R81706 VDD.n1366 VDD.n1222 4.5005
R81707 VDD.n1324 VDD.n1222 4.5005
R81708 VDD.n1368 VDD.n1222 4.5005
R81709 VDD.n1323 VDD.n1222 4.5005
R81710 VDD.n1369 VDD.n1222 4.5005
R81711 VDD.n1322 VDD.n1222 4.5005
R81712 VDD.n1371 VDD.n1222 4.5005
R81713 VDD.n1321 VDD.n1222 4.5005
R81714 VDD.n1372 VDD.n1222 4.5005
R81715 VDD.n1320 VDD.n1222 4.5005
R81716 VDD.n1374 VDD.n1222 4.5005
R81717 VDD.n1319 VDD.n1222 4.5005
R81718 VDD.n1375 VDD.n1222 4.5005
R81719 VDD.n1318 VDD.n1222 4.5005
R81720 VDD.n1376 VDD.n1222 4.5005
R81721 VDD.n1316 VDD.n1222 4.5005
R81722 VDD.n1377 VDD.n1222 4.5005
R81723 VDD.n1315 VDD.n1222 4.5005
R81724 VDD.n1378 VDD.n1222 4.5005
R81725 VDD.n1313 VDD.n1222 4.5005
R81726 VDD.n1379 VDD.n1222 4.5005
R81727 VDD.n1312 VDD.n1222 4.5005
R81728 VDD.n1380 VDD.n1222 4.5005
R81729 VDD.n1310 VDD.n1222 4.5005
R81730 VDD.n1381 VDD.n1222 4.5005
R81731 VDD.n1309 VDD.n1222 4.5005
R81732 VDD.n1382 VDD.n1222 4.5005
R81733 VDD.n1307 VDD.n1222 4.5005
R81734 VDD.n1383 VDD.n1222 4.5005
R81735 VDD.n1306 VDD.n1222 4.5005
R81736 VDD.n1384 VDD.n1222 4.5005
R81737 VDD.n1304 VDD.n1222 4.5005
R81738 VDD.n1385 VDD.n1222 4.5005
R81739 VDD.n1303 VDD.n1222 4.5005
R81740 VDD.n1386 VDD.n1222 4.5005
R81741 VDD.n1301 VDD.n1222 4.5005
R81742 VDD.n1387 VDD.n1222 4.5005
R81743 VDD.n1300 VDD.n1222 4.5005
R81744 VDD.n1388 VDD.n1222 4.5005
R81745 VDD.n1298 VDD.n1222 4.5005
R81746 VDD.n1389 VDD.n1222 4.5005
R81747 VDD.n1297 VDD.n1222 4.5005
R81748 VDD.n1390 VDD.n1222 4.5005
R81749 VDD.n1295 VDD.n1222 4.5005
R81750 VDD.n1391 VDD.n1222 4.5005
R81751 VDD.n1294 VDD.n1222 4.5005
R81752 VDD.n1392 VDD.n1222 4.5005
R81753 VDD.n1292 VDD.n1222 4.5005
R81754 VDD.n1393 VDD.n1222 4.5005
R81755 VDD.n1291 VDD.n1222 4.5005
R81756 VDD.n1394 VDD.n1222 4.5005
R81757 VDD.n1289 VDD.n1222 4.5005
R81758 VDD.n1395 VDD.n1222 4.5005
R81759 VDD.n1288 VDD.n1222 4.5005
R81760 VDD.n1396 VDD.n1222 4.5005
R81761 VDD.n1286 VDD.n1222 4.5005
R81762 VDD.n1397 VDD.n1222 4.5005
R81763 VDD.n1285 VDD.n1222 4.5005
R81764 VDD.n1398 VDD.n1222 4.5005
R81765 VDD.n1283 VDD.n1222 4.5005
R81766 VDD.n1399 VDD.n1222 4.5005
R81767 VDD.n1282 VDD.n1222 4.5005
R81768 VDD.n1400 VDD.n1222 4.5005
R81769 VDD.n1280 VDD.n1222 4.5005
R81770 VDD.n1401 VDD.n1222 4.5005
R81771 VDD.n1279 VDD.n1222 4.5005
R81772 VDD.n1402 VDD.n1222 4.5005
R81773 VDD.n1277 VDD.n1222 4.5005
R81774 VDD.n1403 VDD.n1222 4.5005
R81775 VDD.n1276 VDD.n1222 4.5005
R81776 VDD.n1404 VDD.n1222 4.5005
R81777 VDD.n1274 VDD.n1222 4.5005
R81778 VDD.n1405 VDD.n1222 4.5005
R81779 VDD.n1273 VDD.n1222 4.5005
R81780 VDD.n1406 VDD.n1222 4.5005
R81781 VDD.n1271 VDD.n1222 4.5005
R81782 VDD.n1407 VDD.n1222 4.5005
R81783 VDD.n1270 VDD.n1222 4.5005
R81784 VDD.n1408 VDD.n1222 4.5005
R81785 VDD.n1268 VDD.n1222 4.5005
R81786 VDD.n1409 VDD.n1222 4.5005
R81787 VDD.n1267 VDD.n1222 4.5005
R81788 VDD.n1410 VDD.n1222 4.5005
R81789 VDD.n1265 VDD.n1222 4.5005
R81790 VDD.n1411 VDD.n1222 4.5005
R81791 VDD.n1264 VDD.n1222 4.5005
R81792 VDD.n1412 VDD.n1222 4.5005
R81793 VDD.n1262 VDD.n1222 4.5005
R81794 VDD.n1413 VDD.n1222 4.5005
R81795 VDD.n1261 VDD.n1222 4.5005
R81796 VDD.n1414 VDD.n1222 4.5005
R81797 VDD.n1415 VDD.n1222 4.5005
R81798 VDD.n1674 VDD.n1222 4.5005
R81799 VDD.n1676 VDD.n1167 4.5005
R81800 VDD.n1341 VDD.n1167 4.5005
R81801 VDD.n1342 VDD.n1167 4.5005
R81802 VDD.n1340 VDD.n1167 4.5005
R81803 VDD.n1344 VDD.n1167 4.5005
R81804 VDD.n1339 VDD.n1167 4.5005
R81805 VDD.n1345 VDD.n1167 4.5005
R81806 VDD.n1338 VDD.n1167 4.5005
R81807 VDD.n1347 VDD.n1167 4.5005
R81808 VDD.n1337 VDD.n1167 4.5005
R81809 VDD.n1348 VDD.n1167 4.5005
R81810 VDD.n1336 VDD.n1167 4.5005
R81811 VDD.n1350 VDD.n1167 4.5005
R81812 VDD.n1335 VDD.n1167 4.5005
R81813 VDD.n1351 VDD.n1167 4.5005
R81814 VDD.n1334 VDD.n1167 4.5005
R81815 VDD.n1353 VDD.n1167 4.5005
R81816 VDD.n1333 VDD.n1167 4.5005
R81817 VDD.n1354 VDD.n1167 4.5005
R81818 VDD.n1332 VDD.n1167 4.5005
R81819 VDD.n1356 VDD.n1167 4.5005
R81820 VDD.n1331 VDD.n1167 4.5005
R81821 VDD.n1357 VDD.n1167 4.5005
R81822 VDD.n1330 VDD.n1167 4.5005
R81823 VDD.n1359 VDD.n1167 4.5005
R81824 VDD.n1329 VDD.n1167 4.5005
R81825 VDD.n1360 VDD.n1167 4.5005
R81826 VDD.n1328 VDD.n1167 4.5005
R81827 VDD.n1362 VDD.n1167 4.5005
R81828 VDD.n1327 VDD.n1167 4.5005
R81829 VDD.n1363 VDD.n1167 4.5005
R81830 VDD.n1326 VDD.n1167 4.5005
R81831 VDD.n1365 VDD.n1167 4.5005
R81832 VDD.n1325 VDD.n1167 4.5005
R81833 VDD.n1366 VDD.n1167 4.5005
R81834 VDD.n1324 VDD.n1167 4.5005
R81835 VDD.n1368 VDD.n1167 4.5005
R81836 VDD.n1323 VDD.n1167 4.5005
R81837 VDD.n1369 VDD.n1167 4.5005
R81838 VDD.n1322 VDD.n1167 4.5005
R81839 VDD.n1371 VDD.n1167 4.5005
R81840 VDD.n1321 VDD.n1167 4.5005
R81841 VDD.n1372 VDD.n1167 4.5005
R81842 VDD.n1320 VDD.n1167 4.5005
R81843 VDD.n1374 VDD.n1167 4.5005
R81844 VDD.n1319 VDD.n1167 4.5005
R81845 VDD.n1375 VDD.n1167 4.5005
R81846 VDD.n1318 VDD.n1167 4.5005
R81847 VDD.n1376 VDD.n1167 4.5005
R81848 VDD.n1316 VDD.n1167 4.5005
R81849 VDD.n1377 VDD.n1167 4.5005
R81850 VDD.n1315 VDD.n1167 4.5005
R81851 VDD.n1378 VDD.n1167 4.5005
R81852 VDD.n1313 VDD.n1167 4.5005
R81853 VDD.n1379 VDD.n1167 4.5005
R81854 VDD.n1312 VDD.n1167 4.5005
R81855 VDD.n1380 VDD.n1167 4.5005
R81856 VDD.n1310 VDD.n1167 4.5005
R81857 VDD.n1381 VDD.n1167 4.5005
R81858 VDD.n1309 VDD.n1167 4.5005
R81859 VDD.n1382 VDD.n1167 4.5005
R81860 VDD.n1307 VDD.n1167 4.5005
R81861 VDD.n1383 VDD.n1167 4.5005
R81862 VDD.n1306 VDD.n1167 4.5005
R81863 VDD.n1384 VDD.n1167 4.5005
R81864 VDD.n1304 VDD.n1167 4.5005
R81865 VDD.n1385 VDD.n1167 4.5005
R81866 VDD.n1303 VDD.n1167 4.5005
R81867 VDD.n1386 VDD.n1167 4.5005
R81868 VDD.n1301 VDD.n1167 4.5005
R81869 VDD.n1387 VDD.n1167 4.5005
R81870 VDD.n1300 VDD.n1167 4.5005
R81871 VDD.n1388 VDD.n1167 4.5005
R81872 VDD.n1298 VDD.n1167 4.5005
R81873 VDD.n1389 VDD.n1167 4.5005
R81874 VDD.n1297 VDD.n1167 4.5005
R81875 VDD.n1390 VDD.n1167 4.5005
R81876 VDD.n1295 VDD.n1167 4.5005
R81877 VDD.n1391 VDD.n1167 4.5005
R81878 VDD.n1294 VDD.n1167 4.5005
R81879 VDD.n1392 VDD.n1167 4.5005
R81880 VDD.n1292 VDD.n1167 4.5005
R81881 VDD.n1393 VDD.n1167 4.5005
R81882 VDD.n1291 VDD.n1167 4.5005
R81883 VDD.n1394 VDD.n1167 4.5005
R81884 VDD.n1289 VDD.n1167 4.5005
R81885 VDD.n1395 VDD.n1167 4.5005
R81886 VDD.n1288 VDD.n1167 4.5005
R81887 VDD.n1396 VDD.n1167 4.5005
R81888 VDD.n1286 VDD.n1167 4.5005
R81889 VDD.n1397 VDD.n1167 4.5005
R81890 VDD.n1285 VDD.n1167 4.5005
R81891 VDD.n1398 VDD.n1167 4.5005
R81892 VDD.n1283 VDD.n1167 4.5005
R81893 VDD.n1399 VDD.n1167 4.5005
R81894 VDD.n1282 VDD.n1167 4.5005
R81895 VDD.n1400 VDD.n1167 4.5005
R81896 VDD.n1280 VDD.n1167 4.5005
R81897 VDD.n1401 VDD.n1167 4.5005
R81898 VDD.n1279 VDD.n1167 4.5005
R81899 VDD.n1402 VDD.n1167 4.5005
R81900 VDD.n1277 VDD.n1167 4.5005
R81901 VDD.n1403 VDD.n1167 4.5005
R81902 VDD.n1276 VDD.n1167 4.5005
R81903 VDD.n1404 VDD.n1167 4.5005
R81904 VDD.n1274 VDD.n1167 4.5005
R81905 VDD.n1405 VDD.n1167 4.5005
R81906 VDD.n1273 VDD.n1167 4.5005
R81907 VDD.n1406 VDD.n1167 4.5005
R81908 VDD.n1271 VDD.n1167 4.5005
R81909 VDD.n1407 VDD.n1167 4.5005
R81910 VDD.n1270 VDD.n1167 4.5005
R81911 VDD.n1408 VDD.n1167 4.5005
R81912 VDD.n1268 VDD.n1167 4.5005
R81913 VDD.n1409 VDD.n1167 4.5005
R81914 VDD.n1267 VDD.n1167 4.5005
R81915 VDD.n1410 VDD.n1167 4.5005
R81916 VDD.n1265 VDD.n1167 4.5005
R81917 VDD.n1411 VDD.n1167 4.5005
R81918 VDD.n1264 VDD.n1167 4.5005
R81919 VDD.n1412 VDD.n1167 4.5005
R81920 VDD.n1262 VDD.n1167 4.5005
R81921 VDD.n1413 VDD.n1167 4.5005
R81922 VDD.n1261 VDD.n1167 4.5005
R81923 VDD.n1414 VDD.n1167 4.5005
R81924 VDD.n1415 VDD.n1167 4.5005
R81925 VDD.n1674 VDD.n1167 4.5005
R81926 VDD.n1676 VDD.n1223 4.5005
R81927 VDD.n1341 VDD.n1223 4.5005
R81928 VDD.n1342 VDD.n1223 4.5005
R81929 VDD.n1340 VDD.n1223 4.5005
R81930 VDD.n1344 VDD.n1223 4.5005
R81931 VDD.n1339 VDD.n1223 4.5005
R81932 VDD.n1345 VDD.n1223 4.5005
R81933 VDD.n1338 VDD.n1223 4.5005
R81934 VDD.n1347 VDD.n1223 4.5005
R81935 VDD.n1337 VDD.n1223 4.5005
R81936 VDD.n1348 VDD.n1223 4.5005
R81937 VDD.n1336 VDD.n1223 4.5005
R81938 VDD.n1350 VDD.n1223 4.5005
R81939 VDD.n1335 VDD.n1223 4.5005
R81940 VDD.n1351 VDD.n1223 4.5005
R81941 VDD.n1334 VDD.n1223 4.5005
R81942 VDD.n1353 VDD.n1223 4.5005
R81943 VDD.n1333 VDD.n1223 4.5005
R81944 VDD.n1354 VDD.n1223 4.5005
R81945 VDD.n1332 VDD.n1223 4.5005
R81946 VDD.n1356 VDD.n1223 4.5005
R81947 VDD.n1331 VDD.n1223 4.5005
R81948 VDD.n1357 VDD.n1223 4.5005
R81949 VDD.n1330 VDD.n1223 4.5005
R81950 VDD.n1359 VDD.n1223 4.5005
R81951 VDD.n1329 VDD.n1223 4.5005
R81952 VDD.n1360 VDD.n1223 4.5005
R81953 VDD.n1328 VDD.n1223 4.5005
R81954 VDD.n1362 VDD.n1223 4.5005
R81955 VDD.n1327 VDD.n1223 4.5005
R81956 VDD.n1363 VDD.n1223 4.5005
R81957 VDD.n1326 VDD.n1223 4.5005
R81958 VDD.n1365 VDD.n1223 4.5005
R81959 VDD.n1325 VDD.n1223 4.5005
R81960 VDD.n1366 VDD.n1223 4.5005
R81961 VDD.n1324 VDD.n1223 4.5005
R81962 VDD.n1368 VDD.n1223 4.5005
R81963 VDD.n1323 VDD.n1223 4.5005
R81964 VDD.n1369 VDD.n1223 4.5005
R81965 VDD.n1322 VDD.n1223 4.5005
R81966 VDD.n1371 VDD.n1223 4.5005
R81967 VDD.n1321 VDD.n1223 4.5005
R81968 VDD.n1372 VDD.n1223 4.5005
R81969 VDD.n1320 VDD.n1223 4.5005
R81970 VDD.n1374 VDD.n1223 4.5005
R81971 VDD.n1319 VDD.n1223 4.5005
R81972 VDD.n1375 VDD.n1223 4.5005
R81973 VDD.n1318 VDD.n1223 4.5005
R81974 VDD.n1376 VDD.n1223 4.5005
R81975 VDD.n1316 VDD.n1223 4.5005
R81976 VDD.n1377 VDD.n1223 4.5005
R81977 VDD.n1315 VDD.n1223 4.5005
R81978 VDD.n1378 VDD.n1223 4.5005
R81979 VDD.n1313 VDD.n1223 4.5005
R81980 VDD.n1379 VDD.n1223 4.5005
R81981 VDD.n1312 VDD.n1223 4.5005
R81982 VDD.n1380 VDD.n1223 4.5005
R81983 VDD.n1310 VDD.n1223 4.5005
R81984 VDD.n1381 VDD.n1223 4.5005
R81985 VDD.n1309 VDD.n1223 4.5005
R81986 VDD.n1382 VDD.n1223 4.5005
R81987 VDD.n1307 VDD.n1223 4.5005
R81988 VDD.n1383 VDD.n1223 4.5005
R81989 VDD.n1306 VDD.n1223 4.5005
R81990 VDD.n1384 VDD.n1223 4.5005
R81991 VDD.n1304 VDD.n1223 4.5005
R81992 VDD.n1385 VDD.n1223 4.5005
R81993 VDD.n1303 VDD.n1223 4.5005
R81994 VDD.n1386 VDD.n1223 4.5005
R81995 VDD.n1301 VDD.n1223 4.5005
R81996 VDD.n1387 VDD.n1223 4.5005
R81997 VDD.n1300 VDD.n1223 4.5005
R81998 VDD.n1388 VDD.n1223 4.5005
R81999 VDD.n1298 VDD.n1223 4.5005
R82000 VDD.n1389 VDD.n1223 4.5005
R82001 VDD.n1297 VDD.n1223 4.5005
R82002 VDD.n1390 VDD.n1223 4.5005
R82003 VDD.n1295 VDD.n1223 4.5005
R82004 VDD.n1391 VDD.n1223 4.5005
R82005 VDD.n1294 VDD.n1223 4.5005
R82006 VDD.n1392 VDD.n1223 4.5005
R82007 VDD.n1292 VDD.n1223 4.5005
R82008 VDD.n1393 VDD.n1223 4.5005
R82009 VDD.n1291 VDD.n1223 4.5005
R82010 VDD.n1394 VDD.n1223 4.5005
R82011 VDD.n1289 VDD.n1223 4.5005
R82012 VDD.n1395 VDD.n1223 4.5005
R82013 VDD.n1288 VDD.n1223 4.5005
R82014 VDD.n1396 VDD.n1223 4.5005
R82015 VDD.n1286 VDD.n1223 4.5005
R82016 VDD.n1397 VDD.n1223 4.5005
R82017 VDD.n1285 VDD.n1223 4.5005
R82018 VDD.n1398 VDD.n1223 4.5005
R82019 VDD.n1283 VDD.n1223 4.5005
R82020 VDD.n1399 VDD.n1223 4.5005
R82021 VDD.n1282 VDD.n1223 4.5005
R82022 VDD.n1400 VDD.n1223 4.5005
R82023 VDD.n1280 VDD.n1223 4.5005
R82024 VDD.n1401 VDD.n1223 4.5005
R82025 VDD.n1279 VDD.n1223 4.5005
R82026 VDD.n1402 VDD.n1223 4.5005
R82027 VDD.n1277 VDD.n1223 4.5005
R82028 VDD.n1403 VDD.n1223 4.5005
R82029 VDD.n1276 VDD.n1223 4.5005
R82030 VDD.n1404 VDD.n1223 4.5005
R82031 VDD.n1274 VDD.n1223 4.5005
R82032 VDD.n1405 VDD.n1223 4.5005
R82033 VDD.n1273 VDD.n1223 4.5005
R82034 VDD.n1406 VDD.n1223 4.5005
R82035 VDD.n1271 VDD.n1223 4.5005
R82036 VDD.n1407 VDD.n1223 4.5005
R82037 VDD.n1270 VDD.n1223 4.5005
R82038 VDD.n1408 VDD.n1223 4.5005
R82039 VDD.n1268 VDD.n1223 4.5005
R82040 VDD.n1409 VDD.n1223 4.5005
R82041 VDD.n1267 VDD.n1223 4.5005
R82042 VDD.n1410 VDD.n1223 4.5005
R82043 VDD.n1265 VDD.n1223 4.5005
R82044 VDD.n1411 VDD.n1223 4.5005
R82045 VDD.n1264 VDD.n1223 4.5005
R82046 VDD.n1412 VDD.n1223 4.5005
R82047 VDD.n1262 VDD.n1223 4.5005
R82048 VDD.n1413 VDD.n1223 4.5005
R82049 VDD.n1261 VDD.n1223 4.5005
R82050 VDD.n1414 VDD.n1223 4.5005
R82051 VDD.n1415 VDD.n1223 4.5005
R82052 VDD.n1674 VDD.n1223 4.5005
R82053 VDD.n1676 VDD.n1166 4.5005
R82054 VDD.n1341 VDD.n1166 4.5005
R82055 VDD.n1342 VDD.n1166 4.5005
R82056 VDD.n1340 VDD.n1166 4.5005
R82057 VDD.n1344 VDD.n1166 4.5005
R82058 VDD.n1339 VDD.n1166 4.5005
R82059 VDD.n1345 VDD.n1166 4.5005
R82060 VDD.n1338 VDD.n1166 4.5005
R82061 VDD.n1347 VDD.n1166 4.5005
R82062 VDD.n1337 VDD.n1166 4.5005
R82063 VDD.n1348 VDD.n1166 4.5005
R82064 VDD.n1336 VDD.n1166 4.5005
R82065 VDD.n1350 VDD.n1166 4.5005
R82066 VDD.n1335 VDD.n1166 4.5005
R82067 VDD.n1351 VDD.n1166 4.5005
R82068 VDD.n1334 VDD.n1166 4.5005
R82069 VDD.n1353 VDD.n1166 4.5005
R82070 VDD.n1333 VDD.n1166 4.5005
R82071 VDD.n1354 VDD.n1166 4.5005
R82072 VDD.n1332 VDD.n1166 4.5005
R82073 VDD.n1356 VDD.n1166 4.5005
R82074 VDD.n1331 VDD.n1166 4.5005
R82075 VDD.n1357 VDD.n1166 4.5005
R82076 VDD.n1330 VDD.n1166 4.5005
R82077 VDD.n1359 VDD.n1166 4.5005
R82078 VDD.n1329 VDD.n1166 4.5005
R82079 VDD.n1360 VDD.n1166 4.5005
R82080 VDD.n1328 VDD.n1166 4.5005
R82081 VDD.n1362 VDD.n1166 4.5005
R82082 VDD.n1327 VDD.n1166 4.5005
R82083 VDD.n1363 VDD.n1166 4.5005
R82084 VDD.n1326 VDD.n1166 4.5005
R82085 VDD.n1365 VDD.n1166 4.5005
R82086 VDD.n1325 VDD.n1166 4.5005
R82087 VDD.n1366 VDD.n1166 4.5005
R82088 VDD.n1324 VDD.n1166 4.5005
R82089 VDD.n1368 VDD.n1166 4.5005
R82090 VDD.n1323 VDD.n1166 4.5005
R82091 VDD.n1369 VDD.n1166 4.5005
R82092 VDD.n1322 VDD.n1166 4.5005
R82093 VDD.n1371 VDD.n1166 4.5005
R82094 VDD.n1321 VDD.n1166 4.5005
R82095 VDD.n1372 VDD.n1166 4.5005
R82096 VDD.n1320 VDD.n1166 4.5005
R82097 VDD.n1374 VDD.n1166 4.5005
R82098 VDD.n1319 VDD.n1166 4.5005
R82099 VDD.n1375 VDD.n1166 4.5005
R82100 VDD.n1318 VDD.n1166 4.5005
R82101 VDD.n1376 VDD.n1166 4.5005
R82102 VDD.n1316 VDD.n1166 4.5005
R82103 VDD.n1377 VDD.n1166 4.5005
R82104 VDD.n1315 VDD.n1166 4.5005
R82105 VDD.n1378 VDD.n1166 4.5005
R82106 VDD.n1313 VDD.n1166 4.5005
R82107 VDD.n1379 VDD.n1166 4.5005
R82108 VDD.n1312 VDD.n1166 4.5005
R82109 VDD.n1380 VDD.n1166 4.5005
R82110 VDD.n1310 VDD.n1166 4.5005
R82111 VDD.n1381 VDD.n1166 4.5005
R82112 VDD.n1309 VDD.n1166 4.5005
R82113 VDD.n1382 VDD.n1166 4.5005
R82114 VDD.n1307 VDD.n1166 4.5005
R82115 VDD.n1383 VDD.n1166 4.5005
R82116 VDD.n1306 VDD.n1166 4.5005
R82117 VDD.n1384 VDD.n1166 4.5005
R82118 VDD.n1304 VDD.n1166 4.5005
R82119 VDD.n1385 VDD.n1166 4.5005
R82120 VDD.n1303 VDD.n1166 4.5005
R82121 VDD.n1386 VDD.n1166 4.5005
R82122 VDD.n1301 VDD.n1166 4.5005
R82123 VDD.n1387 VDD.n1166 4.5005
R82124 VDD.n1300 VDD.n1166 4.5005
R82125 VDD.n1388 VDD.n1166 4.5005
R82126 VDD.n1298 VDD.n1166 4.5005
R82127 VDD.n1389 VDD.n1166 4.5005
R82128 VDD.n1297 VDD.n1166 4.5005
R82129 VDD.n1390 VDD.n1166 4.5005
R82130 VDD.n1295 VDD.n1166 4.5005
R82131 VDD.n1391 VDD.n1166 4.5005
R82132 VDD.n1294 VDD.n1166 4.5005
R82133 VDD.n1392 VDD.n1166 4.5005
R82134 VDD.n1292 VDD.n1166 4.5005
R82135 VDD.n1393 VDD.n1166 4.5005
R82136 VDD.n1291 VDD.n1166 4.5005
R82137 VDD.n1394 VDD.n1166 4.5005
R82138 VDD.n1289 VDD.n1166 4.5005
R82139 VDD.n1395 VDD.n1166 4.5005
R82140 VDD.n1288 VDD.n1166 4.5005
R82141 VDD.n1396 VDD.n1166 4.5005
R82142 VDD.n1286 VDD.n1166 4.5005
R82143 VDD.n1397 VDD.n1166 4.5005
R82144 VDD.n1285 VDD.n1166 4.5005
R82145 VDD.n1398 VDD.n1166 4.5005
R82146 VDD.n1283 VDD.n1166 4.5005
R82147 VDD.n1399 VDD.n1166 4.5005
R82148 VDD.n1282 VDD.n1166 4.5005
R82149 VDD.n1400 VDD.n1166 4.5005
R82150 VDD.n1280 VDD.n1166 4.5005
R82151 VDD.n1401 VDD.n1166 4.5005
R82152 VDD.n1279 VDD.n1166 4.5005
R82153 VDD.n1402 VDD.n1166 4.5005
R82154 VDD.n1277 VDD.n1166 4.5005
R82155 VDD.n1403 VDD.n1166 4.5005
R82156 VDD.n1276 VDD.n1166 4.5005
R82157 VDD.n1404 VDD.n1166 4.5005
R82158 VDD.n1274 VDD.n1166 4.5005
R82159 VDD.n1405 VDD.n1166 4.5005
R82160 VDD.n1273 VDD.n1166 4.5005
R82161 VDD.n1406 VDD.n1166 4.5005
R82162 VDD.n1271 VDD.n1166 4.5005
R82163 VDD.n1407 VDD.n1166 4.5005
R82164 VDD.n1270 VDD.n1166 4.5005
R82165 VDD.n1408 VDD.n1166 4.5005
R82166 VDD.n1268 VDD.n1166 4.5005
R82167 VDD.n1409 VDD.n1166 4.5005
R82168 VDD.n1267 VDD.n1166 4.5005
R82169 VDD.n1410 VDD.n1166 4.5005
R82170 VDD.n1265 VDD.n1166 4.5005
R82171 VDD.n1411 VDD.n1166 4.5005
R82172 VDD.n1264 VDD.n1166 4.5005
R82173 VDD.n1412 VDD.n1166 4.5005
R82174 VDD.n1262 VDD.n1166 4.5005
R82175 VDD.n1413 VDD.n1166 4.5005
R82176 VDD.n1261 VDD.n1166 4.5005
R82177 VDD.n1414 VDD.n1166 4.5005
R82178 VDD.n1415 VDD.n1166 4.5005
R82179 VDD.n1674 VDD.n1166 4.5005
R82180 VDD.n1676 VDD.n1224 4.5005
R82181 VDD.n1341 VDD.n1224 4.5005
R82182 VDD.n1342 VDD.n1224 4.5005
R82183 VDD.n1340 VDD.n1224 4.5005
R82184 VDD.n1344 VDD.n1224 4.5005
R82185 VDD.n1339 VDD.n1224 4.5005
R82186 VDD.n1345 VDD.n1224 4.5005
R82187 VDD.n1338 VDD.n1224 4.5005
R82188 VDD.n1347 VDD.n1224 4.5005
R82189 VDD.n1337 VDD.n1224 4.5005
R82190 VDD.n1348 VDD.n1224 4.5005
R82191 VDD.n1336 VDD.n1224 4.5005
R82192 VDD.n1350 VDD.n1224 4.5005
R82193 VDD.n1335 VDD.n1224 4.5005
R82194 VDD.n1351 VDD.n1224 4.5005
R82195 VDD.n1334 VDD.n1224 4.5005
R82196 VDD.n1353 VDD.n1224 4.5005
R82197 VDD.n1333 VDD.n1224 4.5005
R82198 VDD.n1354 VDD.n1224 4.5005
R82199 VDD.n1332 VDD.n1224 4.5005
R82200 VDD.n1356 VDD.n1224 4.5005
R82201 VDD.n1331 VDD.n1224 4.5005
R82202 VDD.n1357 VDD.n1224 4.5005
R82203 VDD.n1330 VDD.n1224 4.5005
R82204 VDD.n1359 VDD.n1224 4.5005
R82205 VDD.n1329 VDD.n1224 4.5005
R82206 VDD.n1360 VDD.n1224 4.5005
R82207 VDD.n1328 VDD.n1224 4.5005
R82208 VDD.n1362 VDD.n1224 4.5005
R82209 VDD.n1327 VDD.n1224 4.5005
R82210 VDD.n1363 VDD.n1224 4.5005
R82211 VDD.n1326 VDD.n1224 4.5005
R82212 VDD.n1365 VDD.n1224 4.5005
R82213 VDD.n1325 VDD.n1224 4.5005
R82214 VDD.n1366 VDD.n1224 4.5005
R82215 VDD.n1324 VDD.n1224 4.5005
R82216 VDD.n1368 VDD.n1224 4.5005
R82217 VDD.n1323 VDD.n1224 4.5005
R82218 VDD.n1369 VDD.n1224 4.5005
R82219 VDD.n1322 VDD.n1224 4.5005
R82220 VDD.n1371 VDD.n1224 4.5005
R82221 VDD.n1321 VDD.n1224 4.5005
R82222 VDD.n1372 VDD.n1224 4.5005
R82223 VDD.n1320 VDD.n1224 4.5005
R82224 VDD.n1374 VDD.n1224 4.5005
R82225 VDD.n1319 VDD.n1224 4.5005
R82226 VDD.n1375 VDD.n1224 4.5005
R82227 VDD.n1318 VDD.n1224 4.5005
R82228 VDD.n1376 VDD.n1224 4.5005
R82229 VDD.n1316 VDD.n1224 4.5005
R82230 VDD.n1377 VDD.n1224 4.5005
R82231 VDD.n1315 VDD.n1224 4.5005
R82232 VDD.n1378 VDD.n1224 4.5005
R82233 VDD.n1313 VDD.n1224 4.5005
R82234 VDD.n1379 VDD.n1224 4.5005
R82235 VDD.n1312 VDD.n1224 4.5005
R82236 VDD.n1380 VDD.n1224 4.5005
R82237 VDD.n1310 VDD.n1224 4.5005
R82238 VDD.n1381 VDD.n1224 4.5005
R82239 VDD.n1309 VDD.n1224 4.5005
R82240 VDD.n1382 VDD.n1224 4.5005
R82241 VDD.n1307 VDD.n1224 4.5005
R82242 VDD.n1383 VDD.n1224 4.5005
R82243 VDD.n1306 VDD.n1224 4.5005
R82244 VDD.n1384 VDD.n1224 4.5005
R82245 VDD.n1304 VDD.n1224 4.5005
R82246 VDD.n1385 VDD.n1224 4.5005
R82247 VDD.n1303 VDD.n1224 4.5005
R82248 VDD.n1386 VDD.n1224 4.5005
R82249 VDD.n1301 VDD.n1224 4.5005
R82250 VDD.n1387 VDD.n1224 4.5005
R82251 VDD.n1300 VDD.n1224 4.5005
R82252 VDD.n1388 VDD.n1224 4.5005
R82253 VDD.n1298 VDD.n1224 4.5005
R82254 VDD.n1389 VDD.n1224 4.5005
R82255 VDD.n1297 VDD.n1224 4.5005
R82256 VDD.n1390 VDD.n1224 4.5005
R82257 VDD.n1295 VDD.n1224 4.5005
R82258 VDD.n1391 VDD.n1224 4.5005
R82259 VDD.n1294 VDD.n1224 4.5005
R82260 VDD.n1392 VDD.n1224 4.5005
R82261 VDD.n1292 VDD.n1224 4.5005
R82262 VDD.n1393 VDD.n1224 4.5005
R82263 VDD.n1291 VDD.n1224 4.5005
R82264 VDD.n1394 VDD.n1224 4.5005
R82265 VDD.n1289 VDD.n1224 4.5005
R82266 VDD.n1395 VDD.n1224 4.5005
R82267 VDD.n1288 VDD.n1224 4.5005
R82268 VDD.n1396 VDD.n1224 4.5005
R82269 VDD.n1286 VDD.n1224 4.5005
R82270 VDD.n1397 VDD.n1224 4.5005
R82271 VDD.n1285 VDD.n1224 4.5005
R82272 VDD.n1398 VDD.n1224 4.5005
R82273 VDD.n1283 VDD.n1224 4.5005
R82274 VDD.n1399 VDD.n1224 4.5005
R82275 VDD.n1282 VDD.n1224 4.5005
R82276 VDD.n1400 VDD.n1224 4.5005
R82277 VDD.n1280 VDD.n1224 4.5005
R82278 VDD.n1401 VDD.n1224 4.5005
R82279 VDD.n1279 VDD.n1224 4.5005
R82280 VDD.n1402 VDD.n1224 4.5005
R82281 VDD.n1277 VDD.n1224 4.5005
R82282 VDD.n1403 VDD.n1224 4.5005
R82283 VDD.n1276 VDD.n1224 4.5005
R82284 VDD.n1404 VDD.n1224 4.5005
R82285 VDD.n1274 VDD.n1224 4.5005
R82286 VDD.n1405 VDD.n1224 4.5005
R82287 VDD.n1273 VDD.n1224 4.5005
R82288 VDD.n1406 VDD.n1224 4.5005
R82289 VDD.n1271 VDD.n1224 4.5005
R82290 VDD.n1407 VDD.n1224 4.5005
R82291 VDD.n1270 VDD.n1224 4.5005
R82292 VDD.n1408 VDD.n1224 4.5005
R82293 VDD.n1268 VDD.n1224 4.5005
R82294 VDD.n1409 VDD.n1224 4.5005
R82295 VDD.n1267 VDD.n1224 4.5005
R82296 VDD.n1410 VDD.n1224 4.5005
R82297 VDD.n1265 VDD.n1224 4.5005
R82298 VDD.n1411 VDD.n1224 4.5005
R82299 VDD.n1264 VDD.n1224 4.5005
R82300 VDD.n1412 VDD.n1224 4.5005
R82301 VDD.n1262 VDD.n1224 4.5005
R82302 VDD.n1413 VDD.n1224 4.5005
R82303 VDD.n1261 VDD.n1224 4.5005
R82304 VDD.n1414 VDD.n1224 4.5005
R82305 VDD.n1415 VDD.n1224 4.5005
R82306 VDD.n1674 VDD.n1224 4.5005
R82307 VDD.n1676 VDD.n1165 4.5005
R82308 VDD.n1341 VDD.n1165 4.5005
R82309 VDD.n1342 VDD.n1165 4.5005
R82310 VDD.n1340 VDD.n1165 4.5005
R82311 VDD.n1344 VDD.n1165 4.5005
R82312 VDD.n1339 VDD.n1165 4.5005
R82313 VDD.n1345 VDD.n1165 4.5005
R82314 VDD.n1338 VDD.n1165 4.5005
R82315 VDD.n1347 VDD.n1165 4.5005
R82316 VDD.n1337 VDD.n1165 4.5005
R82317 VDD.n1348 VDD.n1165 4.5005
R82318 VDD.n1336 VDD.n1165 4.5005
R82319 VDD.n1350 VDD.n1165 4.5005
R82320 VDD.n1335 VDD.n1165 4.5005
R82321 VDD.n1351 VDD.n1165 4.5005
R82322 VDD.n1334 VDD.n1165 4.5005
R82323 VDD.n1353 VDD.n1165 4.5005
R82324 VDD.n1333 VDD.n1165 4.5005
R82325 VDD.n1354 VDD.n1165 4.5005
R82326 VDD.n1332 VDD.n1165 4.5005
R82327 VDD.n1356 VDD.n1165 4.5005
R82328 VDD.n1331 VDD.n1165 4.5005
R82329 VDD.n1357 VDD.n1165 4.5005
R82330 VDD.n1330 VDD.n1165 4.5005
R82331 VDD.n1359 VDD.n1165 4.5005
R82332 VDD.n1329 VDD.n1165 4.5005
R82333 VDD.n1360 VDD.n1165 4.5005
R82334 VDD.n1328 VDD.n1165 4.5005
R82335 VDD.n1362 VDD.n1165 4.5005
R82336 VDD.n1327 VDD.n1165 4.5005
R82337 VDD.n1363 VDD.n1165 4.5005
R82338 VDD.n1326 VDD.n1165 4.5005
R82339 VDD.n1365 VDD.n1165 4.5005
R82340 VDD.n1325 VDD.n1165 4.5005
R82341 VDD.n1366 VDD.n1165 4.5005
R82342 VDD.n1324 VDD.n1165 4.5005
R82343 VDD.n1368 VDD.n1165 4.5005
R82344 VDD.n1323 VDD.n1165 4.5005
R82345 VDD.n1369 VDD.n1165 4.5005
R82346 VDD.n1322 VDD.n1165 4.5005
R82347 VDD.n1371 VDD.n1165 4.5005
R82348 VDD.n1321 VDD.n1165 4.5005
R82349 VDD.n1372 VDD.n1165 4.5005
R82350 VDD.n1320 VDD.n1165 4.5005
R82351 VDD.n1374 VDD.n1165 4.5005
R82352 VDD.n1319 VDD.n1165 4.5005
R82353 VDD.n1375 VDD.n1165 4.5005
R82354 VDD.n1318 VDD.n1165 4.5005
R82355 VDD.n1376 VDD.n1165 4.5005
R82356 VDD.n1316 VDD.n1165 4.5005
R82357 VDD.n1377 VDD.n1165 4.5005
R82358 VDD.n1315 VDD.n1165 4.5005
R82359 VDD.n1378 VDD.n1165 4.5005
R82360 VDD.n1313 VDD.n1165 4.5005
R82361 VDD.n1379 VDD.n1165 4.5005
R82362 VDD.n1312 VDD.n1165 4.5005
R82363 VDD.n1380 VDD.n1165 4.5005
R82364 VDD.n1310 VDD.n1165 4.5005
R82365 VDD.n1381 VDD.n1165 4.5005
R82366 VDD.n1309 VDD.n1165 4.5005
R82367 VDD.n1382 VDD.n1165 4.5005
R82368 VDD.n1307 VDD.n1165 4.5005
R82369 VDD.n1383 VDD.n1165 4.5005
R82370 VDD.n1306 VDD.n1165 4.5005
R82371 VDD.n1384 VDD.n1165 4.5005
R82372 VDD.n1304 VDD.n1165 4.5005
R82373 VDD.n1385 VDD.n1165 4.5005
R82374 VDD.n1303 VDD.n1165 4.5005
R82375 VDD.n1386 VDD.n1165 4.5005
R82376 VDD.n1301 VDD.n1165 4.5005
R82377 VDD.n1387 VDD.n1165 4.5005
R82378 VDD.n1300 VDD.n1165 4.5005
R82379 VDD.n1388 VDD.n1165 4.5005
R82380 VDD.n1298 VDD.n1165 4.5005
R82381 VDD.n1389 VDD.n1165 4.5005
R82382 VDD.n1297 VDD.n1165 4.5005
R82383 VDD.n1390 VDD.n1165 4.5005
R82384 VDD.n1295 VDD.n1165 4.5005
R82385 VDD.n1391 VDD.n1165 4.5005
R82386 VDD.n1294 VDD.n1165 4.5005
R82387 VDD.n1392 VDD.n1165 4.5005
R82388 VDD.n1292 VDD.n1165 4.5005
R82389 VDD.n1393 VDD.n1165 4.5005
R82390 VDD.n1291 VDD.n1165 4.5005
R82391 VDD.n1394 VDD.n1165 4.5005
R82392 VDD.n1289 VDD.n1165 4.5005
R82393 VDD.n1395 VDD.n1165 4.5005
R82394 VDD.n1288 VDD.n1165 4.5005
R82395 VDD.n1396 VDD.n1165 4.5005
R82396 VDD.n1286 VDD.n1165 4.5005
R82397 VDD.n1397 VDD.n1165 4.5005
R82398 VDD.n1285 VDD.n1165 4.5005
R82399 VDD.n1398 VDD.n1165 4.5005
R82400 VDD.n1283 VDD.n1165 4.5005
R82401 VDD.n1399 VDD.n1165 4.5005
R82402 VDD.n1282 VDD.n1165 4.5005
R82403 VDD.n1400 VDD.n1165 4.5005
R82404 VDD.n1280 VDD.n1165 4.5005
R82405 VDD.n1401 VDD.n1165 4.5005
R82406 VDD.n1279 VDD.n1165 4.5005
R82407 VDD.n1402 VDD.n1165 4.5005
R82408 VDD.n1277 VDD.n1165 4.5005
R82409 VDD.n1403 VDD.n1165 4.5005
R82410 VDD.n1276 VDD.n1165 4.5005
R82411 VDD.n1404 VDD.n1165 4.5005
R82412 VDD.n1274 VDD.n1165 4.5005
R82413 VDD.n1405 VDD.n1165 4.5005
R82414 VDD.n1273 VDD.n1165 4.5005
R82415 VDD.n1406 VDD.n1165 4.5005
R82416 VDD.n1271 VDD.n1165 4.5005
R82417 VDD.n1407 VDD.n1165 4.5005
R82418 VDD.n1270 VDD.n1165 4.5005
R82419 VDD.n1408 VDD.n1165 4.5005
R82420 VDD.n1268 VDD.n1165 4.5005
R82421 VDD.n1409 VDD.n1165 4.5005
R82422 VDD.n1267 VDD.n1165 4.5005
R82423 VDD.n1410 VDD.n1165 4.5005
R82424 VDD.n1265 VDD.n1165 4.5005
R82425 VDD.n1411 VDD.n1165 4.5005
R82426 VDD.n1264 VDD.n1165 4.5005
R82427 VDD.n1412 VDD.n1165 4.5005
R82428 VDD.n1262 VDD.n1165 4.5005
R82429 VDD.n1413 VDD.n1165 4.5005
R82430 VDD.n1261 VDD.n1165 4.5005
R82431 VDD.n1414 VDD.n1165 4.5005
R82432 VDD.n1415 VDD.n1165 4.5005
R82433 VDD.n1674 VDD.n1165 4.5005
R82434 VDD.n1676 VDD.n1225 4.5005
R82435 VDD.n1341 VDD.n1225 4.5005
R82436 VDD.n1342 VDD.n1225 4.5005
R82437 VDD.n1340 VDD.n1225 4.5005
R82438 VDD.n1344 VDD.n1225 4.5005
R82439 VDD.n1339 VDD.n1225 4.5005
R82440 VDD.n1345 VDD.n1225 4.5005
R82441 VDD.n1338 VDD.n1225 4.5005
R82442 VDD.n1347 VDD.n1225 4.5005
R82443 VDD.n1337 VDD.n1225 4.5005
R82444 VDD.n1348 VDD.n1225 4.5005
R82445 VDD.n1336 VDD.n1225 4.5005
R82446 VDD.n1350 VDD.n1225 4.5005
R82447 VDD.n1335 VDD.n1225 4.5005
R82448 VDD.n1351 VDD.n1225 4.5005
R82449 VDD.n1334 VDD.n1225 4.5005
R82450 VDD.n1353 VDD.n1225 4.5005
R82451 VDD.n1333 VDD.n1225 4.5005
R82452 VDD.n1354 VDD.n1225 4.5005
R82453 VDD.n1332 VDD.n1225 4.5005
R82454 VDD.n1356 VDD.n1225 4.5005
R82455 VDD.n1331 VDD.n1225 4.5005
R82456 VDD.n1357 VDD.n1225 4.5005
R82457 VDD.n1330 VDD.n1225 4.5005
R82458 VDD.n1359 VDD.n1225 4.5005
R82459 VDD.n1329 VDD.n1225 4.5005
R82460 VDD.n1360 VDD.n1225 4.5005
R82461 VDD.n1328 VDD.n1225 4.5005
R82462 VDD.n1362 VDD.n1225 4.5005
R82463 VDD.n1327 VDD.n1225 4.5005
R82464 VDD.n1363 VDD.n1225 4.5005
R82465 VDD.n1326 VDD.n1225 4.5005
R82466 VDD.n1365 VDD.n1225 4.5005
R82467 VDD.n1325 VDD.n1225 4.5005
R82468 VDD.n1366 VDD.n1225 4.5005
R82469 VDD.n1324 VDD.n1225 4.5005
R82470 VDD.n1368 VDD.n1225 4.5005
R82471 VDD.n1323 VDD.n1225 4.5005
R82472 VDD.n1369 VDD.n1225 4.5005
R82473 VDD.n1322 VDD.n1225 4.5005
R82474 VDD.n1371 VDD.n1225 4.5005
R82475 VDD.n1321 VDD.n1225 4.5005
R82476 VDD.n1372 VDD.n1225 4.5005
R82477 VDD.n1320 VDD.n1225 4.5005
R82478 VDD.n1374 VDD.n1225 4.5005
R82479 VDD.n1319 VDD.n1225 4.5005
R82480 VDD.n1375 VDD.n1225 4.5005
R82481 VDD.n1318 VDD.n1225 4.5005
R82482 VDD.n1376 VDD.n1225 4.5005
R82483 VDD.n1316 VDD.n1225 4.5005
R82484 VDD.n1377 VDD.n1225 4.5005
R82485 VDD.n1315 VDD.n1225 4.5005
R82486 VDD.n1378 VDD.n1225 4.5005
R82487 VDD.n1313 VDD.n1225 4.5005
R82488 VDD.n1379 VDD.n1225 4.5005
R82489 VDD.n1312 VDD.n1225 4.5005
R82490 VDD.n1380 VDD.n1225 4.5005
R82491 VDD.n1310 VDD.n1225 4.5005
R82492 VDD.n1381 VDD.n1225 4.5005
R82493 VDD.n1309 VDD.n1225 4.5005
R82494 VDD.n1382 VDD.n1225 4.5005
R82495 VDD.n1307 VDD.n1225 4.5005
R82496 VDD.n1383 VDD.n1225 4.5005
R82497 VDD.n1306 VDD.n1225 4.5005
R82498 VDD.n1384 VDD.n1225 4.5005
R82499 VDD.n1304 VDD.n1225 4.5005
R82500 VDD.n1385 VDD.n1225 4.5005
R82501 VDD.n1303 VDD.n1225 4.5005
R82502 VDD.n1386 VDD.n1225 4.5005
R82503 VDD.n1301 VDD.n1225 4.5005
R82504 VDD.n1387 VDD.n1225 4.5005
R82505 VDD.n1300 VDD.n1225 4.5005
R82506 VDD.n1388 VDD.n1225 4.5005
R82507 VDD.n1298 VDD.n1225 4.5005
R82508 VDD.n1389 VDD.n1225 4.5005
R82509 VDD.n1297 VDD.n1225 4.5005
R82510 VDD.n1390 VDD.n1225 4.5005
R82511 VDD.n1295 VDD.n1225 4.5005
R82512 VDD.n1391 VDD.n1225 4.5005
R82513 VDD.n1294 VDD.n1225 4.5005
R82514 VDD.n1392 VDD.n1225 4.5005
R82515 VDD.n1292 VDD.n1225 4.5005
R82516 VDD.n1393 VDD.n1225 4.5005
R82517 VDD.n1291 VDD.n1225 4.5005
R82518 VDD.n1394 VDD.n1225 4.5005
R82519 VDD.n1289 VDD.n1225 4.5005
R82520 VDD.n1395 VDD.n1225 4.5005
R82521 VDD.n1288 VDD.n1225 4.5005
R82522 VDD.n1396 VDD.n1225 4.5005
R82523 VDD.n1286 VDD.n1225 4.5005
R82524 VDD.n1397 VDD.n1225 4.5005
R82525 VDD.n1285 VDD.n1225 4.5005
R82526 VDD.n1398 VDD.n1225 4.5005
R82527 VDD.n1283 VDD.n1225 4.5005
R82528 VDD.n1399 VDD.n1225 4.5005
R82529 VDD.n1282 VDD.n1225 4.5005
R82530 VDD.n1400 VDD.n1225 4.5005
R82531 VDD.n1280 VDD.n1225 4.5005
R82532 VDD.n1401 VDD.n1225 4.5005
R82533 VDD.n1279 VDD.n1225 4.5005
R82534 VDD.n1402 VDD.n1225 4.5005
R82535 VDD.n1277 VDD.n1225 4.5005
R82536 VDD.n1403 VDD.n1225 4.5005
R82537 VDD.n1276 VDD.n1225 4.5005
R82538 VDD.n1404 VDD.n1225 4.5005
R82539 VDD.n1274 VDD.n1225 4.5005
R82540 VDD.n1405 VDD.n1225 4.5005
R82541 VDD.n1273 VDD.n1225 4.5005
R82542 VDD.n1406 VDD.n1225 4.5005
R82543 VDD.n1271 VDD.n1225 4.5005
R82544 VDD.n1407 VDD.n1225 4.5005
R82545 VDD.n1270 VDD.n1225 4.5005
R82546 VDD.n1408 VDD.n1225 4.5005
R82547 VDD.n1268 VDD.n1225 4.5005
R82548 VDD.n1409 VDD.n1225 4.5005
R82549 VDD.n1267 VDD.n1225 4.5005
R82550 VDD.n1410 VDD.n1225 4.5005
R82551 VDD.n1265 VDD.n1225 4.5005
R82552 VDD.n1411 VDD.n1225 4.5005
R82553 VDD.n1264 VDD.n1225 4.5005
R82554 VDD.n1412 VDD.n1225 4.5005
R82555 VDD.n1262 VDD.n1225 4.5005
R82556 VDD.n1413 VDD.n1225 4.5005
R82557 VDD.n1261 VDD.n1225 4.5005
R82558 VDD.n1414 VDD.n1225 4.5005
R82559 VDD.n1415 VDD.n1225 4.5005
R82560 VDD.n1674 VDD.n1225 4.5005
R82561 VDD.n1676 VDD.n1164 4.5005
R82562 VDD.n1341 VDD.n1164 4.5005
R82563 VDD.n1342 VDD.n1164 4.5005
R82564 VDD.n1340 VDD.n1164 4.5005
R82565 VDD.n1344 VDD.n1164 4.5005
R82566 VDD.n1339 VDD.n1164 4.5005
R82567 VDD.n1345 VDD.n1164 4.5005
R82568 VDD.n1338 VDD.n1164 4.5005
R82569 VDD.n1347 VDD.n1164 4.5005
R82570 VDD.n1337 VDD.n1164 4.5005
R82571 VDD.n1348 VDD.n1164 4.5005
R82572 VDD.n1336 VDD.n1164 4.5005
R82573 VDD.n1350 VDD.n1164 4.5005
R82574 VDD.n1335 VDD.n1164 4.5005
R82575 VDD.n1351 VDD.n1164 4.5005
R82576 VDD.n1334 VDD.n1164 4.5005
R82577 VDD.n1353 VDD.n1164 4.5005
R82578 VDD.n1333 VDD.n1164 4.5005
R82579 VDD.n1354 VDD.n1164 4.5005
R82580 VDD.n1332 VDD.n1164 4.5005
R82581 VDD.n1356 VDD.n1164 4.5005
R82582 VDD.n1331 VDD.n1164 4.5005
R82583 VDD.n1357 VDD.n1164 4.5005
R82584 VDD.n1330 VDD.n1164 4.5005
R82585 VDD.n1359 VDD.n1164 4.5005
R82586 VDD.n1329 VDD.n1164 4.5005
R82587 VDD.n1360 VDD.n1164 4.5005
R82588 VDD.n1328 VDD.n1164 4.5005
R82589 VDD.n1362 VDD.n1164 4.5005
R82590 VDD.n1327 VDD.n1164 4.5005
R82591 VDD.n1363 VDD.n1164 4.5005
R82592 VDD.n1326 VDD.n1164 4.5005
R82593 VDD.n1365 VDD.n1164 4.5005
R82594 VDD.n1325 VDD.n1164 4.5005
R82595 VDD.n1366 VDD.n1164 4.5005
R82596 VDD.n1324 VDD.n1164 4.5005
R82597 VDD.n1368 VDD.n1164 4.5005
R82598 VDD.n1323 VDD.n1164 4.5005
R82599 VDD.n1369 VDD.n1164 4.5005
R82600 VDD.n1322 VDD.n1164 4.5005
R82601 VDD.n1371 VDD.n1164 4.5005
R82602 VDD.n1321 VDD.n1164 4.5005
R82603 VDD.n1372 VDD.n1164 4.5005
R82604 VDD.n1320 VDD.n1164 4.5005
R82605 VDD.n1374 VDD.n1164 4.5005
R82606 VDD.n1319 VDD.n1164 4.5005
R82607 VDD.n1375 VDD.n1164 4.5005
R82608 VDD.n1318 VDD.n1164 4.5005
R82609 VDD.n1376 VDD.n1164 4.5005
R82610 VDD.n1316 VDD.n1164 4.5005
R82611 VDD.n1377 VDD.n1164 4.5005
R82612 VDD.n1315 VDD.n1164 4.5005
R82613 VDD.n1378 VDD.n1164 4.5005
R82614 VDD.n1313 VDD.n1164 4.5005
R82615 VDD.n1379 VDD.n1164 4.5005
R82616 VDD.n1312 VDD.n1164 4.5005
R82617 VDD.n1380 VDD.n1164 4.5005
R82618 VDD.n1310 VDD.n1164 4.5005
R82619 VDD.n1381 VDD.n1164 4.5005
R82620 VDD.n1309 VDD.n1164 4.5005
R82621 VDD.n1382 VDD.n1164 4.5005
R82622 VDD.n1307 VDD.n1164 4.5005
R82623 VDD.n1383 VDD.n1164 4.5005
R82624 VDD.n1306 VDD.n1164 4.5005
R82625 VDD.n1384 VDD.n1164 4.5005
R82626 VDD.n1304 VDD.n1164 4.5005
R82627 VDD.n1385 VDD.n1164 4.5005
R82628 VDD.n1303 VDD.n1164 4.5005
R82629 VDD.n1386 VDD.n1164 4.5005
R82630 VDD.n1301 VDD.n1164 4.5005
R82631 VDD.n1387 VDD.n1164 4.5005
R82632 VDD.n1300 VDD.n1164 4.5005
R82633 VDD.n1388 VDD.n1164 4.5005
R82634 VDD.n1298 VDD.n1164 4.5005
R82635 VDD.n1389 VDD.n1164 4.5005
R82636 VDD.n1297 VDD.n1164 4.5005
R82637 VDD.n1390 VDD.n1164 4.5005
R82638 VDD.n1295 VDD.n1164 4.5005
R82639 VDD.n1391 VDD.n1164 4.5005
R82640 VDD.n1294 VDD.n1164 4.5005
R82641 VDD.n1392 VDD.n1164 4.5005
R82642 VDD.n1292 VDD.n1164 4.5005
R82643 VDD.n1393 VDD.n1164 4.5005
R82644 VDD.n1291 VDD.n1164 4.5005
R82645 VDD.n1394 VDD.n1164 4.5005
R82646 VDD.n1289 VDD.n1164 4.5005
R82647 VDD.n1395 VDD.n1164 4.5005
R82648 VDD.n1288 VDD.n1164 4.5005
R82649 VDD.n1396 VDD.n1164 4.5005
R82650 VDD.n1286 VDD.n1164 4.5005
R82651 VDD.n1397 VDD.n1164 4.5005
R82652 VDD.n1285 VDD.n1164 4.5005
R82653 VDD.n1398 VDD.n1164 4.5005
R82654 VDD.n1283 VDD.n1164 4.5005
R82655 VDD.n1399 VDD.n1164 4.5005
R82656 VDD.n1282 VDD.n1164 4.5005
R82657 VDD.n1400 VDD.n1164 4.5005
R82658 VDD.n1280 VDD.n1164 4.5005
R82659 VDD.n1401 VDD.n1164 4.5005
R82660 VDD.n1279 VDD.n1164 4.5005
R82661 VDD.n1402 VDD.n1164 4.5005
R82662 VDD.n1277 VDD.n1164 4.5005
R82663 VDD.n1403 VDD.n1164 4.5005
R82664 VDD.n1276 VDD.n1164 4.5005
R82665 VDD.n1404 VDD.n1164 4.5005
R82666 VDD.n1274 VDD.n1164 4.5005
R82667 VDD.n1405 VDD.n1164 4.5005
R82668 VDD.n1273 VDD.n1164 4.5005
R82669 VDD.n1406 VDD.n1164 4.5005
R82670 VDD.n1271 VDD.n1164 4.5005
R82671 VDD.n1407 VDD.n1164 4.5005
R82672 VDD.n1270 VDD.n1164 4.5005
R82673 VDD.n1408 VDD.n1164 4.5005
R82674 VDD.n1268 VDD.n1164 4.5005
R82675 VDD.n1409 VDD.n1164 4.5005
R82676 VDD.n1267 VDD.n1164 4.5005
R82677 VDD.n1410 VDD.n1164 4.5005
R82678 VDD.n1265 VDD.n1164 4.5005
R82679 VDD.n1411 VDD.n1164 4.5005
R82680 VDD.n1264 VDD.n1164 4.5005
R82681 VDD.n1412 VDD.n1164 4.5005
R82682 VDD.n1262 VDD.n1164 4.5005
R82683 VDD.n1413 VDD.n1164 4.5005
R82684 VDD.n1261 VDD.n1164 4.5005
R82685 VDD.n1414 VDD.n1164 4.5005
R82686 VDD.n1415 VDD.n1164 4.5005
R82687 VDD.n1674 VDD.n1164 4.5005
R82688 VDD.n1676 VDD.n1226 4.5005
R82689 VDD.n1341 VDD.n1226 4.5005
R82690 VDD.n1342 VDD.n1226 4.5005
R82691 VDD.n1340 VDD.n1226 4.5005
R82692 VDD.n1344 VDD.n1226 4.5005
R82693 VDD.n1339 VDD.n1226 4.5005
R82694 VDD.n1345 VDD.n1226 4.5005
R82695 VDD.n1338 VDD.n1226 4.5005
R82696 VDD.n1347 VDD.n1226 4.5005
R82697 VDD.n1337 VDD.n1226 4.5005
R82698 VDD.n1348 VDD.n1226 4.5005
R82699 VDD.n1336 VDD.n1226 4.5005
R82700 VDD.n1350 VDD.n1226 4.5005
R82701 VDD.n1335 VDD.n1226 4.5005
R82702 VDD.n1351 VDD.n1226 4.5005
R82703 VDD.n1334 VDD.n1226 4.5005
R82704 VDD.n1353 VDD.n1226 4.5005
R82705 VDD.n1333 VDD.n1226 4.5005
R82706 VDD.n1354 VDD.n1226 4.5005
R82707 VDD.n1332 VDD.n1226 4.5005
R82708 VDD.n1356 VDD.n1226 4.5005
R82709 VDD.n1331 VDD.n1226 4.5005
R82710 VDD.n1357 VDD.n1226 4.5005
R82711 VDD.n1330 VDD.n1226 4.5005
R82712 VDD.n1359 VDD.n1226 4.5005
R82713 VDD.n1329 VDD.n1226 4.5005
R82714 VDD.n1360 VDD.n1226 4.5005
R82715 VDD.n1328 VDD.n1226 4.5005
R82716 VDD.n1362 VDD.n1226 4.5005
R82717 VDD.n1327 VDD.n1226 4.5005
R82718 VDD.n1363 VDD.n1226 4.5005
R82719 VDD.n1326 VDD.n1226 4.5005
R82720 VDD.n1365 VDD.n1226 4.5005
R82721 VDD.n1325 VDD.n1226 4.5005
R82722 VDD.n1366 VDD.n1226 4.5005
R82723 VDD.n1324 VDD.n1226 4.5005
R82724 VDD.n1368 VDD.n1226 4.5005
R82725 VDD.n1323 VDD.n1226 4.5005
R82726 VDD.n1369 VDD.n1226 4.5005
R82727 VDD.n1322 VDD.n1226 4.5005
R82728 VDD.n1371 VDD.n1226 4.5005
R82729 VDD.n1321 VDD.n1226 4.5005
R82730 VDD.n1372 VDD.n1226 4.5005
R82731 VDD.n1320 VDD.n1226 4.5005
R82732 VDD.n1374 VDD.n1226 4.5005
R82733 VDD.n1319 VDD.n1226 4.5005
R82734 VDD.n1375 VDD.n1226 4.5005
R82735 VDD.n1318 VDD.n1226 4.5005
R82736 VDD.n1376 VDD.n1226 4.5005
R82737 VDD.n1316 VDD.n1226 4.5005
R82738 VDD.n1377 VDD.n1226 4.5005
R82739 VDD.n1315 VDD.n1226 4.5005
R82740 VDD.n1378 VDD.n1226 4.5005
R82741 VDD.n1313 VDD.n1226 4.5005
R82742 VDD.n1379 VDD.n1226 4.5005
R82743 VDD.n1312 VDD.n1226 4.5005
R82744 VDD.n1380 VDD.n1226 4.5005
R82745 VDD.n1310 VDD.n1226 4.5005
R82746 VDD.n1381 VDD.n1226 4.5005
R82747 VDD.n1309 VDD.n1226 4.5005
R82748 VDD.n1382 VDD.n1226 4.5005
R82749 VDD.n1307 VDD.n1226 4.5005
R82750 VDD.n1383 VDD.n1226 4.5005
R82751 VDD.n1306 VDD.n1226 4.5005
R82752 VDD.n1384 VDD.n1226 4.5005
R82753 VDD.n1304 VDD.n1226 4.5005
R82754 VDD.n1385 VDD.n1226 4.5005
R82755 VDD.n1303 VDD.n1226 4.5005
R82756 VDD.n1386 VDD.n1226 4.5005
R82757 VDD.n1301 VDD.n1226 4.5005
R82758 VDD.n1387 VDD.n1226 4.5005
R82759 VDD.n1300 VDD.n1226 4.5005
R82760 VDD.n1388 VDD.n1226 4.5005
R82761 VDD.n1298 VDD.n1226 4.5005
R82762 VDD.n1389 VDD.n1226 4.5005
R82763 VDD.n1297 VDD.n1226 4.5005
R82764 VDD.n1390 VDD.n1226 4.5005
R82765 VDD.n1295 VDD.n1226 4.5005
R82766 VDD.n1391 VDD.n1226 4.5005
R82767 VDD.n1294 VDD.n1226 4.5005
R82768 VDD.n1392 VDD.n1226 4.5005
R82769 VDD.n1292 VDD.n1226 4.5005
R82770 VDD.n1393 VDD.n1226 4.5005
R82771 VDD.n1291 VDD.n1226 4.5005
R82772 VDD.n1394 VDD.n1226 4.5005
R82773 VDD.n1289 VDD.n1226 4.5005
R82774 VDD.n1395 VDD.n1226 4.5005
R82775 VDD.n1288 VDD.n1226 4.5005
R82776 VDD.n1396 VDD.n1226 4.5005
R82777 VDD.n1286 VDD.n1226 4.5005
R82778 VDD.n1397 VDD.n1226 4.5005
R82779 VDD.n1285 VDD.n1226 4.5005
R82780 VDD.n1398 VDD.n1226 4.5005
R82781 VDD.n1283 VDD.n1226 4.5005
R82782 VDD.n1399 VDD.n1226 4.5005
R82783 VDD.n1282 VDD.n1226 4.5005
R82784 VDD.n1400 VDD.n1226 4.5005
R82785 VDD.n1280 VDD.n1226 4.5005
R82786 VDD.n1401 VDD.n1226 4.5005
R82787 VDD.n1279 VDD.n1226 4.5005
R82788 VDD.n1402 VDD.n1226 4.5005
R82789 VDD.n1277 VDD.n1226 4.5005
R82790 VDD.n1403 VDD.n1226 4.5005
R82791 VDD.n1276 VDD.n1226 4.5005
R82792 VDD.n1404 VDD.n1226 4.5005
R82793 VDD.n1274 VDD.n1226 4.5005
R82794 VDD.n1405 VDD.n1226 4.5005
R82795 VDD.n1273 VDD.n1226 4.5005
R82796 VDD.n1406 VDD.n1226 4.5005
R82797 VDD.n1271 VDD.n1226 4.5005
R82798 VDD.n1407 VDD.n1226 4.5005
R82799 VDD.n1270 VDD.n1226 4.5005
R82800 VDD.n1408 VDD.n1226 4.5005
R82801 VDD.n1268 VDD.n1226 4.5005
R82802 VDD.n1409 VDD.n1226 4.5005
R82803 VDD.n1267 VDD.n1226 4.5005
R82804 VDD.n1410 VDD.n1226 4.5005
R82805 VDD.n1265 VDD.n1226 4.5005
R82806 VDD.n1411 VDD.n1226 4.5005
R82807 VDD.n1264 VDD.n1226 4.5005
R82808 VDD.n1412 VDD.n1226 4.5005
R82809 VDD.n1262 VDD.n1226 4.5005
R82810 VDD.n1413 VDD.n1226 4.5005
R82811 VDD.n1261 VDD.n1226 4.5005
R82812 VDD.n1414 VDD.n1226 4.5005
R82813 VDD.n1415 VDD.n1226 4.5005
R82814 VDD.n1674 VDD.n1226 4.5005
R82815 VDD.n1676 VDD.n1163 4.5005
R82816 VDD.n1341 VDD.n1163 4.5005
R82817 VDD.n1342 VDD.n1163 4.5005
R82818 VDD.n1340 VDD.n1163 4.5005
R82819 VDD.n1344 VDD.n1163 4.5005
R82820 VDD.n1339 VDD.n1163 4.5005
R82821 VDD.n1345 VDD.n1163 4.5005
R82822 VDD.n1338 VDD.n1163 4.5005
R82823 VDD.n1347 VDD.n1163 4.5005
R82824 VDD.n1337 VDD.n1163 4.5005
R82825 VDD.n1348 VDD.n1163 4.5005
R82826 VDD.n1336 VDD.n1163 4.5005
R82827 VDD.n1350 VDD.n1163 4.5005
R82828 VDD.n1335 VDD.n1163 4.5005
R82829 VDD.n1351 VDD.n1163 4.5005
R82830 VDD.n1334 VDD.n1163 4.5005
R82831 VDD.n1353 VDD.n1163 4.5005
R82832 VDD.n1333 VDD.n1163 4.5005
R82833 VDD.n1354 VDD.n1163 4.5005
R82834 VDD.n1332 VDD.n1163 4.5005
R82835 VDD.n1356 VDD.n1163 4.5005
R82836 VDD.n1331 VDD.n1163 4.5005
R82837 VDD.n1357 VDD.n1163 4.5005
R82838 VDD.n1330 VDD.n1163 4.5005
R82839 VDD.n1359 VDD.n1163 4.5005
R82840 VDD.n1329 VDD.n1163 4.5005
R82841 VDD.n1360 VDD.n1163 4.5005
R82842 VDD.n1328 VDD.n1163 4.5005
R82843 VDD.n1362 VDD.n1163 4.5005
R82844 VDD.n1327 VDD.n1163 4.5005
R82845 VDD.n1363 VDD.n1163 4.5005
R82846 VDD.n1326 VDD.n1163 4.5005
R82847 VDD.n1365 VDD.n1163 4.5005
R82848 VDD.n1325 VDD.n1163 4.5005
R82849 VDD.n1366 VDD.n1163 4.5005
R82850 VDD.n1324 VDD.n1163 4.5005
R82851 VDD.n1368 VDD.n1163 4.5005
R82852 VDD.n1323 VDD.n1163 4.5005
R82853 VDD.n1369 VDD.n1163 4.5005
R82854 VDD.n1322 VDD.n1163 4.5005
R82855 VDD.n1371 VDD.n1163 4.5005
R82856 VDD.n1321 VDD.n1163 4.5005
R82857 VDD.n1372 VDD.n1163 4.5005
R82858 VDD.n1320 VDD.n1163 4.5005
R82859 VDD.n1374 VDD.n1163 4.5005
R82860 VDD.n1319 VDD.n1163 4.5005
R82861 VDD.n1375 VDD.n1163 4.5005
R82862 VDD.n1318 VDD.n1163 4.5005
R82863 VDD.n1376 VDD.n1163 4.5005
R82864 VDD.n1316 VDD.n1163 4.5005
R82865 VDD.n1377 VDD.n1163 4.5005
R82866 VDD.n1315 VDD.n1163 4.5005
R82867 VDD.n1378 VDD.n1163 4.5005
R82868 VDD.n1313 VDD.n1163 4.5005
R82869 VDD.n1379 VDD.n1163 4.5005
R82870 VDD.n1312 VDD.n1163 4.5005
R82871 VDD.n1380 VDD.n1163 4.5005
R82872 VDD.n1310 VDD.n1163 4.5005
R82873 VDD.n1381 VDD.n1163 4.5005
R82874 VDD.n1309 VDD.n1163 4.5005
R82875 VDD.n1382 VDD.n1163 4.5005
R82876 VDD.n1307 VDD.n1163 4.5005
R82877 VDD.n1383 VDD.n1163 4.5005
R82878 VDD.n1306 VDD.n1163 4.5005
R82879 VDD.n1384 VDD.n1163 4.5005
R82880 VDD.n1304 VDD.n1163 4.5005
R82881 VDD.n1385 VDD.n1163 4.5005
R82882 VDD.n1303 VDD.n1163 4.5005
R82883 VDD.n1386 VDD.n1163 4.5005
R82884 VDD.n1301 VDD.n1163 4.5005
R82885 VDD.n1387 VDD.n1163 4.5005
R82886 VDD.n1300 VDD.n1163 4.5005
R82887 VDD.n1388 VDD.n1163 4.5005
R82888 VDD.n1298 VDD.n1163 4.5005
R82889 VDD.n1389 VDD.n1163 4.5005
R82890 VDD.n1297 VDD.n1163 4.5005
R82891 VDD.n1390 VDD.n1163 4.5005
R82892 VDD.n1295 VDD.n1163 4.5005
R82893 VDD.n1391 VDD.n1163 4.5005
R82894 VDD.n1294 VDD.n1163 4.5005
R82895 VDD.n1392 VDD.n1163 4.5005
R82896 VDD.n1292 VDD.n1163 4.5005
R82897 VDD.n1393 VDD.n1163 4.5005
R82898 VDD.n1291 VDD.n1163 4.5005
R82899 VDD.n1394 VDD.n1163 4.5005
R82900 VDD.n1289 VDD.n1163 4.5005
R82901 VDD.n1395 VDD.n1163 4.5005
R82902 VDD.n1288 VDD.n1163 4.5005
R82903 VDD.n1396 VDD.n1163 4.5005
R82904 VDD.n1286 VDD.n1163 4.5005
R82905 VDD.n1397 VDD.n1163 4.5005
R82906 VDD.n1285 VDD.n1163 4.5005
R82907 VDD.n1398 VDD.n1163 4.5005
R82908 VDD.n1283 VDD.n1163 4.5005
R82909 VDD.n1399 VDD.n1163 4.5005
R82910 VDD.n1282 VDD.n1163 4.5005
R82911 VDD.n1400 VDD.n1163 4.5005
R82912 VDD.n1280 VDD.n1163 4.5005
R82913 VDD.n1401 VDD.n1163 4.5005
R82914 VDD.n1279 VDD.n1163 4.5005
R82915 VDD.n1402 VDD.n1163 4.5005
R82916 VDD.n1277 VDD.n1163 4.5005
R82917 VDD.n1403 VDD.n1163 4.5005
R82918 VDD.n1276 VDD.n1163 4.5005
R82919 VDD.n1404 VDD.n1163 4.5005
R82920 VDD.n1274 VDD.n1163 4.5005
R82921 VDD.n1405 VDD.n1163 4.5005
R82922 VDD.n1273 VDD.n1163 4.5005
R82923 VDD.n1406 VDD.n1163 4.5005
R82924 VDD.n1271 VDD.n1163 4.5005
R82925 VDD.n1407 VDD.n1163 4.5005
R82926 VDD.n1270 VDD.n1163 4.5005
R82927 VDD.n1408 VDD.n1163 4.5005
R82928 VDD.n1268 VDD.n1163 4.5005
R82929 VDD.n1409 VDD.n1163 4.5005
R82930 VDD.n1267 VDD.n1163 4.5005
R82931 VDD.n1410 VDD.n1163 4.5005
R82932 VDD.n1265 VDD.n1163 4.5005
R82933 VDD.n1411 VDD.n1163 4.5005
R82934 VDD.n1264 VDD.n1163 4.5005
R82935 VDD.n1412 VDD.n1163 4.5005
R82936 VDD.n1262 VDD.n1163 4.5005
R82937 VDD.n1413 VDD.n1163 4.5005
R82938 VDD.n1261 VDD.n1163 4.5005
R82939 VDD.n1414 VDD.n1163 4.5005
R82940 VDD.n1415 VDD.n1163 4.5005
R82941 VDD.n1674 VDD.n1163 4.5005
R82942 VDD.n1676 VDD.n1227 4.5005
R82943 VDD.n1341 VDD.n1227 4.5005
R82944 VDD.n1342 VDD.n1227 4.5005
R82945 VDD.n1340 VDD.n1227 4.5005
R82946 VDD.n1344 VDD.n1227 4.5005
R82947 VDD.n1339 VDD.n1227 4.5005
R82948 VDD.n1345 VDD.n1227 4.5005
R82949 VDD.n1338 VDD.n1227 4.5005
R82950 VDD.n1347 VDD.n1227 4.5005
R82951 VDD.n1337 VDD.n1227 4.5005
R82952 VDD.n1348 VDD.n1227 4.5005
R82953 VDD.n1336 VDD.n1227 4.5005
R82954 VDD.n1350 VDD.n1227 4.5005
R82955 VDD.n1335 VDD.n1227 4.5005
R82956 VDD.n1351 VDD.n1227 4.5005
R82957 VDD.n1334 VDD.n1227 4.5005
R82958 VDD.n1353 VDD.n1227 4.5005
R82959 VDD.n1333 VDD.n1227 4.5005
R82960 VDD.n1354 VDD.n1227 4.5005
R82961 VDD.n1332 VDD.n1227 4.5005
R82962 VDD.n1356 VDD.n1227 4.5005
R82963 VDD.n1331 VDD.n1227 4.5005
R82964 VDD.n1357 VDD.n1227 4.5005
R82965 VDD.n1330 VDD.n1227 4.5005
R82966 VDD.n1359 VDD.n1227 4.5005
R82967 VDD.n1329 VDD.n1227 4.5005
R82968 VDD.n1360 VDD.n1227 4.5005
R82969 VDD.n1328 VDD.n1227 4.5005
R82970 VDD.n1362 VDD.n1227 4.5005
R82971 VDD.n1327 VDD.n1227 4.5005
R82972 VDD.n1363 VDD.n1227 4.5005
R82973 VDD.n1326 VDD.n1227 4.5005
R82974 VDD.n1365 VDD.n1227 4.5005
R82975 VDD.n1325 VDD.n1227 4.5005
R82976 VDD.n1366 VDD.n1227 4.5005
R82977 VDD.n1324 VDD.n1227 4.5005
R82978 VDD.n1368 VDD.n1227 4.5005
R82979 VDD.n1323 VDD.n1227 4.5005
R82980 VDD.n1369 VDD.n1227 4.5005
R82981 VDD.n1322 VDD.n1227 4.5005
R82982 VDD.n1371 VDD.n1227 4.5005
R82983 VDD.n1321 VDD.n1227 4.5005
R82984 VDD.n1372 VDD.n1227 4.5005
R82985 VDD.n1320 VDD.n1227 4.5005
R82986 VDD.n1374 VDD.n1227 4.5005
R82987 VDD.n1319 VDD.n1227 4.5005
R82988 VDD.n1375 VDD.n1227 4.5005
R82989 VDD.n1318 VDD.n1227 4.5005
R82990 VDD.n1376 VDD.n1227 4.5005
R82991 VDD.n1316 VDD.n1227 4.5005
R82992 VDD.n1377 VDD.n1227 4.5005
R82993 VDD.n1315 VDD.n1227 4.5005
R82994 VDD.n1378 VDD.n1227 4.5005
R82995 VDD.n1313 VDD.n1227 4.5005
R82996 VDD.n1379 VDD.n1227 4.5005
R82997 VDD.n1312 VDD.n1227 4.5005
R82998 VDD.n1380 VDD.n1227 4.5005
R82999 VDD.n1310 VDD.n1227 4.5005
R83000 VDD.n1381 VDD.n1227 4.5005
R83001 VDD.n1309 VDD.n1227 4.5005
R83002 VDD.n1382 VDD.n1227 4.5005
R83003 VDD.n1307 VDD.n1227 4.5005
R83004 VDD.n1383 VDD.n1227 4.5005
R83005 VDD.n1306 VDD.n1227 4.5005
R83006 VDD.n1384 VDD.n1227 4.5005
R83007 VDD.n1304 VDD.n1227 4.5005
R83008 VDD.n1385 VDD.n1227 4.5005
R83009 VDD.n1303 VDD.n1227 4.5005
R83010 VDD.n1386 VDD.n1227 4.5005
R83011 VDD.n1301 VDD.n1227 4.5005
R83012 VDD.n1387 VDD.n1227 4.5005
R83013 VDD.n1300 VDD.n1227 4.5005
R83014 VDD.n1388 VDD.n1227 4.5005
R83015 VDD.n1298 VDD.n1227 4.5005
R83016 VDD.n1389 VDD.n1227 4.5005
R83017 VDD.n1297 VDD.n1227 4.5005
R83018 VDD.n1390 VDD.n1227 4.5005
R83019 VDD.n1295 VDD.n1227 4.5005
R83020 VDD.n1391 VDD.n1227 4.5005
R83021 VDD.n1294 VDD.n1227 4.5005
R83022 VDD.n1392 VDD.n1227 4.5005
R83023 VDD.n1292 VDD.n1227 4.5005
R83024 VDD.n1393 VDD.n1227 4.5005
R83025 VDD.n1291 VDD.n1227 4.5005
R83026 VDD.n1394 VDD.n1227 4.5005
R83027 VDD.n1289 VDD.n1227 4.5005
R83028 VDD.n1395 VDD.n1227 4.5005
R83029 VDD.n1288 VDD.n1227 4.5005
R83030 VDD.n1396 VDD.n1227 4.5005
R83031 VDD.n1286 VDD.n1227 4.5005
R83032 VDD.n1397 VDD.n1227 4.5005
R83033 VDD.n1285 VDD.n1227 4.5005
R83034 VDD.n1398 VDD.n1227 4.5005
R83035 VDD.n1283 VDD.n1227 4.5005
R83036 VDD.n1399 VDD.n1227 4.5005
R83037 VDD.n1282 VDD.n1227 4.5005
R83038 VDD.n1400 VDD.n1227 4.5005
R83039 VDD.n1280 VDD.n1227 4.5005
R83040 VDD.n1401 VDD.n1227 4.5005
R83041 VDD.n1279 VDD.n1227 4.5005
R83042 VDD.n1402 VDD.n1227 4.5005
R83043 VDD.n1277 VDD.n1227 4.5005
R83044 VDD.n1403 VDD.n1227 4.5005
R83045 VDD.n1276 VDD.n1227 4.5005
R83046 VDD.n1404 VDD.n1227 4.5005
R83047 VDD.n1274 VDD.n1227 4.5005
R83048 VDD.n1405 VDD.n1227 4.5005
R83049 VDD.n1273 VDD.n1227 4.5005
R83050 VDD.n1406 VDD.n1227 4.5005
R83051 VDD.n1271 VDD.n1227 4.5005
R83052 VDD.n1407 VDD.n1227 4.5005
R83053 VDD.n1270 VDD.n1227 4.5005
R83054 VDD.n1408 VDD.n1227 4.5005
R83055 VDD.n1268 VDD.n1227 4.5005
R83056 VDD.n1409 VDD.n1227 4.5005
R83057 VDD.n1267 VDD.n1227 4.5005
R83058 VDD.n1410 VDD.n1227 4.5005
R83059 VDD.n1265 VDD.n1227 4.5005
R83060 VDD.n1411 VDD.n1227 4.5005
R83061 VDD.n1264 VDD.n1227 4.5005
R83062 VDD.n1412 VDD.n1227 4.5005
R83063 VDD.n1262 VDD.n1227 4.5005
R83064 VDD.n1413 VDD.n1227 4.5005
R83065 VDD.n1261 VDD.n1227 4.5005
R83066 VDD.n1414 VDD.n1227 4.5005
R83067 VDD.n1415 VDD.n1227 4.5005
R83068 VDD.n1674 VDD.n1227 4.5005
R83069 VDD.n1676 VDD.n1162 4.5005
R83070 VDD.n1341 VDD.n1162 4.5005
R83071 VDD.n1342 VDD.n1162 4.5005
R83072 VDD.n1340 VDD.n1162 4.5005
R83073 VDD.n1344 VDD.n1162 4.5005
R83074 VDD.n1339 VDD.n1162 4.5005
R83075 VDD.n1345 VDD.n1162 4.5005
R83076 VDD.n1338 VDD.n1162 4.5005
R83077 VDD.n1347 VDD.n1162 4.5005
R83078 VDD.n1337 VDD.n1162 4.5005
R83079 VDD.n1348 VDD.n1162 4.5005
R83080 VDD.n1336 VDD.n1162 4.5005
R83081 VDD.n1350 VDD.n1162 4.5005
R83082 VDD.n1335 VDD.n1162 4.5005
R83083 VDD.n1351 VDD.n1162 4.5005
R83084 VDD.n1334 VDD.n1162 4.5005
R83085 VDD.n1353 VDD.n1162 4.5005
R83086 VDD.n1333 VDD.n1162 4.5005
R83087 VDD.n1354 VDD.n1162 4.5005
R83088 VDD.n1332 VDD.n1162 4.5005
R83089 VDD.n1356 VDD.n1162 4.5005
R83090 VDD.n1331 VDD.n1162 4.5005
R83091 VDD.n1357 VDD.n1162 4.5005
R83092 VDD.n1330 VDD.n1162 4.5005
R83093 VDD.n1359 VDD.n1162 4.5005
R83094 VDD.n1329 VDD.n1162 4.5005
R83095 VDD.n1360 VDD.n1162 4.5005
R83096 VDD.n1328 VDD.n1162 4.5005
R83097 VDD.n1362 VDD.n1162 4.5005
R83098 VDD.n1327 VDD.n1162 4.5005
R83099 VDD.n1363 VDD.n1162 4.5005
R83100 VDD.n1326 VDD.n1162 4.5005
R83101 VDD.n1365 VDD.n1162 4.5005
R83102 VDD.n1325 VDD.n1162 4.5005
R83103 VDD.n1366 VDD.n1162 4.5005
R83104 VDD.n1324 VDD.n1162 4.5005
R83105 VDD.n1368 VDD.n1162 4.5005
R83106 VDD.n1323 VDD.n1162 4.5005
R83107 VDD.n1369 VDD.n1162 4.5005
R83108 VDD.n1322 VDD.n1162 4.5005
R83109 VDD.n1371 VDD.n1162 4.5005
R83110 VDD.n1321 VDD.n1162 4.5005
R83111 VDD.n1372 VDD.n1162 4.5005
R83112 VDD.n1320 VDD.n1162 4.5005
R83113 VDD.n1374 VDD.n1162 4.5005
R83114 VDD.n1319 VDD.n1162 4.5005
R83115 VDD.n1375 VDD.n1162 4.5005
R83116 VDD.n1318 VDD.n1162 4.5005
R83117 VDD.n1376 VDD.n1162 4.5005
R83118 VDD.n1316 VDD.n1162 4.5005
R83119 VDD.n1377 VDD.n1162 4.5005
R83120 VDD.n1315 VDD.n1162 4.5005
R83121 VDD.n1378 VDD.n1162 4.5005
R83122 VDD.n1313 VDD.n1162 4.5005
R83123 VDD.n1379 VDD.n1162 4.5005
R83124 VDD.n1312 VDD.n1162 4.5005
R83125 VDD.n1380 VDD.n1162 4.5005
R83126 VDD.n1310 VDD.n1162 4.5005
R83127 VDD.n1381 VDD.n1162 4.5005
R83128 VDD.n1309 VDD.n1162 4.5005
R83129 VDD.n1382 VDD.n1162 4.5005
R83130 VDD.n1307 VDD.n1162 4.5005
R83131 VDD.n1383 VDD.n1162 4.5005
R83132 VDD.n1306 VDD.n1162 4.5005
R83133 VDD.n1384 VDD.n1162 4.5005
R83134 VDD.n1304 VDD.n1162 4.5005
R83135 VDD.n1385 VDD.n1162 4.5005
R83136 VDD.n1303 VDD.n1162 4.5005
R83137 VDD.n1386 VDD.n1162 4.5005
R83138 VDD.n1301 VDD.n1162 4.5005
R83139 VDD.n1387 VDD.n1162 4.5005
R83140 VDD.n1300 VDD.n1162 4.5005
R83141 VDD.n1388 VDD.n1162 4.5005
R83142 VDD.n1298 VDD.n1162 4.5005
R83143 VDD.n1389 VDD.n1162 4.5005
R83144 VDD.n1297 VDD.n1162 4.5005
R83145 VDD.n1390 VDD.n1162 4.5005
R83146 VDD.n1295 VDD.n1162 4.5005
R83147 VDD.n1391 VDD.n1162 4.5005
R83148 VDD.n1294 VDD.n1162 4.5005
R83149 VDD.n1392 VDD.n1162 4.5005
R83150 VDD.n1292 VDD.n1162 4.5005
R83151 VDD.n1393 VDD.n1162 4.5005
R83152 VDD.n1291 VDD.n1162 4.5005
R83153 VDD.n1394 VDD.n1162 4.5005
R83154 VDD.n1289 VDD.n1162 4.5005
R83155 VDD.n1395 VDD.n1162 4.5005
R83156 VDD.n1288 VDD.n1162 4.5005
R83157 VDD.n1396 VDD.n1162 4.5005
R83158 VDD.n1286 VDD.n1162 4.5005
R83159 VDD.n1397 VDD.n1162 4.5005
R83160 VDD.n1285 VDD.n1162 4.5005
R83161 VDD.n1398 VDD.n1162 4.5005
R83162 VDD.n1283 VDD.n1162 4.5005
R83163 VDD.n1399 VDD.n1162 4.5005
R83164 VDD.n1282 VDD.n1162 4.5005
R83165 VDD.n1400 VDD.n1162 4.5005
R83166 VDD.n1280 VDD.n1162 4.5005
R83167 VDD.n1401 VDD.n1162 4.5005
R83168 VDD.n1279 VDD.n1162 4.5005
R83169 VDD.n1402 VDD.n1162 4.5005
R83170 VDD.n1277 VDD.n1162 4.5005
R83171 VDD.n1403 VDD.n1162 4.5005
R83172 VDD.n1276 VDD.n1162 4.5005
R83173 VDD.n1404 VDD.n1162 4.5005
R83174 VDD.n1274 VDD.n1162 4.5005
R83175 VDD.n1405 VDD.n1162 4.5005
R83176 VDD.n1273 VDD.n1162 4.5005
R83177 VDD.n1406 VDD.n1162 4.5005
R83178 VDD.n1271 VDD.n1162 4.5005
R83179 VDD.n1407 VDD.n1162 4.5005
R83180 VDD.n1270 VDD.n1162 4.5005
R83181 VDD.n1408 VDD.n1162 4.5005
R83182 VDD.n1268 VDD.n1162 4.5005
R83183 VDD.n1409 VDD.n1162 4.5005
R83184 VDD.n1267 VDD.n1162 4.5005
R83185 VDD.n1410 VDD.n1162 4.5005
R83186 VDD.n1265 VDD.n1162 4.5005
R83187 VDD.n1411 VDD.n1162 4.5005
R83188 VDD.n1264 VDD.n1162 4.5005
R83189 VDD.n1412 VDD.n1162 4.5005
R83190 VDD.n1262 VDD.n1162 4.5005
R83191 VDD.n1413 VDD.n1162 4.5005
R83192 VDD.n1261 VDD.n1162 4.5005
R83193 VDD.n1414 VDD.n1162 4.5005
R83194 VDD.n1415 VDD.n1162 4.5005
R83195 VDD.n1674 VDD.n1162 4.5005
R83196 VDD.n1676 VDD.n1228 4.5005
R83197 VDD.n1341 VDD.n1228 4.5005
R83198 VDD.n1342 VDD.n1228 4.5005
R83199 VDD.n1340 VDD.n1228 4.5005
R83200 VDD.n1344 VDD.n1228 4.5005
R83201 VDD.n1339 VDD.n1228 4.5005
R83202 VDD.n1345 VDD.n1228 4.5005
R83203 VDD.n1338 VDD.n1228 4.5005
R83204 VDD.n1347 VDD.n1228 4.5005
R83205 VDD.n1337 VDD.n1228 4.5005
R83206 VDD.n1348 VDD.n1228 4.5005
R83207 VDD.n1336 VDD.n1228 4.5005
R83208 VDD.n1350 VDD.n1228 4.5005
R83209 VDD.n1335 VDD.n1228 4.5005
R83210 VDD.n1351 VDD.n1228 4.5005
R83211 VDD.n1334 VDD.n1228 4.5005
R83212 VDD.n1353 VDD.n1228 4.5005
R83213 VDD.n1333 VDD.n1228 4.5005
R83214 VDD.n1354 VDD.n1228 4.5005
R83215 VDD.n1332 VDD.n1228 4.5005
R83216 VDD.n1356 VDD.n1228 4.5005
R83217 VDD.n1331 VDD.n1228 4.5005
R83218 VDD.n1357 VDD.n1228 4.5005
R83219 VDD.n1330 VDD.n1228 4.5005
R83220 VDD.n1359 VDD.n1228 4.5005
R83221 VDD.n1329 VDD.n1228 4.5005
R83222 VDD.n1360 VDD.n1228 4.5005
R83223 VDD.n1328 VDD.n1228 4.5005
R83224 VDD.n1362 VDD.n1228 4.5005
R83225 VDD.n1327 VDD.n1228 4.5005
R83226 VDD.n1363 VDD.n1228 4.5005
R83227 VDD.n1326 VDD.n1228 4.5005
R83228 VDD.n1365 VDD.n1228 4.5005
R83229 VDD.n1325 VDD.n1228 4.5005
R83230 VDD.n1366 VDD.n1228 4.5005
R83231 VDD.n1324 VDD.n1228 4.5005
R83232 VDD.n1368 VDD.n1228 4.5005
R83233 VDD.n1323 VDD.n1228 4.5005
R83234 VDD.n1369 VDD.n1228 4.5005
R83235 VDD.n1322 VDD.n1228 4.5005
R83236 VDD.n1371 VDD.n1228 4.5005
R83237 VDD.n1321 VDD.n1228 4.5005
R83238 VDD.n1372 VDD.n1228 4.5005
R83239 VDD.n1320 VDD.n1228 4.5005
R83240 VDD.n1374 VDD.n1228 4.5005
R83241 VDD.n1319 VDD.n1228 4.5005
R83242 VDD.n1375 VDD.n1228 4.5005
R83243 VDD.n1318 VDD.n1228 4.5005
R83244 VDD.n1376 VDD.n1228 4.5005
R83245 VDD.n1316 VDD.n1228 4.5005
R83246 VDD.n1377 VDD.n1228 4.5005
R83247 VDD.n1315 VDD.n1228 4.5005
R83248 VDD.n1378 VDD.n1228 4.5005
R83249 VDD.n1313 VDD.n1228 4.5005
R83250 VDD.n1379 VDD.n1228 4.5005
R83251 VDD.n1312 VDD.n1228 4.5005
R83252 VDD.n1380 VDD.n1228 4.5005
R83253 VDD.n1310 VDD.n1228 4.5005
R83254 VDD.n1381 VDD.n1228 4.5005
R83255 VDD.n1309 VDD.n1228 4.5005
R83256 VDD.n1382 VDD.n1228 4.5005
R83257 VDD.n1307 VDD.n1228 4.5005
R83258 VDD.n1383 VDD.n1228 4.5005
R83259 VDD.n1306 VDD.n1228 4.5005
R83260 VDD.n1384 VDD.n1228 4.5005
R83261 VDD.n1304 VDD.n1228 4.5005
R83262 VDD.n1385 VDD.n1228 4.5005
R83263 VDD.n1303 VDD.n1228 4.5005
R83264 VDD.n1386 VDD.n1228 4.5005
R83265 VDD.n1301 VDD.n1228 4.5005
R83266 VDD.n1387 VDD.n1228 4.5005
R83267 VDD.n1300 VDD.n1228 4.5005
R83268 VDD.n1388 VDD.n1228 4.5005
R83269 VDD.n1298 VDD.n1228 4.5005
R83270 VDD.n1389 VDD.n1228 4.5005
R83271 VDD.n1297 VDD.n1228 4.5005
R83272 VDD.n1390 VDD.n1228 4.5005
R83273 VDD.n1295 VDD.n1228 4.5005
R83274 VDD.n1391 VDD.n1228 4.5005
R83275 VDD.n1294 VDD.n1228 4.5005
R83276 VDD.n1392 VDD.n1228 4.5005
R83277 VDD.n1292 VDD.n1228 4.5005
R83278 VDD.n1393 VDD.n1228 4.5005
R83279 VDD.n1291 VDD.n1228 4.5005
R83280 VDD.n1394 VDD.n1228 4.5005
R83281 VDD.n1289 VDD.n1228 4.5005
R83282 VDD.n1395 VDD.n1228 4.5005
R83283 VDD.n1288 VDD.n1228 4.5005
R83284 VDD.n1396 VDD.n1228 4.5005
R83285 VDD.n1286 VDD.n1228 4.5005
R83286 VDD.n1397 VDD.n1228 4.5005
R83287 VDD.n1285 VDD.n1228 4.5005
R83288 VDD.n1398 VDD.n1228 4.5005
R83289 VDD.n1283 VDD.n1228 4.5005
R83290 VDD.n1399 VDD.n1228 4.5005
R83291 VDD.n1282 VDD.n1228 4.5005
R83292 VDD.n1400 VDD.n1228 4.5005
R83293 VDD.n1280 VDD.n1228 4.5005
R83294 VDD.n1401 VDD.n1228 4.5005
R83295 VDD.n1279 VDD.n1228 4.5005
R83296 VDD.n1402 VDD.n1228 4.5005
R83297 VDD.n1277 VDD.n1228 4.5005
R83298 VDD.n1403 VDD.n1228 4.5005
R83299 VDD.n1276 VDD.n1228 4.5005
R83300 VDD.n1404 VDD.n1228 4.5005
R83301 VDD.n1274 VDD.n1228 4.5005
R83302 VDD.n1405 VDD.n1228 4.5005
R83303 VDD.n1273 VDD.n1228 4.5005
R83304 VDD.n1406 VDD.n1228 4.5005
R83305 VDD.n1271 VDD.n1228 4.5005
R83306 VDD.n1407 VDD.n1228 4.5005
R83307 VDD.n1270 VDD.n1228 4.5005
R83308 VDD.n1408 VDD.n1228 4.5005
R83309 VDD.n1268 VDD.n1228 4.5005
R83310 VDD.n1409 VDD.n1228 4.5005
R83311 VDD.n1267 VDD.n1228 4.5005
R83312 VDD.n1410 VDD.n1228 4.5005
R83313 VDD.n1265 VDD.n1228 4.5005
R83314 VDD.n1411 VDD.n1228 4.5005
R83315 VDD.n1264 VDD.n1228 4.5005
R83316 VDD.n1412 VDD.n1228 4.5005
R83317 VDD.n1262 VDD.n1228 4.5005
R83318 VDD.n1413 VDD.n1228 4.5005
R83319 VDD.n1261 VDD.n1228 4.5005
R83320 VDD.n1414 VDD.n1228 4.5005
R83321 VDD.n1415 VDD.n1228 4.5005
R83322 VDD.n1674 VDD.n1228 4.5005
R83323 VDD.n1676 VDD.n1161 4.5005
R83324 VDD.n1341 VDD.n1161 4.5005
R83325 VDD.n1342 VDD.n1161 4.5005
R83326 VDD.n1340 VDD.n1161 4.5005
R83327 VDD.n1344 VDD.n1161 4.5005
R83328 VDD.n1339 VDD.n1161 4.5005
R83329 VDD.n1345 VDD.n1161 4.5005
R83330 VDD.n1338 VDD.n1161 4.5005
R83331 VDD.n1347 VDD.n1161 4.5005
R83332 VDD.n1337 VDD.n1161 4.5005
R83333 VDD.n1348 VDD.n1161 4.5005
R83334 VDD.n1336 VDD.n1161 4.5005
R83335 VDD.n1350 VDD.n1161 4.5005
R83336 VDD.n1335 VDD.n1161 4.5005
R83337 VDD.n1351 VDD.n1161 4.5005
R83338 VDD.n1334 VDD.n1161 4.5005
R83339 VDD.n1353 VDD.n1161 4.5005
R83340 VDD.n1333 VDD.n1161 4.5005
R83341 VDD.n1354 VDD.n1161 4.5005
R83342 VDD.n1332 VDD.n1161 4.5005
R83343 VDD.n1356 VDD.n1161 4.5005
R83344 VDD.n1331 VDD.n1161 4.5005
R83345 VDD.n1357 VDD.n1161 4.5005
R83346 VDD.n1330 VDD.n1161 4.5005
R83347 VDD.n1359 VDD.n1161 4.5005
R83348 VDD.n1329 VDD.n1161 4.5005
R83349 VDD.n1360 VDD.n1161 4.5005
R83350 VDD.n1328 VDD.n1161 4.5005
R83351 VDD.n1362 VDD.n1161 4.5005
R83352 VDD.n1327 VDD.n1161 4.5005
R83353 VDD.n1363 VDD.n1161 4.5005
R83354 VDD.n1326 VDD.n1161 4.5005
R83355 VDD.n1365 VDD.n1161 4.5005
R83356 VDD.n1325 VDD.n1161 4.5005
R83357 VDD.n1366 VDD.n1161 4.5005
R83358 VDD.n1324 VDD.n1161 4.5005
R83359 VDD.n1368 VDD.n1161 4.5005
R83360 VDD.n1323 VDD.n1161 4.5005
R83361 VDD.n1369 VDD.n1161 4.5005
R83362 VDD.n1322 VDD.n1161 4.5005
R83363 VDD.n1371 VDD.n1161 4.5005
R83364 VDD.n1321 VDD.n1161 4.5005
R83365 VDD.n1372 VDD.n1161 4.5005
R83366 VDD.n1320 VDD.n1161 4.5005
R83367 VDD.n1374 VDD.n1161 4.5005
R83368 VDD.n1319 VDD.n1161 4.5005
R83369 VDD.n1375 VDD.n1161 4.5005
R83370 VDD.n1318 VDD.n1161 4.5005
R83371 VDD.n1376 VDD.n1161 4.5005
R83372 VDD.n1316 VDD.n1161 4.5005
R83373 VDD.n1377 VDD.n1161 4.5005
R83374 VDD.n1315 VDD.n1161 4.5005
R83375 VDD.n1378 VDD.n1161 4.5005
R83376 VDD.n1313 VDD.n1161 4.5005
R83377 VDD.n1379 VDD.n1161 4.5005
R83378 VDD.n1312 VDD.n1161 4.5005
R83379 VDD.n1380 VDD.n1161 4.5005
R83380 VDD.n1310 VDD.n1161 4.5005
R83381 VDD.n1381 VDD.n1161 4.5005
R83382 VDD.n1309 VDD.n1161 4.5005
R83383 VDD.n1382 VDD.n1161 4.5005
R83384 VDD.n1307 VDD.n1161 4.5005
R83385 VDD.n1383 VDD.n1161 4.5005
R83386 VDD.n1306 VDD.n1161 4.5005
R83387 VDD.n1384 VDD.n1161 4.5005
R83388 VDD.n1304 VDD.n1161 4.5005
R83389 VDD.n1385 VDD.n1161 4.5005
R83390 VDD.n1303 VDD.n1161 4.5005
R83391 VDD.n1386 VDD.n1161 4.5005
R83392 VDD.n1301 VDD.n1161 4.5005
R83393 VDD.n1387 VDD.n1161 4.5005
R83394 VDD.n1300 VDD.n1161 4.5005
R83395 VDD.n1388 VDD.n1161 4.5005
R83396 VDD.n1298 VDD.n1161 4.5005
R83397 VDD.n1389 VDD.n1161 4.5005
R83398 VDD.n1297 VDD.n1161 4.5005
R83399 VDD.n1390 VDD.n1161 4.5005
R83400 VDD.n1295 VDD.n1161 4.5005
R83401 VDD.n1391 VDD.n1161 4.5005
R83402 VDD.n1294 VDD.n1161 4.5005
R83403 VDD.n1392 VDD.n1161 4.5005
R83404 VDD.n1292 VDD.n1161 4.5005
R83405 VDD.n1393 VDD.n1161 4.5005
R83406 VDD.n1291 VDD.n1161 4.5005
R83407 VDD.n1394 VDD.n1161 4.5005
R83408 VDD.n1289 VDD.n1161 4.5005
R83409 VDD.n1395 VDD.n1161 4.5005
R83410 VDD.n1288 VDD.n1161 4.5005
R83411 VDD.n1396 VDD.n1161 4.5005
R83412 VDD.n1286 VDD.n1161 4.5005
R83413 VDD.n1397 VDD.n1161 4.5005
R83414 VDD.n1285 VDD.n1161 4.5005
R83415 VDD.n1398 VDD.n1161 4.5005
R83416 VDD.n1283 VDD.n1161 4.5005
R83417 VDD.n1399 VDD.n1161 4.5005
R83418 VDD.n1282 VDD.n1161 4.5005
R83419 VDD.n1400 VDD.n1161 4.5005
R83420 VDD.n1280 VDD.n1161 4.5005
R83421 VDD.n1401 VDD.n1161 4.5005
R83422 VDD.n1279 VDD.n1161 4.5005
R83423 VDD.n1402 VDD.n1161 4.5005
R83424 VDD.n1277 VDD.n1161 4.5005
R83425 VDD.n1403 VDD.n1161 4.5005
R83426 VDD.n1276 VDD.n1161 4.5005
R83427 VDD.n1404 VDD.n1161 4.5005
R83428 VDD.n1274 VDD.n1161 4.5005
R83429 VDD.n1405 VDD.n1161 4.5005
R83430 VDD.n1273 VDD.n1161 4.5005
R83431 VDD.n1406 VDD.n1161 4.5005
R83432 VDD.n1271 VDD.n1161 4.5005
R83433 VDD.n1407 VDD.n1161 4.5005
R83434 VDD.n1270 VDD.n1161 4.5005
R83435 VDD.n1408 VDD.n1161 4.5005
R83436 VDD.n1268 VDD.n1161 4.5005
R83437 VDD.n1409 VDD.n1161 4.5005
R83438 VDD.n1267 VDD.n1161 4.5005
R83439 VDD.n1410 VDD.n1161 4.5005
R83440 VDD.n1265 VDD.n1161 4.5005
R83441 VDD.n1411 VDD.n1161 4.5005
R83442 VDD.n1264 VDD.n1161 4.5005
R83443 VDD.n1412 VDD.n1161 4.5005
R83444 VDD.n1262 VDD.n1161 4.5005
R83445 VDD.n1413 VDD.n1161 4.5005
R83446 VDD.n1261 VDD.n1161 4.5005
R83447 VDD.n1414 VDD.n1161 4.5005
R83448 VDD.n1415 VDD.n1161 4.5005
R83449 VDD.n1674 VDD.n1161 4.5005
R83450 VDD.n1676 VDD.n1229 4.5005
R83451 VDD.n1341 VDD.n1229 4.5005
R83452 VDD.n1342 VDD.n1229 4.5005
R83453 VDD.n1340 VDD.n1229 4.5005
R83454 VDD.n1344 VDD.n1229 4.5005
R83455 VDD.n1339 VDD.n1229 4.5005
R83456 VDD.n1345 VDD.n1229 4.5005
R83457 VDD.n1338 VDD.n1229 4.5005
R83458 VDD.n1347 VDD.n1229 4.5005
R83459 VDD.n1337 VDD.n1229 4.5005
R83460 VDD.n1348 VDD.n1229 4.5005
R83461 VDD.n1336 VDD.n1229 4.5005
R83462 VDD.n1350 VDD.n1229 4.5005
R83463 VDD.n1335 VDD.n1229 4.5005
R83464 VDD.n1351 VDD.n1229 4.5005
R83465 VDD.n1334 VDD.n1229 4.5005
R83466 VDD.n1353 VDD.n1229 4.5005
R83467 VDD.n1333 VDD.n1229 4.5005
R83468 VDD.n1354 VDD.n1229 4.5005
R83469 VDD.n1332 VDD.n1229 4.5005
R83470 VDD.n1356 VDD.n1229 4.5005
R83471 VDD.n1331 VDD.n1229 4.5005
R83472 VDD.n1357 VDD.n1229 4.5005
R83473 VDD.n1330 VDD.n1229 4.5005
R83474 VDD.n1359 VDD.n1229 4.5005
R83475 VDD.n1329 VDD.n1229 4.5005
R83476 VDD.n1360 VDD.n1229 4.5005
R83477 VDD.n1328 VDD.n1229 4.5005
R83478 VDD.n1362 VDD.n1229 4.5005
R83479 VDD.n1327 VDD.n1229 4.5005
R83480 VDD.n1363 VDD.n1229 4.5005
R83481 VDD.n1326 VDD.n1229 4.5005
R83482 VDD.n1365 VDD.n1229 4.5005
R83483 VDD.n1325 VDD.n1229 4.5005
R83484 VDD.n1366 VDD.n1229 4.5005
R83485 VDD.n1324 VDD.n1229 4.5005
R83486 VDD.n1368 VDD.n1229 4.5005
R83487 VDD.n1323 VDD.n1229 4.5005
R83488 VDD.n1369 VDD.n1229 4.5005
R83489 VDD.n1322 VDD.n1229 4.5005
R83490 VDD.n1371 VDD.n1229 4.5005
R83491 VDD.n1321 VDD.n1229 4.5005
R83492 VDD.n1372 VDD.n1229 4.5005
R83493 VDD.n1320 VDD.n1229 4.5005
R83494 VDD.n1374 VDD.n1229 4.5005
R83495 VDD.n1319 VDD.n1229 4.5005
R83496 VDD.n1375 VDD.n1229 4.5005
R83497 VDD.n1318 VDD.n1229 4.5005
R83498 VDD.n1376 VDD.n1229 4.5005
R83499 VDD.n1316 VDD.n1229 4.5005
R83500 VDD.n1377 VDD.n1229 4.5005
R83501 VDD.n1315 VDD.n1229 4.5005
R83502 VDD.n1378 VDD.n1229 4.5005
R83503 VDD.n1313 VDD.n1229 4.5005
R83504 VDD.n1379 VDD.n1229 4.5005
R83505 VDD.n1312 VDD.n1229 4.5005
R83506 VDD.n1380 VDD.n1229 4.5005
R83507 VDD.n1310 VDD.n1229 4.5005
R83508 VDD.n1381 VDD.n1229 4.5005
R83509 VDD.n1309 VDD.n1229 4.5005
R83510 VDD.n1382 VDD.n1229 4.5005
R83511 VDD.n1307 VDD.n1229 4.5005
R83512 VDD.n1383 VDD.n1229 4.5005
R83513 VDD.n1306 VDD.n1229 4.5005
R83514 VDD.n1384 VDD.n1229 4.5005
R83515 VDD.n1304 VDD.n1229 4.5005
R83516 VDD.n1385 VDD.n1229 4.5005
R83517 VDD.n1303 VDD.n1229 4.5005
R83518 VDD.n1386 VDD.n1229 4.5005
R83519 VDD.n1301 VDD.n1229 4.5005
R83520 VDD.n1387 VDD.n1229 4.5005
R83521 VDD.n1300 VDD.n1229 4.5005
R83522 VDD.n1388 VDD.n1229 4.5005
R83523 VDD.n1298 VDD.n1229 4.5005
R83524 VDD.n1389 VDD.n1229 4.5005
R83525 VDD.n1297 VDD.n1229 4.5005
R83526 VDD.n1390 VDD.n1229 4.5005
R83527 VDD.n1295 VDD.n1229 4.5005
R83528 VDD.n1391 VDD.n1229 4.5005
R83529 VDD.n1294 VDD.n1229 4.5005
R83530 VDD.n1392 VDD.n1229 4.5005
R83531 VDD.n1292 VDD.n1229 4.5005
R83532 VDD.n1393 VDD.n1229 4.5005
R83533 VDD.n1291 VDD.n1229 4.5005
R83534 VDD.n1394 VDD.n1229 4.5005
R83535 VDD.n1289 VDD.n1229 4.5005
R83536 VDD.n1395 VDD.n1229 4.5005
R83537 VDD.n1288 VDD.n1229 4.5005
R83538 VDD.n1396 VDD.n1229 4.5005
R83539 VDD.n1286 VDD.n1229 4.5005
R83540 VDD.n1397 VDD.n1229 4.5005
R83541 VDD.n1285 VDD.n1229 4.5005
R83542 VDD.n1398 VDD.n1229 4.5005
R83543 VDD.n1283 VDD.n1229 4.5005
R83544 VDD.n1399 VDD.n1229 4.5005
R83545 VDD.n1282 VDD.n1229 4.5005
R83546 VDD.n1400 VDD.n1229 4.5005
R83547 VDD.n1280 VDD.n1229 4.5005
R83548 VDD.n1401 VDD.n1229 4.5005
R83549 VDD.n1279 VDD.n1229 4.5005
R83550 VDD.n1402 VDD.n1229 4.5005
R83551 VDD.n1277 VDD.n1229 4.5005
R83552 VDD.n1403 VDD.n1229 4.5005
R83553 VDD.n1276 VDD.n1229 4.5005
R83554 VDD.n1404 VDD.n1229 4.5005
R83555 VDD.n1274 VDD.n1229 4.5005
R83556 VDD.n1405 VDD.n1229 4.5005
R83557 VDD.n1273 VDD.n1229 4.5005
R83558 VDD.n1406 VDD.n1229 4.5005
R83559 VDD.n1271 VDD.n1229 4.5005
R83560 VDD.n1407 VDD.n1229 4.5005
R83561 VDD.n1270 VDD.n1229 4.5005
R83562 VDD.n1408 VDD.n1229 4.5005
R83563 VDD.n1268 VDD.n1229 4.5005
R83564 VDD.n1409 VDD.n1229 4.5005
R83565 VDD.n1267 VDD.n1229 4.5005
R83566 VDD.n1410 VDD.n1229 4.5005
R83567 VDD.n1265 VDD.n1229 4.5005
R83568 VDD.n1411 VDD.n1229 4.5005
R83569 VDD.n1264 VDD.n1229 4.5005
R83570 VDD.n1412 VDD.n1229 4.5005
R83571 VDD.n1262 VDD.n1229 4.5005
R83572 VDD.n1413 VDD.n1229 4.5005
R83573 VDD.n1261 VDD.n1229 4.5005
R83574 VDD.n1414 VDD.n1229 4.5005
R83575 VDD.n1415 VDD.n1229 4.5005
R83576 VDD.n1674 VDD.n1229 4.5005
R83577 VDD.n1676 VDD.n1160 4.5005
R83578 VDD.n1341 VDD.n1160 4.5005
R83579 VDD.n1342 VDD.n1160 4.5005
R83580 VDD.n1340 VDD.n1160 4.5005
R83581 VDD.n1344 VDD.n1160 4.5005
R83582 VDD.n1339 VDD.n1160 4.5005
R83583 VDD.n1345 VDD.n1160 4.5005
R83584 VDD.n1338 VDD.n1160 4.5005
R83585 VDD.n1347 VDD.n1160 4.5005
R83586 VDD.n1337 VDD.n1160 4.5005
R83587 VDD.n1348 VDD.n1160 4.5005
R83588 VDD.n1336 VDD.n1160 4.5005
R83589 VDD.n1350 VDD.n1160 4.5005
R83590 VDD.n1335 VDD.n1160 4.5005
R83591 VDD.n1351 VDD.n1160 4.5005
R83592 VDD.n1334 VDD.n1160 4.5005
R83593 VDD.n1353 VDD.n1160 4.5005
R83594 VDD.n1333 VDD.n1160 4.5005
R83595 VDD.n1354 VDD.n1160 4.5005
R83596 VDD.n1332 VDD.n1160 4.5005
R83597 VDD.n1356 VDD.n1160 4.5005
R83598 VDD.n1331 VDD.n1160 4.5005
R83599 VDD.n1357 VDD.n1160 4.5005
R83600 VDD.n1330 VDD.n1160 4.5005
R83601 VDD.n1359 VDD.n1160 4.5005
R83602 VDD.n1329 VDD.n1160 4.5005
R83603 VDD.n1360 VDD.n1160 4.5005
R83604 VDD.n1328 VDD.n1160 4.5005
R83605 VDD.n1362 VDD.n1160 4.5005
R83606 VDD.n1327 VDD.n1160 4.5005
R83607 VDD.n1363 VDD.n1160 4.5005
R83608 VDD.n1326 VDD.n1160 4.5005
R83609 VDD.n1365 VDD.n1160 4.5005
R83610 VDD.n1325 VDD.n1160 4.5005
R83611 VDD.n1366 VDD.n1160 4.5005
R83612 VDD.n1324 VDD.n1160 4.5005
R83613 VDD.n1368 VDD.n1160 4.5005
R83614 VDD.n1323 VDD.n1160 4.5005
R83615 VDD.n1369 VDD.n1160 4.5005
R83616 VDD.n1322 VDD.n1160 4.5005
R83617 VDD.n1371 VDD.n1160 4.5005
R83618 VDD.n1321 VDD.n1160 4.5005
R83619 VDD.n1372 VDD.n1160 4.5005
R83620 VDD.n1320 VDD.n1160 4.5005
R83621 VDD.n1374 VDD.n1160 4.5005
R83622 VDD.n1319 VDD.n1160 4.5005
R83623 VDD.n1375 VDD.n1160 4.5005
R83624 VDD.n1318 VDD.n1160 4.5005
R83625 VDD.n1376 VDD.n1160 4.5005
R83626 VDD.n1316 VDD.n1160 4.5005
R83627 VDD.n1377 VDD.n1160 4.5005
R83628 VDD.n1315 VDD.n1160 4.5005
R83629 VDD.n1378 VDD.n1160 4.5005
R83630 VDD.n1313 VDD.n1160 4.5005
R83631 VDD.n1379 VDD.n1160 4.5005
R83632 VDD.n1312 VDD.n1160 4.5005
R83633 VDD.n1380 VDD.n1160 4.5005
R83634 VDD.n1310 VDD.n1160 4.5005
R83635 VDD.n1381 VDD.n1160 4.5005
R83636 VDD.n1309 VDD.n1160 4.5005
R83637 VDD.n1382 VDD.n1160 4.5005
R83638 VDD.n1307 VDD.n1160 4.5005
R83639 VDD.n1383 VDD.n1160 4.5005
R83640 VDD.n1306 VDD.n1160 4.5005
R83641 VDD.n1384 VDD.n1160 4.5005
R83642 VDD.n1304 VDD.n1160 4.5005
R83643 VDD.n1385 VDD.n1160 4.5005
R83644 VDD.n1303 VDD.n1160 4.5005
R83645 VDD.n1386 VDD.n1160 4.5005
R83646 VDD.n1301 VDD.n1160 4.5005
R83647 VDD.n1387 VDD.n1160 4.5005
R83648 VDD.n1300 VDD.n1160 4.5005
R83649 VDD.n1388 VDD.n1160 4.5005
R83650 VDD.n1298 VDD.n1160 4.5005
R83651 VDD.n1389 VDD.n1160 4.5005
R83652 VDD.n1297 VDD.n1160 4.5005
R83653 VDD.n1390 VDD.n1160 4.5005
R83654 VDD.n1295 VDD.n1160 4.5005
R83655 VDD.n1391 VDD.n1160 4.5005
R83656 VDD.n1294 VDD.n1160 4.5005
R83657 VDD.n1392 VDD.n1160 4.5005
R83658 VDD.n1292 VDD.n1160 4.5005
R83659 VDD.n1393 VDD.n1160 4.5005
R83660 VDD.n1291 VDD.n1160 4.5005
R83661 VDD.n1394 VDD.n1160 4.5005
R83662 VDD.n1289 VDD.n1160 4.5005
R83663 VDD.n1395 VDD.n1160 4.5005
R83664 VDD.n1288 VDD.n1160 4.5005
R83665 VDD.n1396 VDD.n1160 4.5005
R83666 VDD.n1286 VDD.n1160 4.5005
R83667 VDD.n1397 VDD.n1160 4.5005
R83668 VDD.n1285 VDD.n1160 4.5005
R83669 VDD.n1398 VDD.n1160 4.5005
R83670 VDD.n1283 VDD.n1160 4.5005
R83671 VDD.n1399 VDD.n1160 4.5005
R83672 VDD.n1282 VDD.n1160 4.5005
R83673 VDD.n1400 VDD.n1160 4.5005
R83674 VDD.n1280 VDD.n1160 4.5005
R83675 VDD.n1401 VDD.n1160 4.5005
R83676 VDD.n1279 VDD.n1160 4.5005
R83677 VDD.n1402 VDD.n1160 4.5005
R83678 VDD.n1277 VDD.n1160 4.5005
R83679 VDD.n1403 VDD.n1160 4.5005
R83680 VDD.n1276 VDD.n1160 4.5005
R83681 VDD.n1404 VDD.n1160 4.5005
R83682 VDD.n1274 VDD.n1160 4.5005
R83683 VDD.n1405 VDD.n1160 4.5005
R83684 VDD.n1273 VDD.n1160 4.5005
R83685 VDD.n1406 VDD.n1160 4.5005
R83686 VDD.n1271 VDD.n1160 4.5005
R83687 VDD.n1407 VDD.n1160 4.5005
R83688 VDD.n1270 VDD.n1160 4.5005
R83689 VDD.n1408 VDD.n1160 4.5005
R83690 VDD.n1268 VDD.n1160 4.5005
R83691 VDD.n1409 VDD.n1160 4.5005
R83692 VDD.n1267 VDD.n1160 4.5005
R83693 VDD.n1410 VDD.n1160 4.5005
R83694 VDD.n1265 VDD.n1160 4.5005
R83695 VDD.n1411 VDD.n1160 4.5005
R83696 VDD.n1264 VDD.n1160 4.5005
R83697 VDD.n1412 VDD.n1160 4.5005
R83698 VDD.n1262 VDD.n1160 4.5005
R83699 VDD.n1413 VDD.n1160 4.5005
R83700 VDD.n1261 VDD.n1160 4.5005
R83701 VDD.n1414 VDD.n1160 4.5005
R83702 VDD.n1415 VDD.n1160 4.5005
R83703 VDD.n1674 VDD.n1160 4.5005
R83704 VDD.n1676 VDD.n1230 4.5005
R83705 VDD.n1341 VDD.n1230 4.5005
R83706 VDD.n1342 VDD.n1230 4.5005
R83707 VDD.n1340 VDD.n1230 4.5005
R83708 VDD.n1344 VDD.n1230 4.5005
R83709 VDD.n1339 VDD.n1230 4.5005
R83710 VDD.n1345 VDD.n1230 4.5005
R83711 VDD.n1338 VDD.n1230 4.5005
R83712 VDD.n1347 VDD.n1230 4.5005
R83713 VDD.n1337 VDD.n1230 4.5005
R83714 VDD.n1348 VDD.n1230 4.5005
R83715 VDD.n1336 VDD.n1230 4.5005
R83716 VDD.n1350 VDD.n1230 4.5005
R83717 VDD.n1335 VDD.n1230 4.5005
R83718 VDD.n1351 VDD.n1230 4.5005
R83719 VDD.n1334 VDD.n1230 4.5005
R83720 VDD.n1353 VDD.n1230 4.5005
R83721 VDD.n1333 VDD.n1230 4.5005
R83722 VDD.n1354 VDD.n1230 4.5005
R83723 VDD.n1332 VDD.n1230 4.5005
R83724 VDD.n1356 VDD.n1230 4.5005
R83725 VDD.n1331 VDD.n1230 4.5005
R83726 VDD.n1357 VDD.n1230 4.5005
R83727 VDD.n1330 VDD.n1230 4.5005
R83728 VDD.n1359 VDD.n1230 4.5005
R83729 VDD.n1329 VDD.n1230 4.5005
R83730 VDD.n1360 VDD.n1230 4.5005
R83731 VDD.n1328 VDD.n1230 4.5005
R83732 VDD.n1362 VDD.n1230 4.5005
R83733 VDD.n1327 VDD.n1230 4.5005
R83734 VDD.n1363 VDD.n1230 4.5005
R83735 VDD.n1326 VDD.n1230 4.5005
R83736 VDD.n1365 VDD.n1230 4.5005
R83737 VDD.n1325 VDD.n1230 4.5005
R83738 VDD.n1366 VDD.n1230 4.5005
R83739 VDD.n1324 VDD.n1230 4.5005
R83740 VDD.n1368 VDD.n1230 4.5005
R83741 VDD.n1323 VDD.n1230 4.5005
R83742 VDD.n1369 VDD.n1230 4.5005
R83743 VDD.n1322 VDD.n1230 4.5005
R83744 VDD.n1371 VDD.n1230 4.5005
R83745 VDD.n1321 VDD.n1230 4.5005
R83746 VDD.n1372 VDD.n1230 4.5005
R83747 VDD.n1320 VDD.n1230 4.5005
R83748 VDD.n1374 VDD.n1230 4.5005
R83749 VDD.n1319 VDD.n1230 4.5005
R83750 VDD.n1375 VDD.n1230 4.5005
R83751 VDD.n1318 VDD.n1230 4.5005
R83752 VDD.n1376 VDD.n1230 4.5005
R83753 VDD.n1316 VDD.n1230 4.5005
R83754 VDD.n1377 VDD.n1230 4.5005
R83755 VDD.n1315 VDD.n1230 4.5005
R83756 VDD.n1378 VDD.n1230 4.5005
R83757 VDD.n1313 VDD.n1230 4.5005
R83758 VDD.n1379 VDD.n1230 4.5005
R83759 VDD.n1312 VDD.n1230 4.5005
R83760 VDD.n1380 VDD.n1230 4.5005
R83761 VDD.n1310 VDD.n1230 4.5005
R83762 VDD.n1381 VDD.n1230 4.5005
R83763 VDD.n1309 VDD.n1230 4.5005
R83764 VDD.n1382 VDD.n1230 4.5005
R83765 VDD.n1307 VDD.n1230 4.5005
R83766 VDD.n1383 VDD.n1230 4.5005
R83767 VDD.n1306 VDD.n1230 4.5005
R83768 VDD.n1384 VDD.n1230 4.5005
R83769 VDD.n1304 VDD.n1230 4.5005
R83770 VDD.n1385 VDD.n1230 4.5005
R83771 VDD.n1303 VDD.n1230 4.5005
R83772 VDD.n1386 VDD.n1230 4.5005
R83773 VDD.n1301 VDD.n1230 4.5005
R83774 VDD.n1387 VDD.n1230 4.5005
R83775 VDD.n1300 VDD.n1230 4.5005
R83776 VDD.n1388 VDD.n1230 4.5005
R83777 VDD.n1298 VDD.n1230 4.5005
R83778 VDD.n1389 VDD.n1230 4.5005
R83779 VDD.n1297 VDD.n1230 4.5005
R83780 VDD.n1390 VDD.n1230 4.5005
R83781 VDD.n1295 VDD.n1230 4.5005
R83782 VDD.n1391 VDD.n1230 4.5005
R83783 VDD.n1294 VDD.n1230 4.5005
R83784 VDD.n1392 VDD.n1230 4.5005
R83785 VDD.n1292 VDD.n1230 4.5005
R83786 VDD.n1393 VDD.n1230 4.5005
R83787 VDD.n1291 VDD.n1230 4.5005
R83788 VDD.n1394 VDD.n1230 4.5005
R83789 VDD.n1289 VDD.n1230 4.5005
R83790 VDD.n1395 VDD.n1230 4.5005
R83791 VDD.n1288 VDD.n1230 4.5005
R83792 VDD.n1396 VDD.n1230 4.5005
R83793 VDD.n1286 VDD.n1230 4.5005
R83794 VDD.n1397 VDD.n1230 4.5005
R83795 VDD.n1285 VDD.n1230 4.5005
R83796 VDD.n1398 VDD.n1230 4.5005
R83797 VDD.n1283 VDD.n1230 4.5005
R83798 VDD.n1399 VDD.n1230 4.5005
R83799 VDD.n1282 VDD.n1230 4.5005
R83800 VDD.n1400 VDD.n1230 4.5005
R83801 VDD.n1280 VDD.n1230 4.5005
R83802 VDD.n1401 VDD.n1230 4.5005
R83803 VDD.n1279 VDD.n1230 4.5005
R83804 VDD.n1402 VDD.n1230 4.5005
R83805 VDD.n1277 VDD.n1230 4.5005
R83806 VDD.n1403 VDD.n1230 4.5005
R83807 VDD.n1276 VDD.n1230 4.5005
R83808 VDD.n1404 VDD.n1230 4.5005
R83809 VDD.n1274 VDD.n1230 4.5005
R83810 VDD.n1405 VDD.n1230 4.5005
R83811 VDD.n1273 VDD.n1230 4.5005
R83812 VDD.n1406 VDD.n1230 4.5005
R83813 VDD.n1271 VDD.n1230 4.5005
R83814 VDD.n1407 VDD.n1230 4.5005
R83815 VDD.n1270 VDD.n1230 4.5005
R83816 VDD.n1408 VDD.n1230 4.5005
R83817 VDD.n1268 VDD.n1230 4.5005
R83818 VDD.n1409 VDD.n1230 4.5005
R83819 VDD.n1267 VDD.n1230 4.5005
R83820 VDD.n1410 VDD.n1230 4.5005
R83821 VDD.n1265 VDD.n1230 4.5005
R83822 VDD.n1411 VDD.n1230 4.5005
R83823 VDD.n1264 VDD.n1230 4.5005
R83824 VDD.n1412 VDD.n1230 4.5005
R83825 VDD.n1262 VDD.n1230 4.5005
R83826 VDD.n1413 VDD.n1230 4.5005
R83827 VDD.n1261 VDD.n1230 4.5005
R83828 VDD.n1414 VDD.n1230 4.5005
R83829 VDD.n1415 VDD.n1230 4.5005
R83830 VDD.n1674 VDD.n1230 4.5005
R83831 VDD.n1676 VDD.n1159 4.5005
R83832 VDD.n1341 VDD.n1159 4.5005
R83833 VDD.n1342 VDD.n1159 4.5005
R83834 VDD.n1340 VDD.n1159 4.5005
R83835 VDD.n1344 VDD.n1159 4.5005
R83836 VDD.n1339 VDD.n1159 4.5005
R83837 VDD.n1345 VDD.n1159 4.5005
R83838 VDD.n1338 VDD.n1159 4.5005
R83839 VDD.n1347 VDD.n1159 4.5005
R83840 VDD.n1337 VDD.n1159 4.5005
R83841 VDD.n1348 VDD.n1159 4.5005
R83842 VDD.n1336 VDD.n1159 4.5005
R83843 VDD.n1350 VDD.n1159 4.5005
R83844 VDD.n1335 VDD.n1159 4.5005
R83845 VDD.n1351 VDD.n1159 4.5005
R83846 VDD.n1334 VDD.n1159 4.5005
R83847 VDD.n1353 VDD.n1159 4.5005
R83848 VDD.n1333 VDD.n1159 4.5005
R83849 VDD.n1354 VDD.n1159 4.5005
R83850 VDD.n1332 VDD.n1159 4.5005
R83851 VDD.n1356 VDD.n1159 4.5005
R83852 VDD.n1331 VDD.n1159 4.5005
R83853 VDD.n1357 VDD.n1159 4.5005
R83854 VDD.n1330 VDD.n1159 4.5005
R83855 VDD.n1359 VDD.n1159 4.5005
R83856 VDD.n1329 VDD.n1159 4.5005
R83857 VDD.n1360 VDD.n1159 4.5005
R83858 VDD.n1328 VDD.n1159 4.5005
R83859 VDD.n1362 VDD.n1159 4.5005
R83860 VDD.n1327 VDD.n1159 4.5005
R83861 VDD.n1363 VDD.n1159 4.5005
R83862 VDD.n1326 VDD.n1159 4.5005
R83863 VDD.n1365 VDD.n1159 4.5005
R83864 VDD.n1325 VDD.n1159 4.5005
R83865 VDD.n1366 VDD.n1159 4.5005
R83866 VDD.n1324 VDD.n1159 4.5005
R83867 VDD.n1368 VDD.n1159 4.5005
R83868 VDD.n1323 VDD.n1159 4.5005
R83869 VDD.n1369 VDD.n1159 4.5005
R83870 VDD.n1322 VDD.n1159 4.5005
R83871 VDD.n1371 VDD.n1159 4.5005
R83872 VDD.n1321 VDD.n1159 4.5005
R83873 VDD.n1372 VDD.n1159 4.5005
R83874 VDD.n1320 VDD.n1159 4.5005
R83875 VDD.n1374 VDD.n1159 4.5005
R83876 VDD.n1319 VDD.n1159 4.5005
R83877 VDD.n1375 VDD.n1159 4.5005
R83878 VDD.n1318 VDD.n1159 4.5005
R83879 VDD.n1376 VDD.n1159 4.5005
R83880 VDD.n1316 VDD.n1159 4.5005
R83881 VDD.n1377 VDD.n1159 4.5005
R83882 VDD.n1315 VDD.n1159 4.5005
R83883 VDD.n1378 VDD.n1159 4.5005
R83884 VDD.n1313 VDD.n1159 4.5005
R83885 VDD.n1379 VDD.n1159 4.5005
R83886 VDD.n1312 VDD.n1159 4.5005
R83887 VDD.n1380 VDD.n1159 4.5005
R83888 VDD.n1310 VDD.n1159 4.5005
R83889 VDD.n1381 VDD.n1159 4.5005
R83890 VDD.n1309 VDD.n1159 4.5005
R83891 VDD.n1382 VDD.n1159 4.5005
R83892 VDD.n1307 VDD.n1159 4.5005
R83893 VDD.n1383 VDD.n1159 4.5005
R83894 VDD.n1306 VDD.n1159 4.5005
R83895 VDD.n1384 VDD.n1159 4.5005
R83896 VDD.n1304 VDD.n1159 4.5005
R83897 VDD.n1385 VDD.n1159 4.5005
R83898 VDD.n1303 VDD.n1159 4.5005
R83899 VDD.n1386 VDD.n1159 4.5005
R83900 VDD.n1301 VDD.n1159 4.5005
R83901 VDD.n1387 VDD.n1159 4.5005
R83902 VDD.n1300 VDD.n1159 4.5005
R83903 VDD.n1388 VDD.n1159 4.5005
R83904 VDD.n1298 VDD.n1159 4.5005
R83905 VDD.n1389 VDD.n1159 4.5005
R83906 VDD.n1297 VDD.n1159 4.5005
R83907 VDD.n1390 VDD.n1159 4.5005
R83908 VDD.n1295 VDD.n1159 4.5005
R83909 VDD.n1391 VDD.n1159 4.5005
R83910 VDD.n1294 VDD.n1159 4.5005
R83911 VDD.n1392 VDD.n1159 4.5005
R83912 VDD.n1292 VDD.n1159 4.5005
R83913 VDD.n1393 VDD.n1159 4.5005
R83914 VDD.n1291 VDD.n1159 4.5005
R83915 VDD.n1394 VDD.n1159 4.5005
R83916 VDD.n1289 VDD.n1159 4.5005
R83917 VDD.n1395 VDD.n1159 4.5005
R83918 VDD.n1288 VDD.n1159 4.5005
R83919 VDD.n1396 VDD.n1159 4.5005
R83920 VDD.n1286 VDD.n1159 4.5005
R83921 VDD.n1397 VDD.n1159 4.5005
R83922 VDD.n1285 VDD.n1159 4.5005
R83923 VDD.n1398 VDD.n1159 4.5005
R83924 VDD.n1283 VDD.n1159 4.5005
R83925 VDD.n1399 VDD.n1159 4.5005
R83926 VDD.n1282 VDD.n1159 4.5005
R83927 VDD.n1400 VDD.n1159 4.5005
R83928 VDD.n1280 VDD.n1159 4.5005
R83929 VDD.n1401 VDD.n1159 4.5005
R83930 VDD.n1279 VDD.n1159 4.5005
R83931 VDD.n1402 VDD.n1159 4.5005
R83932 VDD.n1277 VDD.n1159 4.5005
R83933 VDD.n1403 VDD.n1159 4.5005
R83934 VDD.n1276 VDD.n1159 4.5005
R83935 VDD.n1404 VDD.n1159 4.5005
R83936 VDD.n1274 VDD.n1159 4.5005
R83937 VDD.n1405 VDD.n1159 4.5005
R83938 VDD.n1273 VDD.n1159 4.5005
R83939 VDD.n1406 VDD.n1159 4.5005
R83940 VDD.n1271 VDD.n1159 4.5005
R83941 VDD.n1407 VDD.n1159 4.5005
R83942 VDD.n1270 VDD.n1159 4.5005
R83943 VDD.n1408 VDD.n1159 4.5005
R83944 VDD.n1268 VDD.n1159 4.5005
R83945 VDD.n1409 VDD.n1159 4.5005
R83946 VDD.n1267 VDD.n1159 4.5005
R83947 VDD.n1410 VDD.n1159 4.5005
R83948 VDD.n1265 VDD.n1159 4.5005
R83949 VDD.n1411 VDD.n1159 4.5005
R83950 VDD.n1264 VDD.n1159 4.5005
R83951 VDD.n1412 VDD.n1159 4.5005
R83952 VDD.n1262 VDD.n1159 4.5005
R83953 VDD.n1413 VDD.n1159 4.5005
R83954 VDD.n1261 VDD.n1159 4.5005
R83955 VDD.n1414 VDD.n1159 4.5005
R83956 VDD.n1415 VDD.n1159 4.5005
R83957 VDD.n1674 VDD.n1159 4.5005
R83958 VDD.n1676 VDD.n1231 4.5005
R83959 VDD.n1341 VDD.n1231 4.5005
R83960 VDD.n1342 VDD.n1231 4.5005
R83961 VDD.n1340 VDD.n1231 4.5005
R83962 VDD.n1344 VDD.n1231 4.5005
R83963 VDD.n1339 VDD.n1231 4.5005
R83964 VDD.n1345 VDD.n1231 4.5005
R83965 VDD.n1338 VDD.n1231 4.5005
R83966 VDD.n1347 VDD.n1231 4.5005
R83967 VDD.n1337 VDD.n1231 4.5005
R83968 VDD.n1348 VDD.n1231 4.5005
R83969 VDD.n1336 VDD.n1231 4.5005
R83970 VDD.n1350 VDD.n1231 4.5005
R83971 VDD.n1335 VDD.n1231 4.5005
R83972 VDD.n1351 VDD.n1231 4.5005
R83973 VDD.n1334 VDD.n1231 4.5005
R83974 VDD.n1353 VDD.n1231 4.5005
R83975 VDD.n1333 VDD.n1231 4.5005
R83976 VDD.n1354 VDD.n1231 4.5005
R83977 VDD.n1332 VDD.n1231 4.5005
R83978 VDD.n1356 VDD.n1231 4.5005
R83979 VDD.n1331 VDD.n1231 4.5005
R83980 VDD.n1357 VDD.n1231 4.5005
R83981 VDD.n1330 VDD.n1231 4.5005
R83982 VDD.n1359 VDD.n1231 4.5005
R83983 VDD.n1329 VDD.n1231 4.5005
R83984 VDD.n1360 VDD.n1231 4.5005
R83985 VDD.n1328 VDD.n1231 4.5005
R83986 VDD.n1362 VDD.n1231 4.5005
R83987 VDD.n1327 VDD.n1231 4.5005
R83988 VDD.n1363 VDD.n1231 4.5005
R83989 VDD.n1326 VDD.n1231 4.5005
R83990 VDD.n1365 VDD.n1231 4.5005
R83991 VDD.n1325 VDD.n1231 4.5005
R83992 VDD.n1366 VDD.n1231 4.5005
R83993 VDD.n1324 VDD.n1231 4.5005
R83994 VDD.n1368 VDD.n1231 4.5005
R83995 VDD.n1323 VDD.n1231 4.5005
R83996 VDD.n1369 VDD.n1231 4.5005
R83997 VDD.n1322 VDD.n1231 4.5005
R83998 VDD.n1371 VDD.n1231 4.5005
R83999 VDD.n1321 VDD.n1231 4.5005
R84000 VDD.n1372 VDD.n1231 4.5005
R84001 VDD.n1320 VDD.n1231 4.5005
R84002 VDD.n1374 VDD.n1231 4.5005
R84003 VDD.n1319 VDD.n1231 4.5005
R84004 VDD.n1375 VDD.n1231 4.5005
R84005 VDD.n1318 VDD.n1231 4.5005
R84006 VDD.n1376 VDD.n1231 4.5005
R84007 VDD.n1316 VDD.n1231 4.5005
R84008 VDD.n1377 VDD.n1231 4.5005
R84009 VDD.n1315 VDD.n1231 4.5005
R84010 VDD.n1378 VDD.n1231 4.5005
R84011 VDD.n1313 VDD.n1231 4.5005
R84012 VDD.n1379 VDD.n1231 4.5005
R84013 VDD.n1312 VDD.n1231 4.5005
R84014 VDD.n1380 VDD.n1231 4.5005
R84015 VDD.n1310 VDD.n1231 4.5005
R84016 VDD.n1381 VDD.n1231 4.5005
R84017 VDD.n1309 VDD.n1231 4.5005
R84018 VDD.n1382 VDD.n1231 4.5005
R84019 VDD.n1307 VDD.n1231 4.5005
R84020 VDD.n1383 VDD.n1231 4.5005
R84021 VDD.n1306 VDD.n1231 4.5005
R84022 VDD.n1384 VDD.n1231 4.5005
R84023 VDD.n1304 VDD.n1231 4.5005
R84024 VDD.n1385 VDD.n1231 4.5005
R84025 VDD.n1303 VDD.n1231 4.5005
R84026 VDD.n1386 VDD.n1231 4.5005
R84027 VDD.n1301 VDD.n1231 4.5005
R84028 VDD.n1387 VDD.n1231 4.5005
R84029 VDD.n1300 VDD.n1231 4.5005
R84030 VDD.n1388 VDD.n1231 4.5005
R84031 VDD.n1298 VDD.n1231 4.5005
R84032 VDD.n1389 VDD.n1231 4.5005
R84033 VDD.n1297 VDD.n1231 4.5005
R84034 VDD.n1390 VDD.n1231 4.5005
R84035 VDD.n1295 VDD.n1231 4.5005
R84036 VDD.n1391 VDD.n1231 4.5005
R84037 VDD.n1294 VDD.n1231 4.5005
R84038 VDD.n1392 VDD.n1231 4.5005
R84039 VDD.n1292 VDD.n1231 4.5005
R84040 VDD.n1393 VDD.n1231 4.5005
R84041 VDD.n1291 VDD.n1231 4.5005
R84042 VDD.n1394 VDD.n1231 4.5005
R84043 VDD.n1289 VDD.n1231 4.5005
R84044 VDD.n1395 VDD.n1231 4.5005
R84045 VDD.n1288 VDD.n1231 4.5005
R84046 VDD.n1396 VDD.n1231 4.5005
R84047 VDD.n1286 VDD.n1231 4.5005
R84048 VDD.n1397 VDD.n1231 4.5005
R84049 VDD.n1285 VDD.n1231 4.5005
R84050 VDD.n1398 VDD.n1231 4.5005
R84051 VDD.n1283 VDD.n1231 4.5005
R84052 VDD.n1399 VDD.n1231 4.5005
R84053 VDD.n1282 VDD.n1231 4.5005
R84054 VDD.n1400 VDD.n1231 4.5005
R84055 VDD.n1280 VDD.n1231 4.5005
R84056 VDD.n1401 VDD.n1231 4.5005
R84057 VDD.n1279 VDD.n1231 4.5005
R84058 VDD.n1402 VDD.n1231 4.5005
R84059 VDD.n1277 VDD.n1231 4.5005
R84060 VDD.n1403 VDD.n1231 4.5005
R84061 VDD.n1276 VDD.n1231 4.5005
R84062 VDD.n1404 VDD.n1231 4.5005
R84063 VDD.n1274 VDD.n1231 4.5005
R84064 VDD.n1405 VDD.n1231 4.5005
R84065 VDD.n1273 VDD.n1231 4.5005
R84066 VDD.n1406 VDD.n1231 4.5005
R84067 VDD.n1271 VDD.n1231 4.5005
R84068 VDD.n1407 VDD.n1231 4.5005
R84069 VDD.n1270 VDD.n1231 4.5005
R84070 VDD.n1408 VDD.n1231 4.5005
R84071 VDD.n1268 VDD.n1231 4.5005
R84072 VDD.n1409 VDD.n1231 4.5005
R84073 VDD.n1267 VDD.n1231 4.5005
R84074 VDD.n1410 VDD.n1231 4.5005
R84075 VDD.n1265 VDD.n1231 4.5005
R84076 VDD.n1411 VDD.n1231 4.5005
R84077 VDD.n1264 VDD.n1231 4.5005
R84078 VDD.n1412 VDD.n1231 4.5005
R84079 VDD.n1262 VDD.n1231 4.5005
R84080 VDD.n1413 VDD.n1231 4.5005
R84081 VDD.n1261 VDD.n1231 4.5005
R84082 VDD.n1414 VDD.n1231 4.5005
R84083 VDD.n1415 VDD.n1231 4.5005
R84084 VDD.n1674 VDD.n1231 4.5005
R84085 VDD.n1676 VDD.n1158 4.5005
R84086 VDD.n1341 VDD.n1158 4.5005
R84087 VDD.n1342 VDD.n1158 4.5005
R84088 VDD.n1340 VDD.n1158 4.5005
R84089 VDD.n1344 VDD.n1158 4.5005
R84090 VDD.n1339 VDD.n1158 4.5005
R84091 VDD.n1345 VDD.n1158 4.5005
R84092 VDD.n1338 VDD.n1158 4.5005
R84093 VDD.n1347 VDD.n1158 4.5005
R84094 VDD.n1337 VDD.n1158 4.5005
R84095 VDD.n1348 VDD.n1158 4.5005
R84096 VDD.n1336 VDD.n1158 4.5005
R84097 VDD.n1350 VDD.n1158 4.5005
R84098 VDD.n1335 VDD.n1158 4.5005
R84099 VDD.n1351 VDD.n1158 4.5005
R84100 VDD.n1334 VDD.n1158 4.5005
R84101 VDD.n1353 VDD.n1158 4.5005
R84102 VDD.n1333 VDD.n1158 4.5005
R84103 VDD.n1354 VDD.n1158 4.5005
R84104 VDD.n1332 VDD.n1158 4.5005
R84105 VDD.n1356 VDD.n1158 4.5005
R84106 VDD.n1331 VDD.n1158 4.5005
R84107 VDD.n1357 VDD.n1158 4.5005
R84108 VDD.n1330 VDD.n1158 4.5005
R84109 VDD.n1359 VDD.n1158 4.5005
R84110 VDD.n1329 VDD.n1158 4.5005
R84111 VDD.n1360 VDD.n1158 4.5005
R84112 VDD.n1328 VDD.n1158 4.5005
R84113 VDD.n1362 VDD.n1158 4.5005
R84114 VDD.n1327 VDD.n1158 4.5005
R84115 VDD.n1363 VDD.n1158 4.5005
R84116 VDD.n1326 VDD.n1158 4.5005
R84117 VDD.n1365 VDD.n1158 4.5005
R84118 VDD.n1325 VDD.n1158 4.5005
R84119 VDD.n1366 VDD.n1158 4.5005
R84120 VDD.n1324 VDD.n1158 4.5005
R84121 VDD.n1368 VDD.n1158 4.5005
R84122 VDD.n1323 VDD.n1158 4.5005
R84123 VDD.n1369 VDD.n1158 4.5005
R84124 VDD.n1322 VDD.n1158 4.5005
R84125 VDD.n1371 VDD.n1158 4.5005
R84126 VDD.n1321 VDD.n1158 4.5005
R84127 VDD.n1372 VDD.n1158 4.5005
R84128 VDD.n1320 VDD.n1158 4.5005
R84129 VDD.n1374 VDD.n1158 4.5005
R84130 VDD.n1319 VDD.n1158 4.5005
R84131 VDD.n1375 VDD.n1158 4.5005
R84132 VDD.n1318 VDD.n1158 4.5005
R84133 VDD.n1376 VDD.n1158 4.5005
R84134 VDD.n1316 VDD.n1158 4.5005
R84135 VDD.n1377 VDD.n1158 4.5005
R84136 VDD.n1315 VDD.n1158 4.5005
R84137 VDD.n1378 VDD.n1158 4.5005
R84138 VDD.n1313 VDD.n1158 4.5005
R84139 VDD.n1379 VDD.n1158 4.5005
R84140 VDD.n1312 VDD.n1158 4.5005
R84141 VDD.n1380 VDD.n1158 4.5005
R84142 VDD.n1310 VDD.n1158 4.5005
R84143 VDD.n1381 VDD.n1158 4.5005
R84144 VDD.n1309 VDD.n1158 4.5005
R84145 VDD.n1382 VDD.n1158 4.5005
R84146 VDD.n1307 VDD.n1158 4.5005
R84147 VDD.n1383 VDD.n1158 4.5005
R84148 VDD.n1306 VDD.n1158 4.5005
R84149 VDD.n1384 VDD.n1158 4.5005
R84150 VDD.n1304 VDD.n1158 4.5005
R84151 VDD.n1385 VDD.n1158 4.5005
R84152 VDD.n1303 VDD.n1158 4.5005
R84153 VDD.n1386 VDD.n1158 4.5005
R84154 VDD.n1301 VDD.n1158 4.5005
R84155 VDD.n1387 VDD.n1158 4.5005
R84156 VDD.n1300 VDD.n1158 4.5005
R84157 VDD.n1388 VDD.n1158 4.5005
R84158 VDD.n1298 VDD.n1158 4.5005
R84159 VDD.n1389 VDD.n1158 4.5005
R84160 VDD.n1297 VDD.n1158 4.5005
R84161 VDD.n1390 VDD.n1158 4.5005
R84162 VDD.n1295 VDD.n1158 4.5005
R84163 VDD.n1391 VDD.n1158 4.5005
R84164 VDD.n1294 VDD.n1158 4.5005
R84165 VDD.n1392 VDD.n1158 4.5005
R84166 VDD.n1292 VDD.n1158 4.5005
R84167 VDD.n1393 VDD.n1158 4.5005
R84168 VDD.n1291 VDD.n1158 4.5005
R84169 VDD.n1394 VDD.n1158 4.5005
R84170 VDD.n1289 VDD.n1158 4.5005
R84171 VDD.n1395 VDD.n1158 4.5005
R84172 VDD.n1288 VDD.n1158 4.5005
R84173 VDD.n1396 VDD.n1158 4.5005
R84174 VDD.n1286 VDD.n1158 4.5005
R84175 VDD.n1397 VDD.n1158 4.5005
R84176 VDD.n1285 VDD.n1158 4.5005
R84177 VDD.n1398 VDD.n1158 4.5005
R84178 VDD.n1283 VDD.n1158 4.5005
R84179 VDD.n1399 VDD.n1158 4.5005
R84180 VDD.n1282 VDD.n1158 4.5005
R84181 VDD.n1400 VDD.n1158 4.5005
R84182 VDD.n1280 VDD.n1158 4.5005
R84183 VDD.n1401 VDD.n1158 4.5005
R84184 VDD.n1279 VDD.n1158 4.5005
R84185 VDD.n1402 VDD.n1158 4.5005
R84186 VDD.n1277 VDD.n1158 4.5005
R84187 VDD.n1403 VDD.n1158 4.5005
R84188 VDD.n1276 VDD.n1158 4.5005
R84189 VDD.n1404 VDD.n1158 4.5005
R84190 VDD.n1274 VDD.n1158 4.5005
R84191 VDD.n1405 VDD.n1158 4.5005
R84192 VDD.n1273 VDD.n1158 4.5005
R84193 VDD.n1406 VDD.n1158 4.5005
R84194 VDD.n1271 VDD.n1158 4.5005
R84195 VDD.n1407 VDD.n1158 4.5005
R84196 VDD.n1270 VDD.n1158 4.5005
R84197 VDD.n1408 VDD.n1158 4.5005
R84198 VDD.n1268 VDD.n1158 4.5005
R84199 VDD.n1409 VDD.n1158 4.5005
R84200 VDD.n1267 VDD.n1158 4.5005
R84201 VDD.n1410 VDD.n1158 4.5005
R84202 VDD.n1265 VDD.n1158 4.5005
R84203 VDD.n1411 VDD.n1158 4.5005
R84204 VDD.n1264 VDD.n1158 4.5005
R84205 VDD.n1412 VDD.n1158 4.5005
R84206 VDD.n1262 VDD.n1158 4.5005
R84207 VDD.n1413 VDD.n1158 4.5005
R84208 VDD.n1261 VDD.n1158 4.5005
R84209 VDD.n1414 VDD.n1158 4.5005
R84210 VDD.n1415 VDD.n1158 4.5005
R84211 VDD.n1674 VDD.n1158 4.5005
R84212 VDD.n1676 VDD.n1232 4.5005
R84213 VDD.n1341 VDD.n1232 4.5005
R84214 VDD.n1342 VDD.n1232 4.5005
R84215 VDD.n1340 VDD.n1232 4.5005
R84216 VDD.n1344 VDD.n1232 4.5005
R84217 VDD.n1339 VDD.n1232 4.5005
R84218 VDD.n1345 VDD.n1232 4.5005
R84219 VDD.n1338 VDD.n1232 4.5005
R84220 VDD.n1347 VDD.n1232 4.5005
R84221 VDD.n1337 VDD.n1232 4.5005
R84222 VDD.n1348 VDD.n1232 4.5005
R84223 VDD.n1336 VDD.n1232 4.5005
R84224 VDD.n1350 VDD.n1232 4.5005
R84225 VDD.n1335 VDD.n1232 4.5005
R84226 VDD.n1351 VDD.n1232 4.5005
R84227 VDD.n1334 VDD.n1232 4.5005
R84228 VDD.n1353 VDD.n1232 4.5005
R84229 VDD.n1333 VDD.n1232 4.5005
R84230 VDD.n1354 VDD.n1232 4.5005
R84231 VDD.n1332 VDD.n1232 4.5005
R84232 VDD.n1356 VDD.n1232 4.5005
R84233 VDD.n1331 VDD.n1232 4.5005
R84234 VDD.n1357 VDD.n1232 4.5005
R84235 VDD.n1330 VDD.n1232 4.5005
R84236 VDD.n1359 VDD.n1232 4.5005
R84237 VDD.n1329 VDD.n1232 4.5005
R84238 VDD.n1360 VDD.n1232 4.5005
R84239 VDD.n1328 VDD.n1232 4.5005
R84240 VDD.n1362 VDD.n1232 4.5005
R84241 VDD.n1327 VDD.n1232 4.5005
R84242 VDD.n1363 VDD.n1232 4.5005
R84243 VDD.n1326 VDD.n1232 4.5005
R84244 VDD.n1365 VDD.n1232 4.5005
R84245 VDD.n1325 VDD.n1232 4.5005
R84246 VDD.n1366 VDD.n1232 4.5005
R84247 VDD.n1324 VDD.n1232 4.5005
R84248 VDD.n1368 VDD.n1232 4.5005
R84249 VDD.n1323 VDD.n1232 4.5005
R84250 VDD.n1369 VDD.n1232 4.5005
R84251 VDD.n1322 VDD.n1232 4.5005
R84252 VDD.n1371 VDD.n1232 4.5005
R84253 VDD.n1321 VDD.n1232 4.5005
R84254 VDD.n1372 VDD.n1232 4.5005
R84255 VDD.n1320 VDD.n1232 4.5005
R84256 VDD.n1374 VDD.n1232 4.5005
R84257 VDD.n1319 VDD.n1232 4.5005
R84258 VDD.n1375 VDD.n1232 4.5005
R84259 VDD.n1318 VDD.n1232 4.5005
R84260 VDD.n1376 VDD.n1232 4.5005
R84261 VDD.n1316 VDD.n1232 4.5005
R84262 VDD.n1377 VDD.n1232 4.5005
R84263 VDD.n1315 VDD.n1232 4.5005
R84264 VDD.n1378 VDD.n1232 4.5005
R84265 VDD.n1313 VDD.n1232 4.5005
R84266 VDD.n1379 VDD.n1232 4.5005
R84267 VDD.n1312 VDD.n1232 4.5005
R84268 VDD.n1380 VDD.n1232 4.5005
R84269 VDD.n1310 VDD.n1232 4.5005
R84270 VDD.n1381 VDD.n1232 4.5005
R84271 VDD.n1309 VDD.n1232 4.5005
R84272 VDD.n1382 VDD.n1232 4.5005
R84273 VDD.n1307 VDD.n1232 4.5005
R84274 VDD.n1383 VDD.n1232 4.5005
R84275 VDD.n1306 VDD.n1232 4.5005
R84276 VDD.n1384 VDD.n1232 4.5005
R84277 VDD.n1304 VDD.n1232 4.5005
R84278 VDD.n1385 VDD.n1232 4.5005
R84279 VDD.n1303 VDD.n1232 4.5005
R84280 VDD.n1386 VDD.n1232 4.5005
R84281 VDD.n1301 VDD.n1232 4.5005
R84282 VDD.n1387 VDD.n1232 4.5005
R84283 VDD.n1300 VDD.n1232 4.5005
R84284 VDD.n1388 VDD.n1232 4.5005
R84285 VDD.n1298 VDD.n1232 4.5005
R84286 VDD.n1389 VDD.n1232 4.5005
R84287 VDD.n1297 VDD.n1232 4.5005
R84288 VDD.n1390 VDD.n1232 4.5005
R84289 VDD.n1295 VDD.n1232 4.5005
R84290 VDD.n1391 VDD.n1232 4.5005
R84291 VDD.n1294 VDD.n1232 4.5005
R84292 VDD.n1392 VDD.n1232 4.5005
R84293 VDD.n1292 VDD.n1232 4.5005
R84294 VDD.n1393 VDD.n1232 4.5005
R84295 VDD.n1291 VDD.n1232 4.5005
R84296 VDD.n1394 VDD.n1232 4.5005
R84297 VDD.n1289 VDD.n1232 4.5005
R84298 VDD.n1395 VDD.n1232 4.5005
R84299 VDD.n1288 VDD.n1232 4.5005
R84300 VDD.n1396 VDD.n1232 4.5005
R84301 VDD.n1286 VDD.n1232 4.5005
R84302 VDD.n1397 VDD.n1232 4.5005
R84303 VDD.n1285 VDD.n1232 4.5005
R84304 VDD.n1398 VDD.n1232 4.5005
R84305 VDD.n1283 VDD.n1232 4.5005
R84306 VDD.n1399 VDD.n1232 4.5005
R84307 VDD.n1282 VDD.n1232 4.5005
R84308 VDD.n1400 VDD.n1232 4.5005
R84309 VDD.n1280 VDD.n1232 4.5005
R84310 VDD.n1401 VDD.n1232 4.5005
R84311 VDD.n1279 VDD.n1232 4.5005
R84312 VDD.n1402 VDD.n1232 4.5005
R84313 VDD.n1277 VDD.n1232 4.5005
R84314 VDD.n1403 VDD.n1232 4.5005
R84315 VDD.n1276 VDD.n1232 4.5005
R84316 VDD.n1404 VDD.n1232 4.5005
R84317 VDD.n1274 VDD.n1232 4.5005
R84318 VDD.n1405 VDD.n1232 4.5005
R84319 VDD.n1273 VDD.n1232 4.5005
R84320 VDD.n1406 VDD.n1232 4.5005
R84321 VDD.n1271 VDD.n1232 4.5005
R84322 VDD.n1407 VDD.n1232 4.5005
R84323 VDD.n1270 VDD.n1232 4.5005
R84324 VDD.n1408 VDD.n1232 4.5005
R84325 VDD.n1268 VDD.n1232 4.5005
R84326 VDD.n1409 VDD.n1232 4.5005
R84327 VDD.n1267 VDD.n1232 4.5005
R84328 VDD.n1410 VDD.n1232 4.5005
R84329 VDD.n1265 VDD.n1232 4.5005
R84330 VDD.n1411 VDD.n1232 4.5005
R84331 VDD.n1264 VDD.n1232 4.5005
R84332 VDD.n1412 VDD.n1232 4.5005
R84333 VDD.n1262 VDD.n1232 4.5005
R84334 VDD.n1413 VDD.n1232 4.5005
R84335 VDD.n1261 VDD.n1232 4.5005
R84336 VDD.n1414 VDD.n1232 4.5005
R84337 VDD.n1415 VDD.n1232 4.5005
R84338 VDD.n1674 VDD.n1232 4.5005
R84339 VDD.n1676 VDD.n1157 4.5005
R84340 VDD.n1341 VDD.n1157 4.5005
R84341 VDD.n1342 VDD.n1157 4.5005
R84342 VDD.n1340 VDD.n1157 4.5005
R84343 VDD.n1344 VDD.n1157 4.5005
R84344 VDD.n1339 VDD.n1157 4.5005
R84345 VDD.n1345 VDD.n1157 4.5005
R84346 VDD.n1338 VDD.n1157 4.5005
R84347 VDD.n1347 VDD.n1157 4.5005
R84348 VDD.n1337 VDD.n1157 4.5005
R84349 VDD.n1348 VDD.n1157 4.5005
R84350 VDD.n1336 VDD.n1157 4.5005
R84351 VDD.n1350 VDD.n1157 4.5005
R84352 VDD.n1335 VDD.n1157 4.5005
R84353 VDD.n1351 VDD.n1157 4.5005
R84354 VDD.n1334 VDD.n1157 4.5005
R84355 VDD.n1353 VDD.n1157 4.5005
R84356 VDD.n1333 VDD.n1157 4.5005
R84357 VDD.n1354 VDD.n1157 4.5005
R84358 VDD.n1332 VDD.n1157 4.5005
R84359 VDD.n1356 VDD.n1157 4.5005
R84360 VDD.n1331 VDD.n1157 4.5005
R84361 VDD.n1357 VDD.n1157 4.5005
R84362 VDD.n1330 VDD.n1157 4.5005
R84363 VDD.n1359 VDD.n1157 4.5005
R84364 VDD.n1329 VDD.n1157 4.5005
R84365 VDD.n1360 VDD.n1157 4.5005
R84366 VDD.n1328 VDD.n1157 4.5005
R84367 VDD.n1362 VDD.n1157 4.5005
R84368 VDD.n1327 VDD.n1157 4.5005
R84369 VDD.n1363 VDD.n1157 4.5005
R84370 VDD.n1326 VDD.n1157 4.5005
R84371 VDD.n1365 VDD.n1157 4.5005
R84372 VDD.n1325 VDD.n1157 4.5005
R84373 VDD.n1366 VDD.n1157 4.5005
R84374 VDD.n1324 VDD.n1157 4.5005
R84375 VDD.n1368 VDD.n1157 4.5005
R84376 VDD.n1323 VDD.n1157 4.5005
R84377 VDD.n1369 VDD.n1157 4.5005
R84378 VDD.n1322 VDD.n1157 4.5005
R84379 VDD.n1371 VDD.n1157 4.5005
R84380 VDD.n1321 VDD.n1157 4.5005
R84381 VDD.n1372 VDD.n1157 4.5005
R84382 VDD.n1320 VDD.n1157 4.5005
R84383 VDD.n1374 VDD.n1157 4.5005
R84384 VDD.n1319 VDD.n1157 4.5005
R84385 VDD.n1375 VDD.n1157 4.5005
R84386 VDD.n1318 VDD.n1157 4.5005
R84387 VDD.n1376 VDD.n1157 4.5005
R84388 VDD.n1316 VDD.n1157 4.5005
R84389 VDD.n1377 VDD.n1157 4.5005
R84390 VDD.n1315 VDD.n1157 4.5005
R84391 VDD.n1378 VDD.n1157 4.5005
R84392 VDD.n1313 VDD.n1157 4.5005
R84393 VDD.n1379 VDD.n1157 4.5005
R84394 VDD.n1312 VDD.n1157 4.5005
R84395 VDD.n1380 VDD.n1157 4.5005
R84396 VDD.n1310 VDD.n1157 4.5005
R84397 VDD.n1381 VDD.n1157 4.5005
R84398 VDD.n1309 VDD.n1157 4.5005
R84399 VDD.n1382 VDD.n1157 4.5005
R84400 VDD.n1307 VDD.n1157 4.5005
R84401 VDD.n1383 VDD.n1157 4.5005
R84402 VDD.n1306 VDD.n1157 4.5005
R84403 VDD.n1384 VDD.n1157 4.5005
R84404 VDD.n1304 VDD.n1157 4.5005
R84405 VDD.n1385 VDD.n1157 4.5005
R84406 VDD.n1303 VDD.n1157 4.5005
R84407 VDD.n1386 VDD.n1157 4.5005
R84408 VDD.n1301 VDD.n1157 4.5005
R84409 VDD.n1387 VDD.n1157 4.5005
R84410 VDD.n1300 VDD.n1157 4.5005
R84411 VDD.n1388 VDD.n1157 4.5005
R84412 VDD.n1298 VDD.n1157 4.5005
R84413 VDD.n1389 VDD.n1157 4.5005
R84414 VDD.n1297 VDD.n1157 4.5005
R84415 VDD.n1390 VDD.n1157 4.5005
R84416 VDD.n1295 VDD.n1157 4.5005
R84417 VDD.n1391 VDD.n1157 4.5005
R84418 VDD.n1294 VDD.n1157 4.5005
R84419 VDD.n1392 VDD.n1157 4.5005
R84420 VDD.n1292 VDD.n1157 4.5005
R84421 VDD.n1393 VDD.n1157 4.5005
R84422 VDD.n1291 VDD.n1157 4.5005
R84423 VDD.n1394 VDD.n1157 4.5005
R84424 VDD.n1289 VDD.n1157 4.5005
R84425 VDD.n1395 VDD.n1157 4.5005
R84426 VDD.n1288 VDD.n1157 4.5005
R84427 VDD.n1396 VDD.n1157 4.5005
R84428 VDD.n1286 VDD.n1157 4.5005
R84429 VDD.n1397 VDD.n1157 4.5005
R84430 VDD.n1285 VDD.n1157 4.5005
R84431 VDD.n1398 VDD.n1157 4.5005
R84432 VDD.n1283 VDD.n1157 4.5005
R84433 VDD.n1399 VDD.n1157 4.5005
R84434 VDD.n1282 VDD.n1157 4.5005
R84435 VDD.n1400 VDD.n1157 4.5005
R84436 VDD.n1280 VDD.n1157 4.5005
R84437 VDD.n1401 VDD.n1157 4.5005
R84438 VDD.n1279 VDD.n1157 4.5005
R84439 VDD.n1402 VDD.n1157 4.5005
R84440 VDD.n1277 VDD.n1157 4.5005
R84441 VDD.n1403 VDD.n1157 4.5005
R84442 VDD.n1276 VDD.n1157 4.5005
R84443 VDD.n1404 VDD.n1157 4.5005
R84444 VDD.n1274 VDD.n1157 4.5005
R84445 VDD.n1405 VDD.n1157 4.5005
R84446 VDD.n1273 VDD.n1157 4.5005
R84447 VDD.n1406 VDD.n1157 4.5005
R84448 VDD.n1271 VDD.n1157 4.5005
R84449 VDD.n1407 VDD.n1157 4.5005
R84450 VDD.n1270 VDD.n1157 4.5005
R84451 VDD.n1408 VDD.n1157 4.5005
R84452 VDD.n1268 VDD.n1157 4.5005
R84453 VDD.n1409 VDD.n1157 4.5005
R84454 VDD.n1267 VDD.n1157 4.5005
R84455 VDD.n1410 VDD.n1157 4.5005
R84456 VDD.n1265 VDD.n1157 4.5005
R84457 VDD.n1411 VDD.n1157 4.5005
R84458 VDD.n1264 VDD.n1157 4.5005
R84459 VDD.n1412 VDD.n1157 4.5005
R84460 VDD.n1262 VDD.n1157 4.5005
R84461 VDD.n1413 VDD.n1157 4.5005
R84462 VDD.n1261 VDD.n1157 4.5005
R84463 VDD.n1414 VDD.n1157 4.5005
R84464 VDD.n1415 VDD.n1157 4.5005
R84465 VDD.n1674 VDD.n1157 4.5005
R84466 VDD.n1676 VDD.n1233 4.5005
R84467 VDD.n1341 VDD.n1233 4.5005
R84468 VDD.n1342 VDD.n1233 4.5005
R84469 VDD.n1340 VDD.n1233 4.5005
R84470 VDD.n1344 VDD.n1233 4.5005
R84471 VDD.n1339 VDD.n1233 4.5005
R84472 VDD.n1345 VDD.n1233 4.5005
R84473 VDD.n1338 VDD.n1233 4.5005
R84474 VDD.n1347 VDD.n1233 4.5005
R84475 VDD.n1337 VDD.n1233 4.5005
R84476 VDD.n1348 VDD.n1233 4.5005
R84477 VDD.n1336 VDD.n1233 4.5005
R84478 VDD.n1350 VDD.n1233 4.5005
R84479 VDD.n1335 VDD.n1233 4.5005
R84480 VDD.n1351 VDD.n1233 4.5005
R84481 VDD.n1334 VDD.n1233 4.5005
R84482 VDD.n1353 VDD.n1233 4.5005
R84483 VDD.n1333 VDD.n1233 4.5005
R84484 VDD.n1354 VDD.n1233 4.5005
R84485 VDD.n1332 VDD.n1233 4.5005
R84486 VDD.n1356 VDD.n1233 4.5005
R84487 VDD.n1331 VDD.n1233 4.5005
R84488 VDD.n1357 VDD.n1233 4.5005
R84489 VDD.n1330 VDD.n1233 4.5005
R84490 VDD.n1359 VDD.n1233 4.5005
R84491 VDD.n1329 VDD.n1233 4.5005
R84492 VDD.n1360 VDD.n1233 4.5005
R84493 VDD.n1328 VDD.n1233 4.5005
R84494 VDD.n1362 VDD.n1233 4.5005
R84495 VDD.n1327 VDD.n1233 4.5005
R84496 VDD.n1363 VDD.n1233 4.5005
R84497 VDD.n1326 VDD.n1233 4.5005
R84498 VDD.n1365 VDD.n1233 4.5005
R84499 VDD.n1325 VDD.n1233 4.5005
R84500 VDD.n1366 VDD.n1233 4.5005
R84501 VDD.n1324 VDD.n1233 4.5005
R84502 VDD.n1368 VDD.n1233 4.5005
R84503 VDD.n1323 VDD.n1233 4.5005
R84504 VDD.n1369 VDD.n1233 4.5005
R84505 VDD.n1322 VDD.n1233 4.5005
R84506 VDD.n1371 VDD.n1233 4.5005
R84507 VDD.n1321 VDD.n1233 4.5005
R84508 VDD.n1372 VDD.n1233 4.5005
R84509 VDD.n1320 VDD.n1233 4.5005
R84510 VDD.n1374 VDD.n1233 4.5005
R84511 VDD.n1319 VDD.n1233 4.5005
R84512 VDD.n1375 VDD.n1233 4.5005
R84513 VDD.n1318 VDD.n1233 4.5005
R84514 VDD.n1376 VDD.n1233 4.5005
R84515 VDD.n1316 VDD.n1233 4.5005
R84516 VDD.n1377 VDD.n1233 4.5005
R84517 VDD.n1315 VDD.n1233 4.5005
R84518 VDD.n1378 VDD.n1233 4.5005
R84519 VDD.n1313 VDD.n1233 4.5005
R84520 VDD.n1379 VDD.n1233 4.5005
R84521 VDD.n1312 VDD.n1233 4.5005
R84522 VDD.n1380 VDD.n1233 4.5005
R84523 VDD.n1310 VDD.n1233 4.5005
R84524 VDD.n1381 VDD.n1233 4.5005
R84525 VDD.n1309 VDD.n1233 4.5005
R84526 VDD.n1382 VDD.n1233 4.5005
R84527 VDD.n1307 VDD.n1233 4.5005
R84528 VDD.n1383 VDD.n1233 4.5005
R84529 VDD.n1306 VDD.n1233 4.5005
R84530 VDD.n1384 VDD.n1233 4.5005
R84531 VDD.n1304 VDD.n1233 4.5005
R84532 VDD.n1385 VDD.n1233 4.5005
R84533 VDD.n1303 VDD.n1233 4.5005
R84534 VDD.n1386 VDD.n1233 4.5005
R84535 VDD.n1301 VDD.n1233 4.5005
R84536 VDD.n1387 VDD.n1233 4.5005
R84537 VDD.n1300 VDD.n1233 4.5005
R84538 VDD.n1388 VDD.n1233 4.5005
R84539 VDD.n1298 VDD.n1233 4.5005
R84540 VDD.n1389 VDD.n1233 4.5005
R84541 VDD.n1297 VDD.n1233 4.5005
R84542 VDD.n1390 VDD.n1233 4.5005
R84543 VDD.n1295 VDD.n1233 4.5005
R84544 VDD.n1391 VDD.n1233 4.5005
R84545 VDD.n1294 VDD.n1233 4.5005
R84546 VDD.n1392 VDD.n1233 4.5005
R84547 VDD.n1292 VDD.n1233 4.5005
R84548 VDD.n1393 VDD.n1233 4.5005
R84549 VDD.n1291 VDD.n1233 4.5005
R84550 VDD.n1394 VDD.n1233 4.5005
R84551 VDD.n1289 VDD.n1233 4.5005
R84552 VDD.n1395 VDD.n1233 4.5005
R84553 VDD.n1288 VDD.n1233 4.5005
R84554 VDD.n1396 VDD.n1233 4.5005
R84555 VDD.n1286 VDD.n1233 4.5005
R84556 VDD.n1397 VDD.n1233 4.5005
R84557 VDD.n1285 VDD.n1233 4.5005
R84558 VDD.n1398 VDD.n1233 4.5005
R84559 VDD.n1283 VDD.n1233 4.5005
R84560 VDD.n1399 VDD.n1233 4.5005
R84561 VDD.n1282 VDD.n1233 4.5005
R84562 VDD.n1400 VDD.n1233 4.5005
R84563 VDD.n1280 VDD.n1233 4.5005
R84564 VDD.n1401 VDD.n1233 4.5005
R84565 VDD.n1279 VDD.n1233 4.5005
R84566 VDD.n1402 VDD.n1233 4.5005
R84567 VDD.n1277 VDD.n1233 4.5005
R84568 VDD.n1403 VDD.n1233 4.5005
R84569 VDD.n1276 VDD.n1233 4.5005
R84570 VDD.n1404 VDD.n1233 4.5005
R84571 VDD.n1274 VDD.n1233 4.5005
R84572 VDD.n1405 VDD.n1233 4.5005
R84573 VDD.n1273 VDD.n1233 4.5005
R84574 VDD.n1406 VDD.n1233 4.5005
R84575 VDD.n1271 VDD.n1233 4.5005
R84576 VDD.n1407 VDD.n1233 4.5005
R84577 VDD.n1270 VDD.n1233 4.5005
R84578 VDD.n1408 VDD.n1233 4.5005
R84579 VDD.n1268 VDD.n1233 4.5005
R84580 VDD.n1409 VDD.n1233 4.5005
R84581 VDD.n1267 VDD.n1233 4.5005
R84582 VDD.n1410 VDD.n1233 4.5005
R84583 VDD.n1265 VDD.n1233 4.5005
R84584 VDD.n1411 VDD.n1233 4.5005
R84585 VDD.n1264 VDD.n1233 4.5005
R84586 VDD.n1412 VDD.n1233 4.5005
R84587 VDD.n1262 VDD.n1233 4.5005
R84588 VDD.n1413 VDD.n1233 4.5005
R84589 VDD.n1261 VDD.n1233 4.5005
R84590 VDD.n1414 VDD.n1233 4.5005
R84591 VDD.n1415 VDD.n1233 4.5005
R84592 VDD.n1674 VDD.n1233 4.5005
R84593 VDD.n1676 VDD.n1156 4.5005
R84594 VDD.n1341 VDD.n1156 4.5005
R84595 VDD.n1342 VDD.n1156 4.5005
R84596 VDD.n1340 VDD.n1156 4.5005
R84597 VDD.n1344 VDD.n1156 4.5005
R84598 VDD.n1339 VDD.n1156 4.5005
R84599 VDD.n1345 VDD.n1156 4.5005
R84600 VDD.n1338 VDD.n1156 4.5005
R84601 VDD.n1347 VDD.n1156 4.5005
R84602 VDD.n1337 VDD.n1156 4.5005
R84603 VDD.n1348 VDD.n1156 4.5005
R84604 VDD.n1336 VDD.n1156 4.5005
R84605 VDD.n1350 VDD.n1156 4.5005
R84606 VDD.n1335 VDD.n1156 4.5005
R84607 VDD.n1351 VDD.n1156 4.5005
R84608 VDD.n1334 VDD.n1156 4.5005
R84609 VDD.n1353 VDD.n1156 4.5005
R84610 VDD.n1333 VDD.n1156 4.5005
R84611 VDD.n1354 VDD.n1156 4.5005
R84612 VDD.n1332 VDD.n1156 4.5005
R84613 VDD.n1356 VDD.n1156 4.5005
R84614 VDD.n1331 VDD.n1156 4.5005
R84615 VDD.n1357 VDD.n1156 4.5005
R84616 VDD.n1330 VDD.n1156 4.5005
R84617 VDD.n1359 VDD.n1156 4.5005
R84618 VDD.n1329 VDD.n1156 4.5005
R84619 VDD.n1360 VDD.n1156 4.5005
R84620 VDD.n1328 VDD.n1156 4.5005
R84621 VDD.n1362 VDD.n1156 4.5005
R84622 VDD.n1327 VDD.n1156 4.5005
R84623 VDD.n1363 VDD.n1156 4.5005
R84624 VDD.n1326 VDD.n1156 4.5005
R84625 VDD.n1365 VDD.n1156 4.5005
R84626 VDD.n1325 VDD.n1156 4.5005
R84627 VDD.n1366 VDD.n1156 4.5005
R84628 VDD.n1324 VDD.n1156 4.5005
R84629 VDD.n1368 VDD.n1156 4.5005
R84630 VDD.n1323 VDD.n1156 4.5005
R84631 VDD.n1369 VDD.n1156 4.5005
R84632 VDD.n1322 VDD.n1156 4.5005
R84633 VDD.n1371 VDD.n1156 4.5005
R84634 VDD.n1321 VDD.n1156 4.5005
R84635 VDD.n1372 VDD.n1156 4.5005
R84636 VDD.n1320 VDD.n1156 4.5005
R84637 VDD.n1374 VDD.n1156 4.5005
R84638 VDD.n1319 VDD.n1156 4.5005
R84639 VDD.n1375 VDD.n1156 4.5005
R84640 VDD.n1318 VDD.n1156 4.5005
R84641 VDD.n1376 VDD.n1156 4.5005
R84642 VDD.n1316 VDD.n1156 4.5005
R84643 VDD.n1377 VDD.n1156 4.5005
R84644 VDD.n1315 VDD.n1156 4.5005
R84645 VDD.n1378 VDD.n1156 4.5005
R84646 VDD.n1313 VDD.n1156 4.5005
R84647 VDD.n1379 VDD.n1156 4.5005
R84648 VDD.n1312 VDD.n1156 4.5005
R84649 VDD.n1380 VDD.n1156 4.5005
R84650 VDD.n1310 VDD.n1156 4.5005
R84651 VDD.n1381 VDD.n1156 4.5005
R84652 VDD.n1309 VDD.n1156 4.5005
R84653 VDD.n1382 VDD.n1156 4.5005
R84654 VDD.n1307 VDD.n1156 4.5005
R84655 VDD.n1383 VDD.n1156 4.5005
R84656 VDD.n1306 VDD.n1156 4.5005
R84657 VDD.n1384 VDD.n1156 4.5005
R84658 VDD.n1304 VDD.n1156 4.5005
R84659 VDD.n1385 VDD.n1156 4.5005
R84660 VDD.n1303 VDD.n1156 4.5005
R84661 VDD.n1386 VDD.n1156 4.5005
R84662 VDD.n1301 VDD.n1156 4.5005
R84663 VDD.n1387 VDD.n1156 4.5005
R84664 VDD.n1300 VDD.n1156 4.5005
R84665 VDD.n1388 VDD.n1156 4.5005
R84666 VDD.n1298 VDD.n1156 4.5005
R84667 VDD.n1389 VDD.n1156 4.5005
R84668 VDD.n1297 VDD.n1156 4.5005
R84669 VDD.n1390 VDD.n1156 4.5005
R84670 VDD.n1295 VDD.n1156 4.5005
R84671 VDD.n1391 VDD.n1156 4.5005
R84672 VDD.n1294 VDD.n1156 4.5005
R84673 VDD.n1392 VDD.n1156 4.5005
R84674 VDD.n1292 VDD.n1156 4.5005
R84675 VDD.n1393 VDD.n1156 4.5005
R84676 VDD.n1291 VDD.n1156 4.5005
R84677 VDD.n1394 VDD.n1156 4.5005
R84678 VDD.n1289 VDD.n1156 4.5005
R84679 VDD.n1395 VDD.n1156 4.5005
R84680 VDD.n1288 VDD.n1156 4.5005
R84681 VDD.n1396 VDD.n1156 4.5005
R84682 VDD.n1286 VDD.n1156 4.5005
R84683 VDD.n1397 VDD.n1156 4.5005
R84684 VDD.n1285 VDD.n1156 4.5005
R84685 VDD.n1398 VDD.n1156 4.5005
R84686 VDD.n1283 VDD.n1156 4.5005
R84687 VDD.n1399 VDD.n1156 4.5005
R84688 VDD.n1282 VDD.n1156 4.5005
R84689 VDD.n1400 VDD.n1156 4.5005
R84690 VDD.n1280 VDD.n1156 4.5005
R84691 VDD.n1401 VDD.n1156 4.5005
R84692 VDD.n1279 VDD.n1156 4.5005
R84693 VDD.n1402 VDD.n1156 4.5005
R84694 VDD.n1277 VDD.n1156 4.5005
R84695 VDD.n1403 VDD.n1156 4.5005
R84696 VDD.n1276 VDD.n1156 4.5005
R84697 VDD.n1404 VDD.n1156 4.5005
R84698 VDD.n1274 VDD.n1156 4.5005
R84699 VDD.n1405 VDD.n1156 4.5005
R84700 VDD.n1273 VDD.n1156 4.5005
R84701 VDD.n1406 VDD.n1156 4.5005
R84702 VDD.n1271 VDD.n1156 4.5005
R84703 VDD.n1407 VDD.n1156 4.5005
R84704 VDD.n1270 VDD.n1156 4.5005
R84705 VDD.n1408 VDD.n1156 4.5005
R84706 VDD.n1268 VDD.n1156 4.5005
R84707 VDD.n1409 VDD.n1156 4.5005
R84708 VDD.n1267 VDD.n1156 4.5005
R84709 VDD.n1410 VDD.n1156 4.5005
R84710 VDD.n1265 VDD.n1156 4.5005
R84711 VDD.n1411 VDD.n1156 4.5005
R84712 VDD.n1264 VDD.n1156 4.5005
R84713 VDD.n1412 VDD.n1156 4.5005
R84714 VDD.n1262 VDD.n1156 4.5005
R84715 VDD.n1413 VDD.n1156 4.5005
R84716 VDD.n1261 VDD.n1156 4.5005
R84717 VDD.n1414 VDD.n1156 4.5005
R84718 VDD.n1415 VDD.n1156 4.5005
R84719 VDD.n1674 VDD.n1156 4.5005
R84720 VDD.n1676 VDD.n1234 4.5005
R84721 VDD.n1341 VDD.n1234 4.5005
R84722 VDD.n1342 VDD.n1234 4.5005
R84723 VDD.n1340 VDD.n1234 4.5005
R84724 VDD.n1344 VDD.n1234 4.5005
R84725 VDD.n1339 VDD.n1234 4.5005
R84726 VDD.n1345 VDD.n1234 4.5005
R84727 VDD.n1338 VDD.n1234 4.5005
R84728 VDD.n1347 VDD.n1234 4.5005
R84729 VDD.n1337 VDD.n1234 4.5005
R84730 VDD.n1348 VDD.n1234 4.5005
R84731 VDD.n1336 VDD.n1234 4.5005
R84732 VDD.n1350 VDD.n1234 4.5005
R84733 VDD.n1335 VDD.n1234 4.5005
R84734 VDD.n1351 VDD.n1234 4.5005
R84735 VDD.n1334 VDD.n1234 4.5005
R84736 VDD.n1353 VDD.n1234 4.5005
R84737 VDD.n1333 VDD.n1234 4.5005
R84738 VDD.n1354 VDD.n1234 4.5005
R84739 VDD.n1332 VDD.n1234 4.5005
R84740 VDD.n1356 VDD.n1234 4.5005
R84741 VDD.n1331 VDD.n1234 4.5005
R84742 VDD.n1357 VDD.n1234 4.5005
R84743 VDD.n1330 VDD.n1234 4.5005
R84744 VDD.n1359 VDD.n1234 4.5005
R84745 VDD.n1329 VDD.n1234 4.5005
R84746 VDD.n1360 VDD.n1234 4.5005
R84747 VDD.n1328 VDD.n1234 4.5005
R84748 VDD.n1362 VDD.n1234 4.5005
R84749 VDD.n1327 VDD.n1234 4.5005
R84750 VDD.n1363 VDD.n1234 4.5005
R84751 VDD.n1326 VDD.n1234 4.5005
R84752 VDD.n1365 VDD.n1234 4.5005
R84753 VDD.n1325 VDD.n1234 4.5005
R84754 VDD.n1366 VDD.n1234 4.5005
R84755 VDD.n1324 VDD.n1234 4.5005
R84756 VDD.n1368 VDD.n1234 4.5005
R84757 VDD.n1323 VDD.n1234 4.5005
R84758 VDD.n1369 VDD.n1234 4.5005
R84759 VDD.n1322 VDD.n1234 4.5005
R84760 VDD.n1371 VDD.n1234 4.5005
R84761 VDD.n1321 VDD.n1234 4.5005
R84762 VDD.n1372 VDD.n1234 4.5005
R84763 VDD.n1320 VDD.n1234 4.5005
R84764 VDD.n1374 VDD.n1234 4.5005
R84765 VDD.n1319 VDD.n1234 4.5005
R84766 VDD.n1375 VDD.n1234 4.5005
R84767 VDD.n1318 VDD.n1234 4.5005
R84768 VDD.n1376 VDD.n1234 4.5005
R84769 VDD.n1316 VDD.n1234 4.5005
R84770 VDD.n1377 VDD.n1234 4.5005
R84771 VDD.n1315 VDD.n1234 4.5005
R84772 VDD.n1378 VDD.n1234 4.5005
R84773 VDD.n1313 VDD.n1234 4.5005
R84774 VDD.n1379 VDD.n1234 4.5005
R84775 VDD.n1312 VDD.n1234 4.5005
R84776 VDD.n1380 VDD.n1234 4.5005
R84777 VDD.n1310 VDD.n1234 4.5005
R84778 VDD.n1381 VDD.n1234 4.5005
R84779 VDD.n1309 VDD.n1234 4.5005
R84780 VDD.n1382 VDD.n1234 4.5005
R84781 VDD.n1307 VDD.n1234 4.5005
R84782 VDD.n1383 VDD.n1234 4.5005
R84783 VDD.n1306 VDD.n1234 4.5005
R84784 VDD.n1384 VDD.n1234 4.5005
R84785 VDD.n1304 VDD.n1234 4.5005
R84786 VDD.n1385 VDD.n1234 4.5005
R84787 VDD.n1303 VDD.n1234 4.5005
R84788 VDD.n1386 VDD.n1234 4.5005
R84789 VDD.n1301 VDD.n1234 4.5005
R84790 VDD.n1387 VDD.n1234 4.5005
R84791 VDD.n1300 VDD.n1234 4.5005
R84792 VDD.n1388 VDD.n1234 4.5005
R84793 VDD.n1298 VDD.n1234 4.5005
R84794 VDD.n1389 VDD.n1234 4.5005
R84795 VDD.n1297 VDD.n1234 4.5005
R84796 VDD.n1390 VDD.n1234 4.5005
R84797 VDD.n1295 VDD.n1234 4.5005
R84798 VDD.n1391 VDD.n1234 4.5005
R84799 VDD.n1294 VDD.n1234 4.5005
R84800 VDD.n1392 VDD.n1234 4.5005
R84801 VDD.n1292 VDD.n1234 4.5005
R84802 VDD.n1393 VDD.n1234 4.5005
R84803 VDD.n1291 VDD.n1234 4.5005
R84804 VDD.n1394 VDD.n1234 4.5005
R84805 VDD.n1289 VDD.n1234 4.5005
R84806 VDD.n1395 VDD.n1234 4.5005
R84807 VDD.n1288 VDD.n1234 4.5005
R84808 VDD.n1396 VDD.n1234 4.5005
R84809 VDD.n1286 VDD.n1234 4.5005
R84810 VDD.n1397 VDD.n1234 4.5005
R84811 VDD.n1285 VDD.n1234 4.5005
R84812 VDD.n1398 VDD.n1234 4.5005
R84813 VDD.n1283 VDD.n1234 4.5005
R84814 VDD.n1399 VDD.n1234 4.5005
R84815 VDD.n1282 VDD.n1234 4.5005
R84816 VDD.n1400 VDD.n1234 4.5005
R84817 VDD.n1280 VDD.n1234 4.5005
R84818 VDD.n1401 VDD.n1234 4.5005
R84819 VDD.n1279 VDD.n1234 4.5005
R84820 VDD.n1402 VDD.n1234 4.5005
R84821 VDD.n1277 VDD.n1234 4.5005
R84822 VDD.n1403 VDD.n1234 4.5005
R84823 VDD.n1276 VDD.n1234 4.5005
R84824 VDD.n1404 VDD.n1234 4.5005
R84825 VDD.n1274 VDD.n1234 4.5005
R84826 VDD.n1405 VDD.n1234 4.5005
R84827 VDD.n1273 VDD.n1234 4.5005
R84828 VDD.n1406 VDD.n1234 4.5005
R84829 VDD.n1271 VDD.n1234 4.5005
R84830 VDD.n1407 VDD.n1234 4.5005
R84831 VDD.n1270 VDD.n1234 4.5005
R84832 VDD.n1408 VDD.n1234 4.5005
R84833 VDD.n1268 VDD.n1234 4.5005
R84834 VDD.n1409 VDD.n1234 4.5005
R84835 VDD.n1267 VDD.n1234 4.5005
R84836 VDD.n1410 VDD.n1234 4.5005
R84837 VDD.n1265 VDD.n1234 4.5005
R84838 VDD.n1411 VDD.n1234 4.5005
R84839 VDD.n1264 VDD.n1234 4.5005
R84840 VDD.n1412 VDD.n1234 4.5005
R84841 VDD.n1262 VDD.n1234 4.5005
R84842 VDD.n1413 VDD.n1234 4.5005
R84843 VDD.n1261 VDD.n1234 4.5005
R84844 VDD.n1414 VDD.n1234 4.5005
R84845 VDD.n1415 VDD.n1234 4.5005
R84846 VDD.n1674 VDD.n1234 4.5005
R84847 VDD.n1676 VDD.n1155 4.5005
R84848 VDD.n1341 VDD.n1155 4.5005
R84849 VDD.n1342 VDD.n1155 4.5005
R84850 VDD.n1340 VDD.n1155 4.5005
R84851 VDD.n1344 VDD.n1155 4.5005
R84852 VDD.n1339 VDD.n1155 4.5005
R84853 VDD.n1345 VDD.n1155 4.5005
R84854 VDD.n1338 VDD.n1155 4.5005
R84855 VDD.n1347 VDD.n1155 4.5005
R84856 VDD.n1337 VDD.n1155 4.5005
R84857 VDD.n1348 VDD.n1155 4.5005
R84858 VDD.n1336 VDD.n1155 4.5005
R84859 VDD.n1350 VDD.n1155 4.5005
R84860 VDD.n1335 VDD.n1155 4.5005
R84861 VDD.n1351 VDD.n1155 4.5005
R84862 VDD.n1334 VDD.n1155 4.5005
R84863 VDD.n1353 VDD.n1155 4.5005
R84864 VDD.n1333 VDD.n1155 4.5005
R84865 VDD.n1354 VDD.n1155 4.5005
R84866 VDD.n1332 VDD.n1155 4.5005
R84867 VDD.n1356 VDD.n1155 4.5005
R84868 VDD.n1331 VDD.n1155 4.5005
R84869 VDD.n1357 VDD.n1155 4.5005
R84870 VDD.n1330 VDD.n1155 4.5005
R84871 VDD.n1359 VDD.n1155 4.5005
R84872 VDD.n1329 VDD.n1155 4.5005
R84873 VDD.n1360 VDD.n1155 4.5005
R84874 VDD.n1328 VDD.n1155 4.5005
R84875 VDD.n1362 VDD.n1155 4.5005
R84876 VDD.n1327 VDD.n1155 4.5005
R84877 VDD.n1363 VDD.n1155 4.5005
R84878 VDD.n1326 VDD.n1155 4.5005
R84879 VDD.n1365 VDD.n1155 4.5005
R84880 VDD.n1325 VDD.n1155 4.5005
R84881 VDD.n1366 VDD.n1155 4.5005
R84882 VDD.n1324 VDD.n1155 4.5005
R84883 VDD.n1368 VDD.n1155 4.5005
R84884 VDD.n1323 VDD.n1155 4.5005
R84885 VDD.n1369 VDD.n1155 4.5005
R84886 VDD.n1322 VDD.n1155 4.5005
R84887 VDD.n1371 VDD.n1155 4.5005
R84888 VDD.n1321 VDD.n1155 4.5005
R84889 VDD.n1372 VDD.n1155 4.5005
R84890 VDD.n1320 VDD.n1155 4.5005
R84891 VDD.n1374 VDD.n1155 4.5005
R84892 VDD.n1319 VDD.n1155 4.5005
R84893 VDD.n1375 VDD.n1155 4.5005
R84894 VDD.n1318 VDD.n1155 4.5005
R84895 VDD.n1376 VDD.n1155 4.5005
R84896 VDD.n1316 VDD.n1155 4.5005
R84897 VDD.n1377 VDD.n1155 4.5005
R84898 VDD.n1315 VDD.n1155 4.5005
R84899 VDD.n1378 VDD.n1155 4.5005
R84900 VDD.n1313 VDD.n1155 4.5005
R84901 VDD.n1379 VDD.n1155 4.5005
R84902 VDD.n1312 VDD.n1155 4.5005
R84903 VDD.n1380 VDD.n1155 4.5005
R84904 VDD.n1310 VDD.n1155 4.5005
R84905 VDD.n1381 VDD.n1155 4.5005
R84906 VDD.n1309 VDD.n1155 4.5005
R84907 VDD.n1382 VDD.n1155 4.5005
R84908 VDD.n1307 VDD.n1155 4.5005
R84909 VDD.n1383 VDD.n1155 4.5005
R84910 VDD.n1306 VDD.n1155 4.5005
R84911 VDD.n1384 VDD.n1155 4.5005
R84912 VDD.n1304 VDD.n1155 4.5005
R84913 VDD.n1385 VDD.n1155 4.5005
R84914 VDD.n1303 VDD.n1155 4.5005
R84915 VDD.n1386 VDD.n1155 4.5005
R84916 VDD.n1301 VDD.n1155 4.5005
R84917 VDD.n1387 VDD.n1155 4.5005
R84918 VDD.n1300 VDD.n1155 4.5005
R84919 VDD.n1388 VDD.n1155 4.5005
R84920 VDD.n1298 VDD.n1155 4.5005
R84921 VDD.n1389 VDD.n1155 4.5005
R84922 VDD.n1297 VDD.n1155 4.5005
R84923 VDD.n1390 VDD.n1155 4.5005
R84924 VDD.n1295 VDD.n1155 4.5005
R84925 VDD.n1391 VDD.n1155 4.5005
R84926 VDD.n1294 VDD.n1155 4.5005
R84927 VDD.n1392 VDD.n1155 4.5005
R84928 VDD.n1292 VDD.n1155 4.5005
R84929 VDD.n1393 VDD.n1155 4.5005
R84930 VDD.n1291 VDD.n1155 4.5005
R84931 VDD.n1394 VDD.n1155 4.5005
R84932 VDD.n1289 VDD.n1155 4.5005
R84933 VDD.n1395 VDD.n1155 4.5005
R84934 VDD.n1288 VDD.n1155 4.5005
R84935 VDD.n1396 VDD.n1155 4.5005
R84936 VDD.n1286 VDD.n1155 4.5005
R84937 VDD.n1397 VDD.n1155 4.5005
R84938 VDD.n1285 VDD.n1155 4.5005
R84939 VDD.n1398 VDD.n1155 4.5005
R84940 VDD.n1283 VDD.n1155 4.5005
R84941 VDD.n1399 VDD.n1155 4.5005
R84942 VDD.n1282 VDD.n1155 4.5005
R84943 VDD.n1400 VDD.n1155 4.5005
R84944 VDD.n1280 VDD.n1155 4.5005
R84945 VDD.n1401 VDD.n1155 4.5005
R84946 VDD.n1279 VDD.n1155 4.5005
R84947 VDD.n1402 VDD.n1155 4.5005
R84948 VDD.n1277 VDD.n1155 4.5005
R84949 VDD.n1403 VDD.n1155 4.5005
R84950 VDD.n1276 VDD.n1155 4.5005
R84951 VDD.n1404 VDD.n1155 4.5005
R84952 VDD.n1274 VDD.n1155 4.5005
R84953 VDD.n1405 VDD.n1155 4.5005
R84954 VDD.n1273 VDD.n1155 4.5005
R84955 VDD.n1406 VDD.n1155 4.5005
R84956 VDD.n1271 VDD.n1155 4.5005
R84957 VDD.n1407 VDD.n1155 4.5005
R84958 VDD.n1270 VDD.n1155 4.5005
R84959 VDD.n1408 VDD.n1155 4.5005
R84960 VDD.n1268 VDD.n1155 4.5005
R84961 VDD.n1409 VDD.n1155 4.5005
R84962 VDD.n1267 VDD.n1155 4.5005
R84963 VDD.n1410 VDD.n1155 4.5005
R84964 VDD.n1265 VDD.n1155 4.5005
R84965 VDD.n1411 VDD.n1155 4.5005
R84966 VDD.n1264 VDD.n1155 4.5005
R84967 VDD.n1412 VDD.n1155 4.5005
R84968 VDD.n1262 VDD.n1155 4.5005
R84969 VDD.n1413 VDD.n1155 4.5005
R84970 VDD.n1261 VDD.n1155 4.5005
R84971 VDD.n1414 VDD.n1155 4.5005
R84972 VDD.n1415 VDD.n1155 4.5005
R84973 VDD.n1674 VDD.n1155 4.5005
R84974 VDD.n1676 VDD.n1235 4.5005
R84975 VDD.n1341 VDD.n1235 4.5005
R84976 VDD.n1342 VDD.n1235 4.5005
R84977 VDD.n1340 VDD.n1235 4.5005
R84978 VDD.n1344 VDD.n1235 4.5005
R84979 VDD.n1339 VDD.n1235 4.5005
R84980 VDD.n1345 VDD.n1235 4.5005
R84981 VDD.n1338 VDD.n1235 4.5005
R84982 VDD.n1347 VDD.n1235 4.5005
R84983 VDD.n1337 VDD.n1235 4.5005
R84984 VDD.n1348 VDD.n1235 4.5005
R84985 VDD.n1336 VDD.n1235 4.5005
R84986 VDD.n1350 VDD.n1235 4.5005
R84987 VDD.n1335 VDD.n1235 4.5005
R84988 VDD.n1351 VDD.n1235 4.5005
R84989 VDD.n1334 VDD.n1235 4.5005
R84990 VDD.n1353 VDD.n1235 4.5005
R84991 VDD.n1333 VDD.n1235 4.5005
R84992 VDD.n1354 VDD.n1235 4.5005
R84993 VDD.n1332 VDD.n1235 4.5005
R84994 VDD.n1356 VDD.n1235 4.5005
R84995 VDD.n1331 VDD.n1235 4.5005
R84996 VDD.n1357 VDD.n1235 4.5005
R84997 VDD.n1330 VDD.n1235 4.5005
R84998 VDD.n1359 VDD.n1235 4.5005
R84999 VDD.n1329 VDD.n1235 4.5005
R85000 VDD.n1360 VDD.n1235 4.5005
R85001 VDD.n1328 VDD.n1235 4.5005
R85002 VDD.n1362 VDD.n1235 4.5005
R85003 VDD.n1327 VDD.n1235 4.5005
R85004 VDD.n1363 VDD.n1235 4.5005
R85005 VDD.n1326 VDD.n1235 4.5005
R85006 VDD.n1365 VDD.n1235 4.5005
R85007 VDD.n1325 VDD.n1235 4.5005
R85008 VDD.n1366 VDD.n1235 4.5005
R85009 VDD.n1324 VDD.n1235 4.5005
R85010 VDD.n1368 VDD.n1235 4.5005
R85011 VDD.n1323 VDD.n1235 4.5005
R85012 VDD.n1369 VDD.n1235 4.5005
R85013 VDD.n1322 VDD.n1235 4.5005
R85014 VDD.n1371 VDD.n1235 4.5005
R85015 VDD.n1321 VDD.n1235 4.5005
R85016 VDD.n1372 VDD.n1235 4.5005
R85017 VDD.n1320 VDD.n1235 4.5005
R85018 VDD.n1374 VDD.n1235 4.5005
R85019 VDD.n1319 VDD.n1235 4.5005
R85020 VDD.n1375 VDD.n1235 4.5005
R85021 VDD.n1318 VDD.n1235 4.5005
R85022 VDD.n1376 VDD.n1235 4.5005
R85023 VDD.n1316 VDD.n1235 4.5005
R85024 VDD.n1377 VDD.n1235 4.5005
R85025 VDD.n1315 VDD.n1235 4.5005
R85026 VDD.n1378 VDD.n1235 4.5005
R85027 VDD.n1313 VDD.n1235 4.5005
R85028 VDD.n1379 VDD.n1235 4.5005
R85029 VDD.n1312 VDD.n1235 4.5005
R85030 VDD.n1380 VDD.n1235 4.5005
R85031 VDD.n1310 VDD.n1235 4.5005
R85032 VDD.n1381 VDD.n1235 4.5005
R85033 VDD.n1309 VDD.n1235 4.5005
R85034 VDD.n1382 VDD.n1235 4.5005
R85035 VDD.n1307 VDD.n1235 4.5005
R85036 VDD.n1383 VDD.n1235 4.5005
R85037 VDD.n1306 VDD.n1235 4.5005
R85038 VDD.n1384 VDD.n1235 4.5005
R85039 VDD.n1304 VDD.n1235 4.5005
R85040 VDD.n1385 VDD.n1235 4.5005
R85041 VDD.n1303 VDD.n1235 4.5005
R85042 VDD.n1386 VDD.n1235 4.5005
R85043 VDD.n1301 VDD.n1235 4.5005
R85044 VDD.n1387 VDD.n1235 4.5005
R85045 VDD.n1300 VDD.n1235 4.5005
R85046 VDD.n1388 VDD.n1235 4.5005
R85047 VDD.n1298 VDD.n1235 4.5005
R85048 VDD.n1389 VDD.n1235 4.5005
R85049 VDD.n1297 VDD.n1235 4.5005
R85050 VDD.n1390 VDD.n1235 4.5005
R85051 VDD.n1295 VDD.n1235 4.5005
R85052 VDD.n1391 VDD.n1235 4.5005
R85053 VDD.n1294 VDD.n1235 4.5005
R85054 VDD.n1392 VDD.n1235 4.5005
R85055 VDD.n1292 VDD.n1235 4.5005
R85056 VDD.n1393 VDD.n1235 4.5005
R85057 VDD.n1291 VDD.n1235 4.5005
R85058 VDD.n1394 VDD.n1235 4.5005
R85059 VDD.n1289 VDD.n1235 4.5005
R85060 VDD.n1395 VDD.n1235 4.5005
R85061 VDD.n1288 VDD.n1235 4.5005
R85062 VDD.n1396 VDD.n1235 4.5005
R85063 VDD.n1286 VDD.n1235 4.5005
R85064 VDD.n1397 VDD.n1235 4.5005
R85065 VDD.n1285 VDD.n1235 4.5005
R85066 VDD.n1398 VDD.n1235 4.5005
R85067 VDD.n1283 VDD.n1235 4.5005
R85068 VDD.n1399 VDD.n1235 4.5005
R85069 VDD.n1282 VDD.n1235 4.5005
R85070 VDD.n1400 VDD.n1235 4.5005
R85071 VDD.n1280 VDD.n1235 4.5005
R85072 VDD.n1401 VDD.n1235 4.5005
R85073 VDD.n1279 VDD.n1235 4.5005
R85074 VDD.n1402 VDD.n1235 4.5005
R85075 VDD.n1277 VDD.n1235 4.5005
R85076 VDD.n1403 VDD.n1235 4.5005
R85077 VDD.n1276 VDD.n1235 4.5005
R85078 VDD.n1404 VDD.n1235 4.5005
R85079 VDD.n1274 VDD.n1235 4.5005
R85080 VDD.n1405 VDD.n1235 4.5005
R85081 VDD.n1273 VDD.n1235 4.5005
R85082 VDD.n1406 VDD.n1235 4.5005
R85083 VDD.n1271 VDD.n1235 4.5005
R85084 VDD.n1407 VDD.n1235 4.5005
R85085 VDD.n1270 VDD.n1235 4.5005
R85086 VDD.n1408 VDD.n1235 4.5005
R85087 VDD.n1268 VDD.n1235 4.5005
R85088 VDD.n1409 VDD.n1235 4.5005
R85089 VDD.n1267 VDD.n1235 4.5005
R85090 VDD.n1410 VDD.n1235 4.5005
R85091 VDD.n1265 VDD.n1235 4.5005
R85092 VDD.n1411 VDD.n1235 4.5005
R85093 VDD.n1264 VDD.n1235 4.5005
R85094 VDD.n1412 VDD.n1235 4.5005
R85095 VDD.n1262 VDD.n1235 4.5005
R85096 VDD.n1413 VDD.n1235 4.5005
R85097 VDD.n1261 VDD.n1235 4.5005
R85098 VDD.n1414 VDD.n1235 4.5005
R85099 VDD.n1415 VDD.n1235 4.5005
R85100 VDD.n1674 VDD.n1235 4.5005
R85101 VDD.n1676 VDD.n1154 4.5005
R85102 VDD.n1341 VDD.n1154 4.5005
R85103 VDD.n1342 VDD.n1154 4.5005
R85104 VDD.n1340 VDD.n1154 4.5005
R85105 VDD.n1344 VDD.n1154 4.5005
R85106 VDD.n1339 VDD.n1154 4.5005
R85107 VDD.n1345 VDD.n1154 4.5005
R85108 VDD.n1338 VDD.n1154 4.5005
R85109 VDD.n1347 VDD.n1154 4.5005
R85110 VDD.n1337 VDD.n1154 4.5005
R85111 VDD.n1348 VDD.n1154 4.5005
R85112 VDD.n1336 VDD.n1154 4.5005
R85113 VDD.n1350 VDD.n1154 4.5005
R85114 VDD.n1335 VDD.n1154 4.5005
R85115 VDD.n1351 VDD.n1154 4.5005
R85116 VDD.n1334 VDD.n1154 4.5005
R85117 VDD.n1353 VDD.n1154 4.5005
R85118 VDD.n1333 VDD.n1154 4.5005
R85119 VDD.n1354 VDD.n1154 4.5005
R85120 VDD.n1332 VDD.n1154 4.5005
R85121 VDD.n1356 VDD.n1154 4.5005
R85122 VDD.n1331 VDD.n1154 4.5005
R85123 VDD.n1357 VDD.n1154 4.5005
R85124 VDD.n1330 VDD.n1154 4.5005
R85125 VDD.n1359 VDD.n1154 4.5005
R85126 VDD.n1329 VDD.n1154 4.5005
R85127 VDD.n1360 VDD.n1154 4.5005
R85128 VDD.n1328 VDD.n1154 4.5005
R85129 VDD.n1362 VDD.n1154 4.5005
R85130 VDD.n1327 VDD.n1154 4.5005
R85131 VDD.n1363 VDD.n1154 4.5005
R85132 VDD.n1326 VDD.n1154 4.5005
R85133 VDD.n1365 VDD.n1154 4.5005
R85134 VDD.n1325 VDD.n1154 4.5005
R85135 VDD.n1366 VDD.n1154 4.5005
R85136 VDD.n1324 VDD.n1154 4.5005
R85137 VDD.n1368 VDD.n1154 4.5005
R85138 VDD.n1323 VDD.n1154 4.5005
R85139 VDD.n1369 VDD.n1154 4.5005
R85140 VDD.n1322 VDD.n1154 4.5005
R85141 VDD.n1371 VDD.n1154 4.5005
R85142 VDD.n1321 VDD.n1154 4.5005
R85143 VDD.n1372 VDD.n1154 4.5005
R85144 VDD.n1320 VDD.n1154 4.5005
R85145 VDD.n1374 VDD.n1154 4.5005
R85146 VDD.n1319 VDD.n1154 4.5005
R85147 VDD.n1375 VDD.n1154 4.5005
R85148 VDD.n1318 VDD.n1154 4.5005
R85149 VDD.n1376 VDD.n1154 4.5005
R85150 VDD.n1316 VDD.n1154 4.5005
R85151 VDD.n1377 VDD.n1154 4.5005
R85152 VDD.n1315 VDD.n1154 4.5005
R85153 VDD.n1378 VDD.n1154 4.5005
R85154 VDD.n1313 VDD.n1154 4.5005
R85155 VDD.n1379 VDD.n1154 4.5005
R85156 VDD.n1312 VDD.n1154 4.5005
R85157 VDD.n1380 VDD.n1154 4.5005
R85158 VDD.n1310 VDD.n1154 4.5005
R85159 VDD.n1381 VDD.n1154 4.5005
R85160 VDD.n1309 VDD.n1154 4.5005
R85161 VDD.n1382 VDD.n1154 4.5005
R85162 VDD.n1307 VDD.n1154 4.5005
R85163 VDD.n1383 VDD.n1154 4.5005
R85164 VDD.n1306 VDD.n1154 4.5005
R85165 VDD.n1384 VDD.n1154 4.5005
R85166 VDD.n1304 VDD.n1154 4.5005
R85167 VDD.n1385 VDD.n1154 4.5005
R85168 VDD.n1303 VDD.n1154 4.5005
R85169 VDD.n1386 VDD.n1154 4.5005
R85170 VDD.n1301 VDD.n1154 4.5005
R85171 VDD.n1387 VDD.n1154 4.5005
R85172 VDD.n1300 VDD.n1154 4.5005
R85173 VDD.n1388 VDD.n1154 4.5005
R85174 VDD.n1298 VDD.n1154 4.5005
R85175 VDD.n1389 VDD.n1154 4.5005
R85176 VDD.n1297 VDD.n1154 4.5005
R85177 VDD.n1390 VDD.n1154 4.5005
R85178 VDD.n1295 VDD.n1154 4.5005
R85179 VDD.n1391 VDD.n1154 4.5005
R85180 VDD.n1294 VDD.n1154 4.5005
R85181 VDD.n1392 VDD.n1154 4.5005
R85182 VDD.n1292 VDD.n1154 4.5005
R85183 VDD.n1393 VDD.n1154 4.5005
R85184 VDD.n1291 VDD.n1154 4.5005
R85185 VDD.n1394 VDD.n1154 4.5005
R85186 VDD.n1289 VDD.n1154 4.5005
R85187 VDD.n1395 VDD.n1154 4.5005
R85188 VDD.n1288 VDD.n1154 4.5005
R85189 VDD.n1396 VDD.n1154 4.5005
R85190 VDD.n1286 VDD.n1154 4.5005
R85191 VDD.n1397 VDD.n1154 4.5005
R85192 VDD.n1285 VDD.n1154 4.5005
R85193 VDD.n1398 VDD.n1154 4.5005
R85194 VDD.n1283 VDD.n1154 4.5005
R85195 VDD.n1399 VDD.n1154 4.5005
R85196 VDD.n1282 VDD.n1154 4.5005
R85197 VDD.n1400 VDD.n1154 4.5005
R85198 VDD.n1280 VDD.n1154 4.5005
R85199 VDD.n1401 VDD.n1154 4.5005
R85200 VDD.n1279 VDD.n1154 4.5005
R85201 VDD.n1402 VDD.n1154 4.5005
R85202 VDD.n1277 VDD.n1154 4.5005
R85203 VDD.n1403 VDD.n1154 4.5005
R85204 VDD.n1276 VDD.n1154 4.5005
R85205 VDD.n1404 VDD.n1154 4.5005
R85206 VDD.n1274 VDD.n1154 4.5005
R85207 VDD.n1405 VDD.n1154 4.5005
R85208 VDD.n1273 VDD.n1154 4.5005
R85209 VDD.n1406 VDD.n1154 4.5005
R85210 VDD.n1271 VDD.n1154 4.5005
R85211 VDD.n1407 VDD.n1154 4.5005
R85212 VDD.n1270 VDD.n1154 4.5005
R85213 VDD.n1408 VDD.n1154 4.5005
R85214 VDD.n1268 VDD.n1154 4.5005
R85215 VDD.n1409 VDD.n1154 4.5005
R85216 VDD.n1267 VDD.n1154 4.5005
R85217 VDD.n1410 VDD.n1154 4.5005
R85218 VDD.n1265 VDD.n1154 4.5005
R85219 VDD.n1411 VDD.n1154 4.5005
R85220 VDD.n1264 VDD.n1154 4.5005
R85221 VDD.n1412 VDD.n1154 4.5005
R85222 VDD.n1262 VDD.n1154 4.5005
R85223 VDD.n1413 VDD.n1154 4.5005
R85224 VDD.n1261 VDD.n1154 4.5005
R85225 VDD.n1414 VDD.n1154 4.5005
R85226 VDD.n1415 VDD.n1154 4.5005
R85227 VDD.n1674 VDD.n1154 4.5005
R85228 VDD.n1676 VDD.n1236 4.5005
R85229 VDD.n1341 VDD.n1236 4.5005
R85230 VDD.n1342 VDD.n1236 4.5005
R85231 VDD.n1340 VDD.n1236 4.5005
R85232 VDD.n1344 VDD.n1236 4.5005
R85233 VDD.n1339 VDD.n1236 4.5005
R85234 VDD.n1345 VDD.n1236 4.5005
R85235 VDD.n1338 VDD.n1236 4.5005
R85236 VDD.n1347 VDD.n1236 4.5005
R85237 VDD.n1337 VDD.n1236 4.5005
R85238 VDD.n1348 VDD.n1236 4.5005
R85239 VDD.n1336 VDD.n1236 4.5005
R85240 VDD.n1350 VDD.n1236 4.5005
R85241 VDD.n1335 VDD.n1236 4.5005
R85242 VDD.n1351 VDD.n1236 4.5005
R85243 VDD.n1334 VDD.n1236 4.5005
R85244 VDD.n1353 VDD.n1236 4.5005
R85245 VDD.n1333 VDD.n1236 4.5005
R85246 VDD.n1354 VDD.n1236 4.5005
R85247 VDD.n1332 VDD.n1236 4.5005
R85248 VDD.n1356 VDD.n1236 4.5005
R85249 VDD.n1331 VDD.n1236 4.5005
R85250 VDD.n1357 VDD.n1236 4.5005
R85251 VDD.n1330 VDD.n1236 4.5005
R85252 VDD.n1359 VDD.n1236 4.5005
R85253 VDD.n1329 VDD.n1236 4.5005
R85254 VDD.n1360 VDD.n1236 4.5005
R85255 VDD.n1328 VDD.n1236 4.5005
R85256 VDD.n1362 VDD.n1236 4.5005
R85257 VDD.n1327 VDD.n1236 4.5005
R85258 VDD.n1363 VDD.n1236 4.5005
R85259 VDD.n1326 VDD.n1236 4.5005
R85260 VDD.n1365 VDD.n1236 4.5005
R85261 VDD.n1325 VDD.n1236 4.5005
R85262 VDD.n1366 VDD.n1236 4.5005
R85263 VDD.n1324 VDD.n1236 4.5005
R85264 VDD.n1368 VDD.n1236 4.5005
R85265 VDD.n1323 VDD.n1236 4.5005
R85266 VDD.n1369 VDD.n1236 4.5005
R85267 VDD.n1322 VDD.n1236 4.5005
R85268 VDD.n1371 VDD.n1236 4.5005
R85269 VDD.n1321 VDD.n1236 4.5005
R85270 VDD.n1372 VDD.n1236 4.5005
R85271 VDD.n1320 VDD.n1236 4.5005
R85272 VDD.n1374 VDD.n1236 4.5005
R85273 VDD.n1319 VDD.n1236 4.5005
R85274 VDD.n1375 VDD.n1236 4.5005
R85275 VDD.n1318 VDD.n1236 4.5005
R85276 VDD.n1376 VDD.n1236 4.5005
R85277 VDD.n1316 VDD.n1236 4.5005
R85278 VDD.n1377 VDD.n1236 4.5005
R85279 VDD.n1315 VDD.n1236 4.5005
R85280 VDD.n1378 VDD.n1236 4.5005
R85281 VDD.n1313 VDD.n1236 4.5005
R85282 VDD.n1379 VDD.n1236 4.5005
R85283 VDD.n1312 VDD.n1236 4.5005
R85284 VDD.n1380 VDD.n1236 4.5005
R85285 VDD.n1310 VDD.n1236 4.5005
R85286 VDD.n1381 VDD.n1236 4.5005
R85287 VDD.n1309 VDD.n1236 4.5005
R85288 VDD.n1382 VDD.n1236 4.5005
R85289 VDD.n1307 VDD.n1236 4.5005
R85290 VDD.n1383 VDD.n1236 4.5005
R85291 VDD.n1306 VDD.n1236 4.5005
R85292 VDD.n1384 VDD.n1236 4.5005
R85293 VDD.n1304 VDD.n1236 4.5005
R85294 VDD.n1385 VDD.n1236 4.5005
R85295 VDD.n1303 VDD.n1236 4.5005
R85296 VDD.n1386 VDD.n1236 4.5005
R85297 VDD.n1301 VDD.n1236 4.5005
R85298 VDD.n1387 VDD.n1236 4.5005
R85299 VDD.n1300 VDD.n1236 4.5005
R85300 VDD.n1388 VDD.n1236 4.5005
R85301 VDD.n1298 VDD.n1236 4.5005
R85302 VDD.n1389 VDD.n1236 4.5005
R85303 VDD.n1297 VDD.n1236 4.5005
R85304 VDD.n1390 VDD.n1236 4.5005
R85305 VDD.n1295 VDD.n1236 4.5005
R85306 VDD.n1391 VDD.n1236 4.5005
R85307 VDD.n1294 VDD.n1236 4.5005
R85308 VDD.n1392 VDD.n1236 4.5005
R85309 VDD.n1292 VDD.n1236 4.5005
R85310 VDD.n1393 VDD.n1236 4.5005
R85311 VDD.n1291 VDD.n1236 4.5005
R85312 VDD.n1394 VDD.n1236 4.5005
R85313 VDD.n1289 VDD.n1236 4.5005
R85314 VDD.n1395 VDD.n1236 4.5005
R85315 VDD.n1288 VDD.n1236 4.5005
R85316 VDD.n1396 VDD.n1236 4.5005
R85317 VDD.n1286 VDD.n1236 4.5005
R85318 VDD.n1397 VDD.n1236 4.5005
R85319 VDD.n1285 VDD.n1236 4.5005
R85320 VDD.n1398 VDD.n1236 4.5005
R85321 VDD.n1283 VDD.n1236 4.5005
R85322 VDD.n1399 VDD.n1236 4.5005
R85323 VDD.n1282 VDD.n1236 4.5005
R85324 VDD.n1400 VDD.n1236 4.5005
R85325 VDD.n1280 VDD.n1236 4.5005
R85326 VDD.n1401 VDD.n1236 4.5005
R85327 VDD.n1279 VDD.n1236 4.5005
R85328 VDD.n1402 VDD.n1236 4.5005
R85329 VDD.n1277 VDD.n1236 4.5005
R85330 VDD.n1403 VDD.n1236 4.5005
R85331 VDD.n1276 VDD.n1236 4.5005
R85332 VDD.n1404 VDD.n1236 4.5005
R85333 VDD.n1274 VDD.n1236 4.5005
R85334 VDD.n1405 VDD.n1236 4.5005
R85335 VDD.n1273 VDD.n1236 4.5005
R85336 VDD.n1406 VDD.n1236 4.5005
R85337 VDD.n1271 VDD.n1236 4.5005
R85338 VDD.n1407 VDD.n1236 4.5005
R85339 VDD.n1270 VDD.n1236 4.5005
R85340 VDD.n1408 VDD.n1236 4.5005
R85341 VDD.n1268 VDD.n1236 4.5005
R85342 VDD.n1409 VDD.n1236 4.5005
R85343 VDD.n1267 VDD.n1236 4.5005
R85344 VDD.n1410 VDD.n1236 4.5005
R85345 VDD.n1265 VDD.n1236 4.5005
R85346 VDD.n1411 VDD.n1236 4.5005
R85347 VDD.n1264 VDD.n1236 4.5005
R85348 VDD.n1412 VDD.n1236 4.5005
R85349 VDD.n1262 VDD.n1236 4.5005
R85350 VDD.n1413 VDD.n1236 4.5005
R85351 VDD.n1261 VDD.n1236 4.5005
R85352 VDD.n1414 VDD.n1236 4.5005
R85353 VDD.n1415 VDD.n1236 4.5005
R85354 VDD.n1674 VDD.n1236 4.5005
R85355 VDD.n1676 VDD.n1153 4.5005
R85356 VDD.n1341 VDD.n1153 4.5005
R85357 VDD.n1342 VDD.n1153 4.5005
R85358 VDD.n1340 VDD.n1153 4.5005
R85359 VDD.n1344 VDD.n1153 4.5005
R85360 VDD.n1339 VDD.n1153 4.5005
R85361 VDD.n1345 VDD.n1153 4.5005
R85362 VDD.n1338 VDD.n1153 4.5005
R85363 VDD.n1347 VDD.n1153 4.5005
R85364 VDD.n1337 VDD.n1153 4.5005
R85365 VDD.n1348 VDD.n1153 4.5005
R85366 VDD.n1336 VDD.n1153 4.5005
R85367 VDD.n1350 VDD.n1153 4.5005
R85368 VDD.n1335 VDD.n1153 4.5005
R85369 VDD.n1351 VDD.n1153 4.5005
R85370 VDD.n1334 VDD.n1153 4.5005
R85371 VDD.n1353 VDD.n1153 4.5005
R85372 VDD.n1333 VDD.n1153 4.5005
R85373 VDD.n1354 VDD.n1153 4.5005
R85374 VDD.n1332 VDD.n1153 4.5005
R85375 VDD.n1356 VDD.n1153 4.5005
R85376 VDD.n1331 VDD.n1153 4.5005
R85377 VDD.n1357 VDD.n1153 4.5005
R85378 VDD.n1330 VDD.n1153 4.5005
R85379 VDD.n1359 VDD.n1153 4.5005
R85380 VDD.n1329 VDD.n1153 4.5005
R85381 VDD.n1360 VDD.n1153 4.5005
R85382 VDD.n1328 VDD.n1153 4.5005
R85383 VDD.n1362 VDD.n1153 4.5005
R85384 VDD.n1327 VDD.n1153 4.5005
R85385 VDD.n1363 VDD.n1153 4.5005
R85386 VDD.n1326 VDD.n1153 4.5005
R85387 VDD.n1365 VDD.n1153 4.5005
R85388 VDD.n1325 VDD.n1153 4.5005
R85389 VDD.n1366 VDD.n1153 4.5005
R85390 VDD.n1324 VDD.n1153 4.5005
R85391 VDD.n1368 VDD.n1153 4.5005
R85392 VDD.n1323 VDD.n1153 4.5005
R85393 VDD.n1369 VDD.n1153 4.5005
R85394 VDD.n1322 VDD.n1153 4.5005
R85395 VDD.n1371 VDD.n1153 4.5005
R85396 VDD.n1321 VDD.n1153 4.5005
R85397 VDD.n1372 VDD.n1153 4.5005
R85398 VDD.n1320 VDD.n1153 4.5005
R85399 VDD.n1374 VDD.n1153 4.5005
R85400 VDD.n1319 VDD.n1153 4.5005
R85401 VDD.n1375 VDD.n1153 4.5005
R85402 VDD.n1318 VDD.n1153 4.5005
R85403 VDD.n1376 VDD.n1153 4.5005
R85404 VDD.n1316 VDD.n1153 4.5005
R85405 VDD.n1377 VDD.n1153 4.5005
R85406 VDD.n1315 VDD.n1153 4.5005
R85407 VDD.n1378 VDD.n1153 4.5005
R85408 VDD.n1313 VDD.n1153 4.5005
R85409 VDD.n1379 VDD.n1153 4.5005
R85410 VDD.n1312 VDD.n1153 4.5005
R85411 VDD.n1380 VDD.n1153 4.5005
R85412 VDD.n1310 VDD.n1153 4.5005
R85413 VDD.n1381 VDD.n1153 4.5005
R85414 VDD.n1309 VDD.n1153 4.5005
R85415 VDD.n1382 VDD.n1153 4.5005
R85416 VDD.n1307 VDD.n1153 4.5005
R85417 VDD.n1383 VDD.n1153 4.5005
R85418 VDD.n1306 VDD.n1153 4.5005
R85419 VDD.n1384 VDD.n1153 4.5005
R85420 VDD.n1304 VDD.n1153 4.5005
R85421 VDD.n1385 VDD.n1153 4.5005
R85422 VDD.n1303 VDD.n1153 4.5005
R85423 VDD.n1386 VDD.n1153 4.5005
R85424 VDD.n1301 VDD.n1153 4.5005
R85425 VDD.n1387 VDD.n1153 4.5005
R85426 VDD.n1300 VDD.n1153 4.5005
R85427 VDD.n1388 VDD.n1153 4.5005
R85428 VDD.n1298 VDD.n1153 4.5005
R85429 VDD.n1389 VDD.n1153 4.5005
R85430 VDD.n1297 VDD.n1153 4.5005
R85431 VDD.n1390 VDD.n1153 4.5005
R85432 VDD.n1295 VDD.n1153 4.5005
R85433 VDD.n1391 VDD.n1153 4.5005
R85434 VDD.n1294 VDD.n1153 4.5005
R85435 VDD.n1392 VDD.n1153 4.5005
R85436 VDD.n1292 VDD.n1153 4.5005
R85437 VDD.n1393 VDD.n1153 4.5005
R85438 VDD.n1291 VDD.n1153 4.5005
R85439 VDD.n1394 VDD.n1153 4.5005
R85440 VDD.n1289 VDD.n1153 4.5005
R85441 VDD.n1395 VDD.n1153 4.5005
R85442 VDD.n1288 VDD.n1153 4.5005
R85443 VDD.n1396 VDD.n1153 4.5005
R85444 VDD.n1286 VDD.n1153 4.5005
R85445 VDD.n1397 VDD.n1153 4.5005
R85446 VDD.n1285 VDD.n1153 4.5005
R85447 VDD.n1398 VDD.n1153 4.5005
R85448 VDD.n1283 VDD.n1153 4.5005
R85449 VDD.n1399 VDD.n1153 4.5005
R85450 VDD.n1282 VDD.n1153 4.5005
R85451 VDD.n1400 VDD.n1153 4.5005
R85452 VDD.n1280 VDD.n1153 4.5005
R85453 VDD.n1401 VDD.n1153 4.5005
R85454 VDD.n1279 VDD.n1153 4.5005
R85455 VDD.n1402 VDD.n1153 4.5005
R85456 VDD.n1277 VDD.n1153 4.5005
R85457 VDD.n1403 VDD.n1153 4.5005
R85458 VDD.n1276 VDD.n1153 4.5005
R85459 VDD.n1404 VDD.n1153 4.5005
R85460 VDD.n1274 VDD.n1153 4.5005
R85461 VDD.n1405 VDD.n1153 4.5005
R85462 VDD.n1273 VDD.n1153 4.5005
R85463 VDD.n1406 VDD.n1153 4.5005
R85464 VDD.n1271 VDD.n1153 4.5005
R85465 VDD.n1407 VDD.n1153 4.5005
R85466 VDD.n1270 VDD.n1153 4.5005
R85467 VDD.n1408 VDD.n1153 4.5005
R85468 VDD.n1268 VDD.n1153 4.5005
R85469 VDD.n1409 VDD.n1153 4.5005
R85470 VDD.n1267 VDD.n1153 4.5005
R85471 VDD.n1410 VDD.n1153 4.5005
R85472 VDD.n1265 VDD.n1153 4.5005
R85473 VDD.n1411 VDD.n1153 4.5005
R85474 VDD.n1264 VDD.n1153 4.5005
R85475 VDD.n1412 VDD.n1153 4.5005
R85476 VDD.n1262 VDD.n1153 4.5005
R85477 VDD.n1413 VDD.n1153 4.5005
R85478 VDD.n1261 VDD.n1153 4.5005
R85479 VDD.n1414 VDD.n1153 4.5005
R85480 VDD.n1415 VDD.n1153 4.5005
R85481 VDD.n1674 VDD.n1153 4.5005
R85482 VDD.n1676 VDD.n1237 4.5005
R85483 VDD.n1341 VDD.n1237 4.5005
R85484 VDD.n1342 VDD.n1237 4.5005
R85485 VDD.n1340 VDD.n1237 4.5005
R85486 VDD.n1344 VDD.n1237 4.5005
R85487 VDD.n1339 VDD.n1237 4.5005
R85488 VDD.n1345 VDD.n1237 4.5005
R85489 VDD.n1338 VDD.n1237 4.5005
R85490 VDD.n1347 VDD.n1237 4.5005
R85491 VDD.n1337 VDD.n1237 4.5005
R85492 VDD.n1348 VDD.n1237 4.5005
R85493 VDD.n1336 VDD.n1237 4.5005
R85494 VDD.n1350 VDD.n1237 4.5005
R85495 VDD.n1335 VDD.n1237 4.5005
R85496 VDD.n1351 VDD.n1237 4.5005
R85497 VDD.n1334 VDD.n1237 4.5005
R85498 VDD.n1353 VDD.n1237 4.5005
R85499 VDD.n1333 VDD.n1237 4.5005
R85500 VDD.n1354 VDD.n1237 4.5005
R85501 VDD.n1332 VDD.n1237 4.5005
R85502 VDD.n1356 VDD.n1237 4.5005
R85503 VDD.n1331 VDD.n1237 4.5005
R85504 VDD.n1357 VDD.n1237 4.5005
R85505 VDD.n1330 VDD.n1237 4.5005
R85506 VDD.n1359 VDD.n1237 4.5005
R85507 VDD.n1329 VDD.n1237 4.5005
R85508 VDD.n1360 VDD.n1237 4.5005
R85509 VDD.n1328 VDD.n1237 4.5005
R85510 VDD.n1362 VDD.n1237 4.5005
R85511 VDD.n1327 VDD.n1237 4.5005
R85512 VDD.n1363 VDD.n1237 4.5005
R85513 VDD.n1326 VDD.n1237 4.5005
R85514 VDD.n1365 VDD.n1237 4.5005
R85515 VDD.n1325 VDD.n1237 4.5005
R85516 VDD.n1366 VDD.n1237 4.5005
R85517 VDD.n1324 VDD.n1237 4.5005
R85518 VDD.n1368 VDD.n1237 4.5005
R85519 VDD.n1323 VDD.n1237 4.5005
R85520 VDD.n1369 VDD.n1237 4.5005
R85521 VDD.n1322 VDD.n1237 4.5005
R85522 VDD.n1371 VDD.n1237 4.5005
R85523 VDD.n1321 VDD.n1237 4.5005
R85524 VDD.n1372 VDD.n1237 4.5005
R85525 VDD.n1320 VDD.n1237 4.5005
R85526 VDD.n1374 VDD.n1237 4.5005
R85527 VDD.n1319 VDD.n1237 4.5005
R85528 VDD.n1375 VDD.n1237 4.5005
R85529 VDD.n1318 VDD.n1237 4.5005
R85530 VDD.n1376 VDD.n1237 4.5005
R85531 VDD.n1316 VDD.n1237 4.5005
R85532 VDD.n1377 VDD.n1237 4.5005
R85533 VDD.n1315 VDD.n1237 4.5005
R85534 VDD.n1378 VDD.n1237 4.5005
R85535 VDD.n1313 VDD.n1237 4.5005
R85536 VDD.n1379 VDD.n1237 4.5005
R85537 VDD.n1312 VDD.n1237 4.5005
R85538 VDD.n1380 VDD.n1237 4.5005
R85539 VDD.n1310 VDD.n1237 4.5005
R85540 VDD.n1381 VDD.n1237 4.5005
R85541 VDD.n1309 VDD.n1237 4.5005
R85542 VDD.n1382 VDD.n1237 4.5005
R85543 VDD.n1307 VDD.n1237 4.5005
R85544 VDD.n1383 VDD.n1237 4.5005
R85545 VDD.n1306 VDD.n1237 4.5005
R85546 VDD.n1384 VDD.n1237 4.5005
R85547 VDD.n1304 VDD.n1237 4.5005
R85548 VDD.n1385 VDD.n1237 4.5005
R85549 VDD.n1303 VDD.n1237 4.5005
R85550 VDD.n1386 VDD.n1237 4.5005
R85551 VDD.n1301 VDD.n1237 4.5005
R85552 VDD.n1387 VDD.n1237 4.5005
R85553 VDD.n1300 VDD.n1237 4.5005
R85554 VDD.n1388 VDD.n1237 4.5005
R85555 VDD.n1298 VDD.n1237 4.5005
R85556 VDD.n1389 VDD.n1237 4.5005
R85557 VDD.n1297 VDD.n1237 4.5005
R85558 VDD.n1390 VDD.n1237 4.5005
R85559 VDD.n1295 VDD.n1237 4.5005
R85560 VDD.n1391 VDD.n1237 4.5005
R85561 VDD.n1294 VDD.n1237 4.5005
R85562 VDD.n1392 VDD.n1237 4.5005
R85563 VDD.n1292 VDD.n1237 4.5005
R85564 VDD.n1393 VDD.n1237 4.5005
R85565 VDD.n1291 VDD.n1237 4.5005
R85566 VDD.n1394 VDD.n1237 4.5005
R85567 VDD.n1289 VDD.n1237 4.5005
R85568 VDD.n1395 VDD.n1237 4.5005
R85569 VDD.n1288 VDD.n1237 4.5005
R85570 VDD.n1396 VDD.n1237 4.5005
R85571 VDD.n1286 VDD.n1237 4.5005
R85572 VDD.n1397 VDD.n1237 4.5005
R85573 VDD.n1285 VDD.n1237 4.5005
R85574 VDD.n1398 VDD.n1237 4.5005
R85575 VDD.n1283 VDD.n1237 4.5005
R85576 VDD.n1399 VDD.n1237 4.5005
R85577 VDD.n1282 VDD.n1237 4.5005
R85578 VDD.n1400 VDD.n1237 4.5005
R85579 VDD.n1280 VDD.n1237 4.5005
R85580 VDD.n1401 VDD.n1237 4.5005
R85581 VDD.n1279 VDD.n1237 4.5005
R85582 VDD.n1402 VDD.n1237 4.5005
R85583 VDD.n1277 VDD.n1237 4.5005
R85584 VDD.n1403 VDD.n1237 4.5005
R85585 VDD.n1276 VDD.n1237 4.5005
R85586 VDD.n1404 VDD.n1237 4.5005
R85587 VDD.n1274 VDD.n1237 4.5005
R85588 VDD.n1405 VDD.n1237 4.5005
R85589 VDD.n1273 VDD.n1237 4.5005
R85590 VDD.n1406 VDD.n1237 4.5005
R85591 VDD.n1271 VDD.n1237 4.5005
R85592 VDD.n1407 VDD.n1237 4.5005
R85593 VDD.n1270 VDD.n1237 4.5005
R85594 VDD.n1408 VDD.n1237 4.5005
R85595 VDD.n1268 VDD.n1237 4.5005
R85596 VDD.n1409 VDD.n1237 4.5005
R85597 VDD.n1267 VDD.n1237 4.5005
R85598 VDD.n1410 VDD.n1237 4.5005
R85599 VDD.n1265 VDD.n1237 4.5005
R85600 VDD.n1411 VDD.n1237 4.5005
R85601 VDD.n1264 VDD.n1237 4.5005
R85602 VDD.n1412 VDD.n1237 4.5005
R85603 VDD.n1262 VDD.n1237 4.5005
R85604 VDD.n1413 VDD.n1237 4.5005
R85605 VDD.n1261 VDD.n1237 4.5005
R85606 VDD.n1414 VDD.n1237 4.5005
R85607 VDD.n1415 VDD.n1237 4.5005
R85608 VDD.n1674 VDD.n1237 4.5005
R85609 VDD.n1676 VDD.n1152 4.5005
R85610 VDD.n1341 VDD.n1152 4.5005
R85611 VDD.n1342 VDD.n1152 4.5005
R85612 VDD.n1340 VDD.n1152 4.5005
R85613 VDD.n1344 VDD.n1152 4.5005
R85614 VDD.n1339 VDD.n1152 4.5005
R85615 VDD.n1345 VDD.n1152 4.5005
R85616 VDD.n1338 VDD.n1152 4.5005
R85617 VDD.n1347 VDD.n1152 4.5005
R85618 VDD.n1337 VDD.n1152 4.5005
R85619 VDD.n1348 VDD.n1152 4.5005
R85620 VDD.n1336 VDD.n1152 4.5005
R85621 VDD.n1350 VDD.n1152 4.5005
R85622 VDD.n1335 VDD.n1152 4.5005
R85623 VDD.n1351 VDD.n1152 4.5005
R85624 VDD.n1334 VDD.n1152 4.5005
R85625 VDD.n1353 VDD.n1152 4.5005
R85626 VDD.n1333 VDD.n1152 4.5005
R85627 VDD.n1354 VDD.n1152 4.5005
R85628 VDD.n1332 VDD.n1152 4.5005
R85629 VDD.n1356 VDD.n1152 4.5005
R85630 VDD.n1331 VDD.n1152 4.5005
R85631 VDD.n1357 VDD.n1152 4.5005
R85632 VDD.n1330 VDD.n1152 4.5005
R85633 VDD.n1359 VDD.n1152 4.5005
R85634 VDD.n1329 VDD.n1152 4.5005
R85635 VDD.n1360 VDD.n1152 4.5005
R85636 VDD.n1328 VDD.n1152 4.5005
R85637 VDD.n1362 VDD.n1152 4.5005
R85638 VDD.n1327 VDD.n1152 4.5005
R85639 VDD.n1363 VDD.n1152 4.5005
R85640 VDD.n1326 VDD.n1152 4.5005
R85641 VDD.n1365 VDD.n1152 4.5005
R85642 VDD.n1325 VDD.n1152 4.5005
R85643 VDD.n1366 VDD.n1152 4.5005
R85644 VDD.n1324 VDD.n1152 4.5005
R85645 VDD.n1368 VDD.n1152 4.5005
R85646 VDD.n1323 VDD.n1152 4.5005
R85647 VDD.n1369 VDD.n1152 4.5005
R85648 VDD.n1322 VDD.n1152 4.5005
R85649 VDD.n1371 VDD.n1152 4.5005
R85650 VDD.n1321 VDD.n1152 4.5005
R85651 VDD.n1372 VDD.n1152 4.5005
R85652 VDD.n1320 VDD.n1152 4.5005
R85653 VDD.n1374 VDD.n1152 4.5005
R85654 VDD.n1319 VDD.n1152 4.5005
R85655 VDD.n1375 VDD.n1152 4.5005
R85656 VDD.n1318 VDD.n1152 4.5005
R85657 VDD.n1376 VDD.n1152 4.5005
R85658 VDD.n1316 VDD.n1152 4.5005
R85659 VDD.n1377 VDD.n1152 4.5005
R85660 VDD.n1315 VDD.n1152 4.5005
R85661 VDD.n1378 VDD.n1152 4.5005
R85662 VDD.n1313 VDD.n1152 4.5005
R85663 VDD.n1379 VDD.n1152 4.5005
R85664 VDD.n1312 VDD.n1152 4.5005
R85665 VDD.n1380 VDD.n1152 4.5005
R85666 VDD.n1310 VDD.n1152 4.5005
R85667 VDD.n1381 VDD.n1152 4.5005
R85668 VDD.n1309 VDD.n1152 4.5005
R85669 VDD.n1382 VDD.n1152 4.5005
R85670 VDD.n1307 VDD.n1152 4.5005
R85671 VDD.n1383 VDD.n1152 4.5005
R85672 VDD.n1306 VDD.n1152 4.5005
R85673 VDD.n1384 VDD.n1152 4.5005
R85674 VDD.n1304 VDD.n1152 4.5005
R85675 VDD.n1385 VDD.n1152 4.5005
R85676 VDD.n1303 VDD.n1152 4.5005
R85677 VDD.n1386 VDD.n1152 4.5005
R85678 VDD.n1301 VDD.n1152 4.5005
R85679 VDD.n1387 VDD.n1152 4.5005
R85680 VDD.n1300 VDD.n1152 4.5005
R85681 VDD.n1388 VDD.n1152 4.5005
R85682 VDD.n1298 VDD.n1152 4.5005
R85683 VDD.n1389 VDD.n1152 4.5005
R85684 VDD.n1297 VDD.n1152 4.5005
R85685 VDD.n1390 VDD.n1152 4.5005
R85686 VDD.n1295 VDD.n1152 4.5005
R85687 VDD.n1391 VDD.n1152 4.5005
R85688 VDD.n1294 VDD.n1152 4.5005
R85689 VDD.n1392 VDD.n1152 4.5005
R85690 VDD.n1292 VDD.n1152 4.5005
R85691 VDD.n1393 VDD.n1152 4.5005
R85692 VDD.n1291 VDD.n1152 4.5005
R85693 VDD.n1394 VDD.n1152 4.5005
R85694 VDD.n1289 VDD.n1152 4.5005
R85695 VDD.n1395 VDD.n1152 4.5005
R85696 VDD.n1288 VDD.n1152 4.5005
R85697 VDD.n1396 VDD.n1152 4.5005
R85698 VDD.n1286 VDD.n1152 4.5005
R85699 VDD.n1397 VDD.n1152 4.5005
R85700 VDD.n1285 VDD.n1152 4.5005
R85701 VDD.n1398 VDD.n1152 4.5005
R85702 VDD.n1283 VDD.n1152 4.5005
R85703 VDD.n1399 VDD.n1152 4.5005
R85704 VDD.n1282 VDD.n1152 4.5005
R85705 VDD.n1400 VDD.n1152 4.5005
R85706 VDD.n1280 VDD.n1152 4.5005
R85707 VDD.n1401 VDD.n1152 4.5005
R85708 VDD.n1279 VDD.n1152 4.5005
R85709 VDD.n1402 VDD.n1152 4.5005
R85710 VDD.n1277 VDD.n1152 4.5005
R85711 VDD.n1403 VDD.n1152 4.5005
R85712 VDD.n1276 VDD.n1152 4.5005
R85713 VDD.n1404 VDD.n1152 4.5005
R85714 VDD.n1274 VDD.n1152 4.5005
R85715 VDD.n1405 VDD.n1152 4.5005
R85716 VDD.n1273 VDD.n1152 4.5005
R85717 VDD.n1406 VDD.n1152 4.5005
R85718 VDD.n1271 VDD.n1152 4.5005
R85719 VDD.n1407 VDD.n1152 4.5005
R85720 VDD.n1270 VDD.n1152 4.5005
R85721 VDD.n1408 VDD.n1152 4.5005
R85722 VDD.n1268 VDD.n1152 4.5005
R85723 VDD.n1409 VDD.n1152 4.5005
R85724 VDD.n1267 VDD.n1152 4.5005
R85725 VDD.n1410 VDD.n1152 4.5005
R85726 VDD.n1265 VDD.n1152 4.5005
R85727 VDD.n1411 VDD.n1152 4.5005
R85728 VDD.n1264 VDD.n1152 4.5005
R85729 VDD.n1412 VDD.n1152 4.5005
R85730 VDD.n1262 VDD.n1152 4.5005
R85731 VDD.n1413 VDD.n1152 4.5005
R85732 VDD.n1261 VDD.n1152 4.5005
R85733 VDD.n1414 VDD.n1152 4.5005
R85734 VDD.n1415 VDD.n1152 4.5005
R85735 VDD.n1674 VDD.n1152 4.5005
R85736 VDD.n1676 VDD.n1238 4.5005
R85737 VDD.n1341 VDD.n1238 4.5005
R85738 VDD.n1342 VDD.n1238 4.5005
R85739 VDD.n1340 VDD.n1238 4.5005
R85740 VDD.n1344 VDD.n1238 4.5005
R85741 VDD.n1339 VDD.n1238 4.5005
R85742 VDD.n1345 VDD.n1238 4.5005
R85743 VDD.n1338 VDD.n1238 4.5005
R85744 VDD.n1347 VDD.n1238 4.5005
R85745 VDD.n1337 VDD.n1238 4.5005
R85746 VDD.n1348 VDD.n1238 4.5005
R85747 VDD.n1336 VDD.n1238 4.5005
R85748 VDD.n1350 VDD.n1238 4.5005
R85749 VDD.n1335 VDD.n1238 4.5005
R85750 VDD.n1351 VDD.n1238 4.5005
R85751 VDD.n1334 VDD.n1238 4.5005
R85752 VDD.n1353 VDD.n1238 4.5005
R85753 VDD.n1333 VDD.n1238 4.5005
R85754 VDD.n1354 VDD.n1238 4.5005
R85755 VDD.n1332 VDD.n1238 4.5005
R85756 VDD.n1356 VDD.n1238 4.5005
R85757 VDD.n1331 VDD.n1238 4.5005
R85758 VDD.n1357 VDD.n1238 4.5005
R85759 VDD.n1330 VDD.n1238 4.5005
R85760 VDD.n1359 VDD.n1238 4.5005
R85761 VDD.n1329 VDD.n1238 4.5005
R85762 VDD.n1360 VDD.n1238 4.5005
R85763 VDD.n1328 VDD.n1238 4.5005
R85764 VDD.n1362 VDD.n1238 4.5005
R85765 VDD.n1327 VDD.n1238 4.5005
R85766 VDD.n1363 VDD.n1238 4.5005
R85767 VDD.n1326 VDD.n1238 4.5005
R85768 VDD.n1365 VDD.n1238 4.5005
R85769 VDD.n1325 VDD.n1238 4.5005
R85770 VDD.n1366 VDD.n1238 4.5005
R85771 VDD.n1324 VDD.n1238 4.5005
R85772 VDD.n1368 VDD.n1238 4.5005
R85773 VDD.n1323 VDD.n1238 4.5005
R85774 VDD.n1369 VDD.n1238 4.5005
R85775 VDD.n1322 VDD.n1238 4.5005
R85776 VDD.n1371 VDD.n1238 4.5005
R85777 VDD.n1321 VDD.n1238 4.5005
R85778 VDD.n1372 VDD.n1238 4.5005
R85779 VDD.n1320 VDD.n1238 4.5005
R85780 VDD.n1374 VDD.n1238 4.5005
R85781 VDD.n1319 VDD.n1238 4.5005
R85782 VDD.n1375 VDD.n1238 4.5005
R85783 VDD.n1318 VDD.n1238 4.5005
R85784 VDD.n1376 VDD.n1238 4.5005
R85785 VDD.n1316 VDD.n1238 4.5005
R85786 VDD.n1377 VDD.n1238 4.5005
R85787 VDD.n1315 VDD.n1238 4.5005
R85788 VDD.n1378 VDD.n1238 4.5005
R85789 VDD.n1313 VDD.n1238 4.5005
R85790 VDD.n1379 VDD.n1238 4.5005
R85791 VDD.n1312 VDD.n1238 4.5005
R85792 VDD.n1380 VDD.n1238 4.5005
R85793 VDD.n1310 VDD.n1238 4.5005
R85794 VDD.n1381 VDD.n1238 4.5005
R85795 VDD.n1309 VDD.n1238 4.5005
R85796 VDD.n1382 VDD.n1238 4.5005
R85797 VDD.n1307 VDD.n1238 4.5005
R85798 VDD.n1383 VDD.n1238 4.5005
R85799 VDD.n1306 VDD.n1238 4.5005
R85800 VDD.n1384 VDD.n1238 4.5005
R85801 VDD.n1304 VDD.n1238 4.5005
R85802 VDD.n1385 VDD.n1238 4.5005
R85803 VDD.n1303 VDD.n1238 4.5005
R85804 VDD.n1386 VDD.n1238 4.5005
R85805 VDD.n1301 VDD.n1238 4.5005
R85806 VDD.n1387 VDD.n1238 4.5005
R85807 VDD.n1300 VDD.n1238 4.5005
R85808 VDD.n1388 VDD.n1238 4.5005
R85809 VDD.n1298 VDD.n1238 4.5005
R85810 VDD.n1389 VDD.n1238 4.5005
R85811 VDD.n1297 VDD.n1238 4.5005
R85812 VDD.n1390 VDD.n1238 4.5005
R85813 VDD.n1295 VDD.n1238 4.5005
R85814 VDD.n1391 VDD.n1238 4.5005
R85815 VDD.n1294 VDD.n1238 4.5005
R85816 VDD.n1392 VDD.n1238 4.5005
R85817 VDD.n1292 VDD.n1238 4.5005
R85818 VDD.n1393 VDD.n1238 4.5005
R85819 VDD.n1291 VDD.n1238 4.5005
R85820 VDD.n1394 VDD.n1238 4.5005
R85821 VDD.n1289 VDD.n1238 4.5005
R85822 VDD.n1395 VDD.n1238 4.5005
R85823 VDD.n1288 VDD.n1238 4.5005
R85824 VDD.n1396 VDD.n1238 4.5005
R85825 VDD.n1286 VDD.n1238 4.5005
R85826 VDD.n1397 VDD.n1238 4.5005
R85827 VDD.n1285 VDD.n1238 4.5005
R85828 VDD.n1398 VDD.n1238 4.5005
R85829 VDD.n1283 VDD.n1238 4.5005
R85830 VDD.n1399 VDD.n1238 4.5005
R85831 VDD.n1282 VDD.n1238 4.5005
R85832 VDD.n1400 VDD.n1238 4.5005
R85833 VDD.n1280 VDD.n1238 4.5005
R85834 VDD.n1401 VDD.n1238 4.5005
R85835 VDD.n1279 VDD.n1238 4.5005
R85836 VDD.n1402 VDD.n1238 4.5005
R85837 VDD.n1277 VDD.n1238 4.5005
R85838 VDD.n1403 VDD.n1238 4.5005
R85839 VDD.n1276 VDD.n1238 4.5005
R85840 VDD.n1404 VDD.n1238 4.5005
R85841 VDD.n1274 VDD.n1238 4.5005
R85842 VDD.n1405 VDD.n1238 4.5005
R85843 VDD.n1273 VDD.n1238 4.5005
R85844 VDD.n1406 VDD.n1238 4.5005
R85845 VDD.n1271 VDD.n1238 4.5005
R85846 VDD.n1407 VDD.n1238 4.5005
R85847 VDD.n1270 VDD.n1238 4.5005
R85848 VDD.n1408 VDD.n1238 4.5005
R85849 VDD.n1268 VDD.n1238 4.5005
R85850 VDD.n1409 VDD.n1238 4.5005
R85851 VDD.n1267 VDD.n1238 4.5005
R85852 VDD.n1410 VDD.n1238 4.5005
R85853 VDD.n1265 VDD.n1238 4.5005
R85854 VDD.n1411 VDD.n1238 4.5005
R85855 VDD.n1264 VDD.n1238 4.5005
R85856 VDD.n1412 VDD.n1238 4.5005
R85857 VDD.n1262 VDD.n1238 4.5005
R85858 VDD.n1413 VDD.n1238 4.5005
R85859 VDD.n1261 VDD.n1238 4.5005
R85860 VDD.n1414 VDD.n1238 4.5005
R85861 VDD.n1415 VDD.n1238 4.5005
R85862 VDD.n1674 VDD.n1238 4.5005
R85863 VDD.n1676 VDD.n1151 4.5005
R85864 VDD.n1341 VDD.n1151 4.5005
R85865 VDD.n1342 VDD.n1151 4.5005
R85866 VDD.n1340 VDD.n1151 4.5005
R85867 VDD.n1344 VDD.n1151 4.5005
R85868 VDD.n1339 VDD.n1151 4.5005
R85869 VDD.n1345 VDD.n1151 4.5005
R85870 VDD.n1338 VDD.n1151 4.5005
R85871 VDD.n1347 VDD.n1151 4.5005
R85872 VDD.n1337 VDD.n1151 4.5005
R85873 VDD.n1348 VDD.n1151 4.5005
R85874 VDD.n1336 VDD.n1151 4.5005
R85875 VDD.n1350 VDD.n1151 4.5005
R85876 VDD.n1335 VDD.n1151 4.5005
R85877 VDD.n1351 VDD.n1151 4.5005
R85878 VDD.n1334 VDD.n1151 4.5005
R85879 VDD.n1353 VDD.n1151 4.5005
R85880 VDD.n1333 VDD.n1151 4.5005
R85881 VDD.n1354 VDD.n1151 4.5005
R85882 VDD.n1332 VDD.n1151 4.5005
R85883 VDD.n1356 VDD.n1151 4.5005
R85884 VDD.n1331 VDD.n1151 4.5005
R85885 VDD.n1357 VDD.n1151 4.5005
R85886 VDD.n1330 VDD.n1151 4.5005
R85887 VDD.n1359 VDD.n1151 4.5005
R85888 VDD.n1329 VDD.n1151 4.5005
R85889 VDD.n1360 VDD.n1151 4.5005
R85890 VDD.n1328 VDD.n1151 4.5005
R85891 VDD.n1362 VDD.n1151 4.5005
R85892 VDD.n1327 VDD.n1151 4.5005
R85893 VDD.n1363 VDD.n1151 4.5005
R85894 VDD.n1326 VDD.n1151 4.5005
R85895 VDD.n1365 VDD.n1151 4.5005
R85896 VDD.n1325 VDD.n1151 4.5005
R85897 VDD.n1366 VDD.n1151 4.5005
R85898 VDD.n1324 VDD.n1151 4.5005
R85899 VDD.n1368 VDD.n1151 4.5005
R85900 VDD.n1323 VDD.n1151 4.5005
R85901 VDD.n1369 VDD.n1151 4.5005
R85902 VDD.n1322 VDD.n1151 4.5005
R85903 VDD.n1371 VDD.n1151 4.5005
R85904 VDD.n1321 VDD.n1151 4.5005
R85905 VDD.n1372 VDD.n1151 4.5005
R85906 VDD.n1320 VDD.n1151 4.5005
R85907 VDD.n1374 VDD.n1151 4.5005
R85908 VDD.n1319 VDD.n1151 4.5005
R85909 VDD.n1375 VDD.n1151 4.5005
R85910 VDD.n1318 VDD.n1151 4.5005
R85911 VDD.n1376 VDD.n1151 4.5005
R85912 VDD.n1316 VDD.n1151 4.5005
R85913 VDD.n1377 VDD.n1151 4.5005
R85914 VDD.n1315 VDD.n1151 4.5005
R85915 VDD.n1378 VDD.n1151 4.5005
R85916 VDD.n1313 VDD.n1151 4.5005
R85917 VDD.n1379 VDD.n1151 4.5005
R85918 VDD.n1312 VDD.n1151 4.5005
R85919 VDD.n1380 VDD.n1151 4.5005
R85920 VDD.n1310 VDD.n1151 4.5005
R85921 VDD.n1381 VDD.n1151 4.5005
R85922 VDD.n1309 VDD.n1151 4.5005
R85923 VDD.n1382 VDD.n1151 4.5005
R85924 VDD.n1307 VDD.n1151 4.5005
R85925 VDD.n1383 VDD.n1151 4.5005
R85926 VDD.n1306 VDD.n1151 4.5005
R85927 VDD.n1384 VDD.n1151 4.5005
R85928 VDD.n1304 VDD.n1151 4.5005
R85929 VDD.n1385 VDD.n1151 4.5005
R85930 VDD.n1303 VDD.n1151 4.5005
R85931 VDD.n1386 VDD.n1151 4.5005
R85932 VDD.n1301 VDD.n1151 4.5005
R85933 VDD.n1387 VDD.n1151 4.5005
R85934 VDD.n1300 VDD.n1151 4.5005
R85935 VDD.n1388 VDD.n1151 4.5005
R85936 VDD.n1298 VDD.n1151 4.5005
R85937 VDD.n1389 VDD.n1151 4.5005
R85938 VDD.n1297 VDD.n1151 4.5005
R85939 VDD.n1390 VDD.n1151 4.5005
R85940 VDD.n1295 VDD.n1151 4.5005
R85941 VDD.n1391 VDD.n1151 4.5005
R85942 VDD.n1294 VDD.n1151 4.5005
R85943 VDD.n1392 VDD.n1151 4.5005
R85944 VDD.n1292 VDD.n1151 4.5005
R85945 VDD.n1393 VDD.n1151 4.5005
R85946 VDD.n1291 VDD.n1151 4.5005
R85947 VDD.n1394 VDD.n1151 4.5005
R85948 VDD.n1289 VDD.n1151 4.5005
R85949 VDD.n1395 VDD.n1151 4.5005
R85950 VDD.n1288 VDD.n1151 4.5005
R85951 VDD.n1396 VDD.n1151 4.5005
R85952 VDD.n1286 VDD.n1151 4.5005
R85953 VDD.n1397 VDD.n1151 4.5005
R85954 VDD.n1285 VDD.n1151 4.5005
R85955 VDD.n1398 VDD.n1151 4.5005
R85956 VDD.n1283 VDD.n1151 4.5005
R85957 VDD.n1399 VDD.n1151 4.5005
R85958 VDD.n1282 VDD.n1151 4.5005
R85959 VDD.n1400 VDD.n1151 4.5005
R85960 VDD.n1280 VDD.n1151 4.5005
R85961 VDD.n1401 VDD.n1151 4.5005
R85962 VDD.n1279 VDD.n1151 4.5005
R85963 VDD.n1402 VDD.n1151 4.5005
R85964 VDD.n1277 VDD.n1151 4.5005
R85965 VDD.n1403 VDD.n1151 4.5005
R85966 VDD.n1276 VDD.n1151 4.5005
R85967 VDD.n1404 VDD.n1151 4.5005
R85968 VDD.n1274 VDD.n1151 4.5005
R85969 VDD.n1405 VDD.n1151 4.5005
R85970 VDD.n1273 VDD.n1151 4.5005
R85971 VDD.n1406 VDD.n1151 4.5005
R85972 VDD.n1271 VDD.n1151 4.5005
R85973 VDD.n1407 VDD.n1151 4.5005
R85974 VDD.n1270 VDD.n1151 4.5005
R85975 VDD.n1408 VDD.n1151 4.5005
R85976 VDD.n1268 VDD.n1151 4.5005
R85977 VDD.n1409 VDD.n1151 4.5005
R85978 VDD.n1267 VDD.n1151 4.5005
R85979 VDD.n1410 VDD.n1151 4.5005
R85980 VDD.n1265 VDD.n1151 4.5005
R85981 VDD.n1411 VDD.n1151 4.5005
R85982 VDD.n1264 VDD.n1151 4.5005
R85983 VDD.n1412 VDD.n1151 4.5005
R85984 VDD.n1262 VDD.n1151 4.5005
R85985 VDD.n1413 VDD.n1151 4.5005
R85986 VDD.n1261 VDD.n1151 4.5005
R85987 VDD.n1414 VDD.n1151 4.5005
R85988 VDD.n1415 VDD.n1151 4.5005
R85989 VDD.n1674 VDD.n1151 4.5005
R85990 VDD.n1676 VDD.n1239 4.5005
R85991 VDD.n1341 VDD.n1239 4.5005
R85992 VDD.n1342 VDD.n1239 4.5005
R85993 VDD.n1340 VDD.n1239 4.5005
R85994 VDD.n1344 VDD.n1239 4.5005
R85995 VDD.n1339 VDD.n1239 4.5005
R85996 VDD.n1345 VDD.n1239 4.5005
R85997 VDD.n1338 VDD.n1239 4.5005
R85998 VDD.n1347 VDD.n1239 4.5005
R85999 VDD.n1337 VDD.n1239 4.5005
R86000 VDD.n1348 VDD.n1239 4.5005
R86001 VDD.n1336 VDD.n1239 4.5005
R86002 VDD.n1350 VDD.n1239 4.5005
R86003 VDD.n1335 VDD.n1239 4.5005
R86004 VDD.n1351 VDD.n1239 4.5005
R86005 VDD.n1334 VDD.n1239 4.5005
R86006 VDD.n1353 VDD.n1239 4.5005
R86007 VDD.n1333 VDD.n1239 4.5005
R86008 VDD.n1354 VDD.n1239 4.5005
R86009 VDD.n1332 VDD.n1239 4.5005
R86010 VDD.n1356 VDD.n1239 4.5005
R86011 VDD.n1331 VDD.n1239 4.5005
R86012 VDD.n1357 VDD.n1239 4.5005
R86013 VDD.n1330 VDD.n1239 4.5005
R86014 VDD.n1359 VDD.n1239 4.5005
R86015 VDD.n1329 VDD.n1239 4.5005
R86016 VDD.n1360 VDD.n1239 4.5005
R86017 VDD.n1328 VDD.n1239 4.5005
R86018 VDD.n1362 VDD.n1239 4.5005
R86019 VDD.n1327 VDD.n1239 4.5005
R86020 VDD.n1363 VDD.n1239 4.5005
R86021 VDD.n1326 VDD.n1239 4.5005
R86022 VDD.n1365 VDD.n1239 4.5005
R86023 VDD.n1325 VDD.n1239 4.5005
R86024 VDD.n1366 VDD.n1239 4.5005
R86025 VDD.n1324 VDD.n1239 4.5005
R86026 VDD.n1368 VDD.n1239 4.5005
R86027 VDD.n1323 VDD.n1239 4.5005
R86028 VDD.n1369 VDD.n1239 4.5005
R86029 VDD.n1322 VDD.n1239 4.5005
R86030 VDD.n1371 VDD.n1239 4.5005
R86031 VDD.n1321 VDD.n1239 4.5005
R86032 VDD.n1372 VDD.n1239 4.5005
R86033 VDD.n1320 VDD.n1239 4.5005
R86034 VDD.n1374 VDD.n1239 4.5005
R86035 VDD.n1319 VDD.n1239 4.5005
R86036 VDD.n1375 VDD.n1239 4.5005
R86037 VDD.n1318 VDD.n1239 4.5005
R86038 VDD.n1376 VDD.n1239 4.5005
R86039 VDD.n1316 VDD.n1239 4.5005
R86040 VDD.n1377 VDD.n1239 4.5005
R86041 VDD.n1315 VDD.n1239 4.5005
R86042 VDD.n1378 VDD.n1239 4.5005
R86043 VDD.n1313 VDD.n1239 4.5005
R86044 VDD.n1379 VDD.n1239 4.5005
R86045 VDD.n1312 VDD.n1239 4.5005
R86046 VDD.n1380 VDD.n1239 4.5005
R86047 VDD.n1310 VDD.n1239 4.5005
R86048 VDD.n1381 VDD.n1239 4.5005
R86049 VDD.n1309 VDD.n1239 4.5005
R86050 VDD.n1382 VDD.n1239 4.5005
R86051 VDD.n1307 VDD.n1239 4.5005
R86052 VDD.n1383 VDD.n1239 4.5005
R86053 VDD.n1306 VDD.n1239 4.5005
R86054 VDD.n1384 VDD.n1239 4.5005
R86055 VDD.n1304 VDD.n1239 4.5005
R86056 VDD.n1385 VDD.n1239 4.5005
R86057 VDD.n1303 VDD.n1239 4.5005
R86058 VDD.n1386 VDD.n1239 4.5005
R86059 VDD.n1301 VDD.n1239 4.5005
R86060 VDD.n1387 VDD.n1239 4.5005
R86061 VDD.n1300 VDD.n1239 4.5005
R86062 VDD.n1388 VDD.n1239 4.5005
R86063 VDD.n1298 VDD.n1239 4.5005
R86064 VDD.n1389 VDD.n1239 4.5005
R86065 VDD.n1297 VDD.n1239 4.5005
R86066 VDD.n1390 VDD.n1239 4.5005
R86067 VDD.n1295 VDD.n1239 4.5005
R86068 VDD.n1391 VDD.n1239 4.5005
R86069 VDD.n1294 VDD.n1239 4.5005
R86070 VDD.n1392 VDD.n1239 4.5005
R86071 VDD.n1292 VDD.n1239 4.5005
R86072 VDD.n1393 VDD.n1239 4.5005
R86073 VDD.n1291 VDD.n1239 4.5005
R86074 VDD.n1394 VDD.n1239 4.5005
R86075 VDD.n1289 VDD.n1239 4.5005
R86076 VDD.n1395 VDD.n1239 4.5005
R86077 VDD.n1288 VDD.n1239 4.5005
R86078 VDD.n1396 VDD.n1239 4.5005
R86079 VDD.n1286 VDD.n1239 4.5005
R86080 VDD.n1397 VDD.n1239 4.5005
R86081 VDD.n1285 VDD.n1239 4.5005
R86082 VDD.n1398 VDD.n1239 4.5005
R86083 VDD.n1283 VDD.n1239 4.5005
R86084 VDD.n1399 VDD.n1239 4.5005
R86085 VDD.n1282 VDD.n1239 4.5005
R86086 VDD.n1400 VDD.n1239 4.5005
R86087 VDD.n1280 VDD.n1239 4.5005
R86088 VDD.n1401 VDD.n1239 4.5005
R86089 VDD.n1279 VDD.n1239 4.5005
R86090 VDD.n1402 VDD.n1239 4.5005
R86091 VDD.n1277 VDD.n1239 4.5005
R86092 VDD.n1403 VDD.n1239 4.5005
R86093 VDD.n1276 VDD.n1239 4.5005
R86094 VDD.n1404 VDD.n1239 4.5005
R86095 VDD.n1274 VDD.n1239 4.5005
R86096 VDD.n1405 VDD.n1239 4.5005
R86097 VDD.n1273 VDD.n1239 4.5005
R86098 VDD.n1406 VDD.n1239 4.5005
R86099 VDD.n1271 VDD.n1239 4.5005
R86100 VDD.n1407 VDD.n1239 4.5005
R86101 VDD.n1270 VDD.n1239 4.5005
R86102 VDD.n1408 VDD.n1239 4.5005
R86103 VDD.n1268 VDD.n1239 4.5005
R86104 VDD.n1409 VDD.n1239 4.5005
R86105 VDD.n1267 VDD.n1239 4.5005
R86106 VDD.n1410 VDD.n1239 4.5005
R86107 VDD.n1265 VDD.n1239 4.5005
R86108 VDD.n1411 VDD.n1239 4.5005
R86109 VDD.n1264 VDD.n1239 4.5005
R86110 VDD.n1412 VDD.n1239 4.5005
R86111 VDD.n1262 VDD.n1239 4.5005
R86112 VDD.n1413 VDD.n1239 4.5005
R86113 VDD.n1261 VDD.n1239 4.5005
R86114 VDD.n1414 VDD.n1239 4.5005
R86115 VDD.n1415 VDD.n1239 4.5005
R86116 VDD.n1674 VDD.n1239 4.5005
R86117 VDD.n1676 VDD.n1150 4.5005
R86118 VDD.n1341 VDD.n1150 4.5005
R86119 VDD.n1342 VDD.n1150 4.5005
R86120 VDD.n1340 VDD.n1150 4.5005
R86121 VDD.n1344 VDD.n1150 4.5005
R86122 VDD.n1339 VDD.n1150 4.5005
R86123 VDD.n1345 VDD.n1150 4.5005
R86124 VDD.n1338 VDD.n1150 4.5005
R86125 VDD.n1347 VDD.n1150 4.5005
R86126 VDD.n1337 VDD.n1150 4.5005
R86127 VDD.n1348 VDD.n1150 4.5005
R86128 VDD.n1336 VDD.n1150 4.5005
R86129 VDD.n1350 VDD.n1150 4.5005
R86130 VDD.n1335 VDD.n1150 4.5005
R86131 VDD.n1351 VDD.n1150 4.5005
R86132 VDD.n1334 VDD.n1150 4.5005
R86133 VDD.n1353 VDD.n1150 4.5005
R86134 VDD.n1333 VDD.n1150 4.5005
R86135 VDD.n1354 VDD.n1150 4.5005
R86136 VDD.n1332 VDD.n1150 4.5005
R86137 VDD.n1356 VDD.n1150 4.5005
R86138 VDD.n1331 VDD.n1150 4.5005
R86139 VDD.n1357 VDD.n1150 4.5005
R86140 VDD.n1330 VDD.n1150 4.5005
R86141 VDD.n1359 VDD.n1150 4.5005
R86142 VDD.n1329 VDD.n1150 4.5005
R86143 VDD.n1360 VDD.n1150 4.5005
R86144 VDD.n1328 VDD.n1150 4.5005
R86145 VDD.n1362 VDD.n1150 4.5005
R86146 VDD.n1327 VDD.n1150 4.5005
R86147 VDD.n1363 VDD.n1150 4.5005
R86148 VDD.n1326 VDD.n1150 4.5005
R86149 VDD.n1365 VDD.n1150 4.5005
R86150 VDD.n1325 VDD.n1150 4.5005
R86151 VDD.n1366 VDD.n1150 4.5005
R86152 VDD.n1324 VDD.n1150 4.5005
R86153 VDD.n1368 VDD.n1150 4.5005
R86154 VDD.n1323 VDD.n1150 4.5005
R86155 VDD.n1369 VDD.n1150 4.5005
R86156 VDD.n1322 VDD.n1150 4.5005
R86157 VDD.n1371 VDD.n1150 4.5005
R86158 VDD.n1321 VDD.n1150 4.5005
R86159 VDD.n1372 VDD.n1150 4.5005
R86160 VDD.n1320 VDD.n1150 4.5005
R86161 VDD.n1374 VDD.n1150 4.5005
R86162 VDD.n1319 VDD.n1150 4.5005
R86163 VDD.n1375 VDD.n1150 4.5005
R86164 VDD.n1318 VDD.n1150 4.5005
R86165 VDD.n1376 VDD.n1150 4.5005
R86166 VDD.n1316 VDD.n1150 4.5005
R86167 VDD.n1377 VDD.n1150 4.5005
R86168 VDD.n1315 VDD.n1150 4.5005
R86169 VDD.n1378 VDD.n1150 4.5005
R86170 VDD.n1313 VDD.n1150 4.5005
R86171 VDD.n1379 VDD.n1150 4.5005
R86172 VDD.n1312 VDD.n1150 4.5005
R86173 VDD.n1380 VDD.n1150 4.5005
R86174 VDD.n1310 VDD.n1150 4.5005
R86175 VDD.n1381 VDD.n1150 4.5005
R86176 VDD.n1309 VDD.n1150 4.5005
R86177 VDD.n1382 VDD.n1150 4.5005
R86178 VDD.n1307 VDD.n1150 4.5005
R86179 VDD.n1383 VDD.n1150 4.5005
R86180 VDD.n1306 VDD.n1150 4.5005
R86181 VDD.n1384 VDD.n1150 4.5005
R86182 VDD.n1304 VDD.n1150 4.5005
R86183 VDD.n1385 VDD.n1150 4.5005
R86184 VDD.n1303 VDD.n1150 4.5005
R86185 VDD.n1386 VDD.n1150 4.5005
R86186 VDD.n1301 VDD.n1150 4.5005
R86187 VDD.n1387 VDD.n1150 4.5005
R86188 VDD.n1300 VDD.n1150 4.5005
R86189 VDD.n1388 VDD.n1150 4.5005
R86190 VDD.n1298 VDD.n1150 4.5005
R86191 VDD.n1389 VDD.n1150 4.5005
R86192 VDD.n1297 VDD.n1150 4.5005
R86193 VDD.n1390 VDD.n1150 4.5005
R86194 VDD.n1295 VDD.n1150 4.5005
R86195 VDD.n1391 VDD.n1150 4.5005
R86196 VDD.n1294 VDD.n1150 4.5005
R86197 VDD.n1392 VDD.n1150 4.5005
R86198 VDD.n1292 VDD.n1150 4.5005
R86199 VDD.n1393 VDD.n1150 4.5005
R86200 VDD.n1291 VDD.n1150 4.5005
R86201 VDD.n1394 VDD.n1150 4.5005
R86202 VDD.n1289 VDD.n1150 4.5005
R86203 VDD.n1395 VDD.n1150 4.5005
R86204 VDD.n1288 VDD.n1150 4.5005
R86205 VDD.n1396 VDD.n1150 4.5005
R86206 VDD.n1286 VDD.n1150 4.5005
R86207 VDD.n1397 VDD.n1150 4.5005
R86208 VDD.n1285 VDD.n1150 4.5005
R86209 VDD.n1398 VDD.n1150 4.5005
R86210 VDD.n1283 VDD.n1150 4.5005
R86211 VDD.n1399 VDD.n1150 4.5005
R86212 VDD.n1282 VDD.n1150 4.5005
R86213 VDD.n1400 VDD.n1150 4.5005
R86214 VDD.n1280 VDD.n1150 4.5005
R86215 VDD.n1401 VDD.n1150 4.5005
R86216 VDD.n1279 VDD.n1150 4.5005
R86217 VDD.n1402 VDD.n1150 4.5005
R86218 VDD.n1277 VDD.n1150 4.5005
R86219 VDD.n1403 VDD.n1150 4.5005
R86220 VDD.n1276 VDD.n1150 4.5005
R86221 VDD.n1404 VDD.n1150 4.5005
R86222 VDD.n1274 VDD.n1150 4.5005
R86223 VDD.n1405 VDD.n1150 4.5005
R86224 VDD.n1273 VDD.n1150 4.5005
R86225 VDD.n1406 VDD.n1150 4.5005
R86226 VDD.n1271 VDD.n1150 4.5005
R86227 VDD.n1407 VDD.n1150 4.5005
R86228 VDD.n1270 VDD.n1150 4.5005
R86229 VDD.n1408 VDD.n1150 4.5005
R86230 VDD.n1268 VDD.n1150 4.5005
R86231 VDD.n1409 VDD.n1150 4.5005
R86232 VDD.n1267 VDD.n1150 4.5005
R86233 VDD.n1410 VDD.n1150 4.5005
R86234 VDD.n1265 VDD.n1150 4.5005
R86235 VDD.n1411 VDD.n1150 4.5005
R86236 VDD.n1264 VDD.n1150 4.5005
R86237 VDD.n1412 VDD.n1150 4.5005
R86238 VDD.n1262 VDD.n1150 4.5005
R86239 VDD.n1413 VDD.n1150 4.5005
R86240 VDD.n1261 VDD.n1150 4.5005
R86241 VDD.n1414 VDD.n1150 4.5005
R86242 VDD.n1415 VDD.n1150 4.5005
R86243 VDD.n1674 VDD.n1150 4.5005
R86244 VDD.n1676 VDD.n1240 4.5005
R86245 VDD.n1341 VDD.n1240 4.5005
R86246 VDD.n1342 VDD.n1240 4.5005
R86247 VDD.n1340 VDD.n1240 4.5005
R86248 VDD.n1344 VDD.n1240 4.5005
R86249 VDD.n1339 VDD.n1240 4.5005
R86250 VDD.n1345 VDD.n1240 4.5005
R86251 VDD.n1338 VDD.n1240 4.5005
R86252 VDD.n1347 VDD.n1240 4.5005
R86253 VDD.n1337 VDD.n1240 4.5005
R86254 VDD.n1348 VDD.n1240 4.5005
R86255 VDD.n1336 VDD.n1240 4.5005
R86256 VDD.n1350 VDD.n1240 4.5005
R86257 VDD.n1335 VDD.n1240 4.5005
R86258 VDD.n1351 VDD.n1240 4.5005
R86259 VDD.n1334 VDD.n1240 4.5005
R86260 VDD.n1353 VDD.n1240 4.5005
R86261 VDD.n1333 VDD.n1240 4.5005
R86262 VDD.n1354 VDD.n1240 4.5005
R86263 VDD.n1332 VDD.n1240 4.5005
R86264 VDD.n1356 VDD.n1240 4.5005
R86265 VDD.n1331 VDD.n1240 4.5005
R86266 VDD.n1357 VDD.n1240 4.5005
R86267 VDD.n1330 VDD.n1240 4.5005
R86268 VDD.n1359 VDD.n1240 4.5005
R86269 VDD.n1329 VDD.n1240 4.5005
R86270 VDD.n1360 VDD.n1240 4.5005
R86271 VDD.n1328 VDD.n1240 4.5005
R86272 VDD.n1362 VDD.n1240 4.5005
R86273 VDD.n1327 VDD.n1240 4.5005
R86274 VDD.n1363 VDD.n1240 4.5005
R86275 VDD.n1326 VDD.n1240 4.5005
R86276 VDD.n1365 VDD.n1240 4.5005
R86277 VDD.n1325 VDD.n1240 4.5005
R86278 VDD.n1366 VDD.n1240 4.5005
R86279 VDD.n1324 VDD.n1240 4.5005
R86280 VDD.n1368 VDD.n1240 4.5005
R86281 VDD.n1323 VDD.n1240 4.5005
R86282 VDD.n1369 VDD.n1240 4.5005
R86283 VDD.n1322 VDD.n1240 4.5005
R86284 VDD.n1371 VDD.n1240 4.5005
R86285 VDD.n1321 VDD.n1240 4.5005
R86286 VDD.n1372 VDD.n1240 4.5005
R86287 VDD.n1320 VDD.n1240 4.5005
R86288 VDD.n1374 VDD.n1240 4.5005
R86289 VDD.n1319 VDD.n1240 4.5005
R86290 VDD.n1375 VDD.n1240 4.5005
R86291 VDD.n1318 VDD.n1240 4.5005
R86292 VDD.n1376 VDD.n1240 4.5005
R86293 VDD.n1316 VDD.n1240 4.5005
R86294 VDD.n1377 VDD.n1240 4.5005
R86295 VDD.n1315 VDD.n1240 4.5005
R86296 VDD.n1378 VDD.n1240 4.5005
R86297 VDD.n1313 VDD.n1240 4.5005
R86298 VDD.n1379 VDD.n1240 4.5005
R86299 VDD.n1312 VDD.n1240 4.5005
R86300 VDD.n1380 VDD.n1240 4.5005
R86301 VDD.n1310 VDD.n1240 4.5005
R86302 VDD.n1381 VDD.n1240 4.5005
R86303 VDD.n1309 VDD.n1240 4.5005
R86304 VDD.n1382 VDD.n1240 4.5005
R86305 VDD.n1307 VDD.n1240 4.5005
R86306 VDD.n1383 VDD.n1240 4.5005
R86307 VDD.n1306 VDD.n1240 4.5005
R86308 VDD.n1384 VDD.n1240 4.5005
R86309 VDD.n1304 VDD.n1240 4.5005
R86310 VDD.n1385 VDD.n1240 4.5005
R86311 VDD.n1303 VDD.n1240 4.5005
R86312 VDD.n1386 VDD.n1240 4.5005
R86313 VDD.n1301 VDD.n1240 4.5005
R86314 VDD.n1387 VDD.n1240 4.5005
R86315 VDD.n1300 VDD.n1240 4.5005
R86316 VDD.n1388 VDD.n1240 4.5005
R86317 VDD.n1298 VDD.n1240 4.5005
R86318 VDD.n1389 VDD.n1240 4.5005
R86319 VDD.n1297 VDD.n1240 4.5005
R86320 VDD.n1390 VDD.n1240 4.5005
R86321 VDD.n1295 VDD.n1240 4.5005
R86322 VDD.n1391 VDD.n1240 4.5005
R86323 VDD.n1294 VDD.n1240 4.5005
R86324 VDD.n1392 VDD.n1240 4.5005
R86325 VDD.n1292 VDD.n1240 4.5005
R86326 VDD.n1393 VDD.n1240 4.5005
R86327 VDD.n1291 VDD.n1240 4.5005
R86328 VDD.n1394 VDD.n1240 4.5005
R86329 VDD.n1289 VDD.n1240 4.5005
R86330 VDD.n1395 VDD.n1240 4.5005
R86331 VDD.n1288 VDD.n1240 4.5005
R86332 VDD.n1396 VDD.n1240 4.5005
R86333 VDD.n1286 VDD.n1240 4.5005
R86334 VDD.n1397 VDD.n1240 4.5005
R86335 VDD.n1285 VDD.n1240 4.5005
R86336 VDD.n1398 VDD.n1240 4.5005
R86337 VDD.n1283 VDD.n1240 4.5005
R86338 VDD.n1399 VDD.n1240 4.5005
R86339 VDD.n1282 VDD.n1240 4.5005
R86340 VDD.n1400 VDD.n1240 4.5005
R86341 VDD.n1280 VDD.n1240 4.5005
R86342 VDD.n1401 VDD.n1240 4.5005
R86343 VDD.n1279 VDD.n1240 4.5005
R86344 VDD.n1402 VDD.n1240 4.5005
R86345 VDD.n1277 VDD.n1240 4.5005
R86346 VDD.n1403 VDD.n1240 4.5005
R86347 VDD.n1276 VDD.n1240 4.5005
R86348 VDD.n1404 VDD.n1240 4.5005
R86349 VDD.n1274 VDD.n1240 4.5005
R86350 VDD.n1405 VDD.n1240 4.5005
R86351 VDD.n1273 VDD.n1240 4.5005
R86352 VDD.n1406 VDD.n1240 4.5005
R86353 VDD.n1271 VDD.n1240 4.5005
R86354 VDD.n1407 VDD.n1240 4.5005
R86355 VDD.n1270 VDD.n1240 4.5005
R86356 VDD.n1408 VDD.n1240 4.5005
R86357 VDD.n1268 VDD.n1240 4.5005
R86358 VDD.n1409 VDD.n1240 4.5005
R86359 VDD.n1267 VDD.n1240 4.5005
R86360 VDD.n1410 VDD.n1240 4.5005
R86361 VDD.n1265 VDD.n1240 4.5005
R86362 VDD.n1411 VDD.n1240 4.5005
R86363 VDD.n1264 VDD.n1240 4.5005
R86364 VDD.n1412 VDD.n1240 4.5005
R86365 VDD.n1262 VDD.n1240 4.5005
R86366 VDD.n1413 VDD.n1240 4.5005
R86367 VDD.n1261 VDD.n1240 4.5005
R86368 VDD.n1414 VDD.n1240 4.5005
R86369 VDD.n1415 VDD.n1240 4.5005
R86370 VDD.n1674 VDD.n1240 4.5005
R86371 VDD.n1676 VDD.n1149 4.5005
R86372 VDD.n1341 VDD.n1149 4.5005
R86373 VDD.n1342 VDD.n1149 4.5005
R86374 VDD.n1340 VDD.n1149 4.5005
R86375 VDD.n1344 VDD.n1149 4.5005
R86376 VDD.n1339 VDD.n1149 4.5005
R86377 VDD.n1345 VDD.n1149 4.5005
R86378 VDD.n1338 VDD.n1149 4.5005
R86379 VDD.n1347 VDD.n1149 4.5005
R86380 VDD.n1337 VDD.n1149 4.5005
R86381 VDD.n1348 VDD.n1149 4.5005
R86382 VDD.n1336 VDD.n1149 4.5005
R86383 VDD.n1350 VDD.n1149 4.5005
R86384 VDD.n1335 VDD.n1149 4.5005
R86385 VDD.n1351 VDD.n1149 4.5005
R86386 VDD.n1334 VDD.n1149 4.5005
R86387 VDD.n1353 VDD.n1149 4.5005
R86388 VDD.n1333 VDD.n1149 4.5005
R86389 VDD.n1354 VDD.n1149 4.5005
R86390 VDD.n1332 VDD.n1149 4.5005
R86391 VDD.n1356 VDD.n1149 4.5005
R86392 VDD.n1331 VDD.n1149 4.5005
R86393 VDD.n1357 VDD.n1149 4.5005
R86394 VDD.n1330 VDD.n1149 4.5005
R86395 VDD.n1359 VDD.n1149 4.5005
R86396 VDD.n1329 VDD.n1149 4.5005
R86397 VDD.n1360 VDD.n1149 4.5005
R86398 VDD.n1328 VDD.n1149 4.5005
R86399 VDD.n1362 VDD.n1149 4.5005
R86400 VDD.n1327 VDD.n1149 4.5005
R86401 VDD.n1363 VDD.n1149 4.5005
R86402 VDD.n1326 VDD.n1149 4.5005
R86403 VDD.n1365 VDD.n1149 4.5005
R86404 VDD.n1325 VDD.n1149 4.5005
R86405 VDD.n1366 VDD.n1149 4.5005
R86406 VDD.n1324 VDD.n1149 4.5005
R86407 VDD.n1368 VDD.n1149 4.5005
R86408 VDD.n1323 VDD.n1149 4.5005
R86409 VDD.n1369 VDD.n1149 4.5005
R86410 VDD.n1322 VDD.n1149 4.5005
R86411 VDD.n1371 VDD.n1149 4.5005
R86412 VDD.n1321 VDD.n1149 4.5005
R86413 VDD.n1372 VDD.n1149 4.5005
R86414 VDD.n1320 VDD.n1149 4.5005
R86415 VDD.n1374 VDD.n1149 4.5005
R86416 VDD.n1319 VDD.n1149 4.5005
R86417 VDD.n1375 VDD.n1149 4.5005
R86418 VDD.n1318 VDD.n1149 4.5005
R86419 VDD.n1376 VDD.n1149 4.5005
R86420 VDD.n1316 VDD.n1149 4.5005
R86421 VDD.n1377 VDD.n1149 4.5005
R86422 VDD.n1315 VDD.n1149 4.5005
R86423 VDD.n1378 VDD.n1149 4.5005
R86424 VDD.n1313 VDD.n1149 4.5005
R86425 VDD.n1379 VDD.n1149 4.5005
R86426 VDD.n1312 VDD.n1149 4.5005
R86427 VDD.n1380 VDD.n1149 4.5005
R86428 VDD.n1310 VDD.n1149 4.5005
R86429 VDD.n1381 VDD.n1149 4.5005
R86430 VDD.n1309 VDD.n1149 4.5005
R86431 VDD.n1382 VDD.n1149 4.5005
R86432 VDD.n1307 VDD.n1149 4.5005
R86433 VDD.n1383 VDD.n1149 4.5005
R86434 VDD.n1306 VDD.n1149 4.5005
R86435 VDD.n1384 VDD.n1149 4.5005
R86436 VDD.n1304 VDD.n1149 4.5005
R86437 VDD.n1385 VDD.n1149 4.5005
R86438 VDD.n1303 VDD.n1149 4.5005
R86439 VDD.n1386 VDD.n1149 4.5005
R86440 VDD.n1301 VDD.n1149 4.5005
R86441 VDD.n1387 VDD.n1149 4.5005
R86442 VDD.n1300 VDD.n1149 4.5005
R86443 VDD.n1388 VDD.n1149 4.5005
R86444 VDD.n1298 VDD.n1149 4.5005
R86445 VDD.n1389 VDD.n1149 4.5005
R86446 VDD.n1297 VDD.n1149 4.5005
R86447 VDD.n1390 VDD.n1149 4.5005
R86448 VDD.n1295 VDD.n1149 4.5005
R86449 VDD.n1391 VDD.n1149 4.5005
R86450 VDD.n1294 VDD.n1149 4.5005
R86451 VDD.n1392 VDD.n1149 4.5005
R86452 VDD.n1292 VDD.n1149 4.5005
R86453 VDD.n1393 VDD.n1149 4.5005
R86454 VDD.n1291 VDD.n1149 4.5005
R86455 VDD.n1394 VDD.n1149 4.5005
R86456 VDD.n1289 VDD.n1149 4.5005
R86457 VDD.n1395 VDD.n1149 4.5005
R86458 VDD.n1288 VDD.n1149 4.5005
R86459 VDD.n1396 VDD.n1149 4.5005
R86460 VDD.n1286 VDD.n1149 4.5005
R86461 VDD.n1397 VDD.n1149 4.5005
R86462 VDD.n1285 VDD.n1149 4.5005
R86463 VDD.n1398 VDD.n1149 4.5005
R86464 VDD.n1283 VDD.n1149 4.5005
R86465 VDD.n1399 VDD.n1149 4.5005
R86466 VDD.n1282 VDD.n1149 4.5005
R86467 VDD.n1400 VDD.n1149 4.5005
R86468 VDD.n1280 VDD.n1149 4.5005
R86469 VDD.n1401 VDD.n1149 4.5005
R86470 VDD.n1279 VDD.n1149 4.5005
R86471 VDD.n1402 VDD.n1149 4.5005
R86472 VDD.n1277 VDD.n1149 4.5005
R86473 VDD.n1403 VDD.n1149 4.5005
R86474 VDD.n1276 VDD.n1149 4.5005
R86475 VDD.n1404 VDD.n1149 4.5005
R86476 VDD.n1274 VDD.n1149 4.5005
R86477 VDD.n1405 VDD.n1149 4.5005
R86478 VDD.n1273 VDD.n1149 4.5005
R86479 VDD.n1406 VDD.n1149 4.5005
R86480 VDD.n1271 VDD.n1149 4.5005
R86481 VDD.n1407 VDD.n1149 4.5005
R86482 VDD.n1270 VDD.n1149 4.5005
R86483 VDD.n1408 VDD.n1149 4.5005
R86484 VDD.n1268 VDD.n1149 4.5005
R86485 VDD.n1409 VDD.n1149 4.5005
R86486 VDD.n1267 VDD.n1149 4.5005
R86487 VDD.n1410 VDD.n1149 4.5005
R86488 VDD.n1265 VDD.n1149 4.5005
R86489 VDD.n1411 VDD.n1149 4.5005
R86490 VDD.n1264 VDD.n1149 4.5005
R86491 VDD.n1412 VDD.n1149 4.5005
R86492 VDD.n1262 VDD.n1149 4.5005
R86493 VDD.n1413 VDD.n1149 4.5005
R86494 VDD.n1261 VDD.n1149 4.5005
R86495 VDD.n1414 VDD.n1149 4.5005
R86496 VDD.n1415 VDD.n1149 4.5005
R86497 VDD.n1674 VDD.n1149 4.5005
R86498 VDD.n1676 VDD.n1241 4.5005
R86499 VDD.n1341 VDD.n1241 4.5005
R86500 VDD.n1342 VDD.n1241 4.5005
R86501 VDD.n1340 VDD.n1241 4.5005
R86502 VDD.n1344 VDD.n1241 4.5005
R86503 VDD.n1339 VDD.n1241 4.5005
R86504 VDD.n1345 VDD.n1241 4.5005
R86505 VDD.n1338 VDD.n1241 4.5005
R86506 VDD.n1347 VDD.n1241 4.5005
R86507 VDD.n1337 VDD.n1241 4.5005
R86508 VDD.n1348 VDD.n1241 4.5005
R86509 VDD.n1336 VDD.n1241 4.5005
R86510 VDD.n1350 VDD.n1241 4.5005
R86511 VDD.n1335 VDD.n1241 4.5005
R86512 VDD.n1351 VDD.n1241 4.5005
R86513 VDD.n1334 VDD.n1241 4.5005
R86514 VDD.n1353 VDD.n1241 4.5005
R86515 VDD.n1333 VDD.n1241 4.5005
R86516 VDD.n1354 VDD.n1241 4.5005
R86517 VDD.n1332 VDD.n1241 4.5005
R86518 VDD.n1356 VDD.n1241 4.5005
R86519 VDD.n1331 VDD.n1241 4.5005
R86520 VDD.n1357 VDD.n1241 4.5005
R86521 VDD.n1330 VDD.n1241 4.5005
R86522 VDD.n1359 VDD.n1241 4.5005
R86523 VDD.n1329 VDD.n1241 4.5005
R86524 VDD.n1360 VDD.n1241 4.5005
R86525 VDD.n1328 VDD.n1241 4.5005
R86526 VDD.n1362 VDD.n1241 4.5005
R86527 VDD.n1327 VDD.n1241 4.5005
R86528 VDD.n1363 VDD.n1241 4.5005
R86529 VDD.n1326 VDD.n1241 4.5005
R86530 VDD.n1365 VDD.n1241 4.5005
R86531 VDD.n1325 VDD.n1241 4.5005
R86532 VDD.n1366 VDD.n1241 4.5005
R86533 VDD.n1324 VDD.n1241 4.5005
R86534 VDD.n1368 VDD.n1241 4.5005
R86535 VDD.n1323 VDD.n1241 4.5005
R86536 VDD.n1369 VDD.n1241 4.5005
R86537 VDD.n1322 VDD.n1241 4.5005
R86538 VDD.n1371 VDD.n1241 4.5005
R86539 VDD.n1321 VDD.n1241 4.5005
R86540 VDD.n1372 VDD.n1241 4.5005
R86541 VDD.n1320 VDD.n1241 4.5005
R86542 VDD.n1374 VDD.n1241 4.5005
R86543 VDD.n1319 VDD.n1241 4.5005
R86544 VDD.n1375 VDD.n1241 4.5005
R86545 VDD.n1318 VDD.n1241 4.5005
R86546 VDD.n1376 VDD.n1241 4.5005
R86547 VDD.n1316 VDD.n1241 4.5005
R86548 VDD.n1377 VDD.n1241 4.5005
R86549 VDD.n1315 VDD.n1241 4.5005
R86550 VDD.n1378 VDD.n1241 4.5005
R86551 VDD.n1313 VDD.n1241 4.5005
R86552 VDD.n1379 VDD.n1241 4.5005
R86553 VDD.n1312 VDD.n1241 4.5005
R86554 VDD.n1380 VDD.n1241 4.5005
R86555 VDD.n1310 VDD.n1241 4.5005
R86556 VDD.n1381 VDD.n1241 4.5005
R86557 VDD.n1309 VDD.n1241 4.5005
R86558 VDD.n1382 VDD.n1241 4.5005
R86559 VDD.n1307 VDD.n1241 4.5005
R86560 VDD.n1383 VDD.n1241 4.5005
R86561 VDD.n1306 VDD.n1241 4.5005
R86562 VDD.n1384 VDD.n1241 4.5005
R86563 VDD.n1304 VDD.n1241 4.5005
R86564 VDD.n1385 VDD.n1241 4.5005
R86565 VDD.n1303 VDD.n1241 4.5005
R86566 VDD.n1386 VDD.n1241 4.5005
R86567 VDD.n1301 VDD.n1241 4.5005
R86568 VDD.n1387 VDD.n1241 4.5005
R86569 VDD.n1300 VDD.n1241 4.5005
R86570 VDD.n1388 VDD.n1241 4.5005
R86571 VDD.n1298 VDD.n1241 4.5005
R86572 VDD.n1389 VDD.n1241 4.5005
R86573 VDD.n1297 VDD.n1241 4.5005
R86574 VDD.n1390 VDD.n1241 4.5005
R86575 VDD.n1295 VDD.n1241 4.5005
R86576 VDD.n1391 VDD.n1241 4.5005
R86577 VDD.n1294 VDD.n1241 4.5005
R86578 VDD.n1392 VDD.n1241 4.5005
R86579 VDD.n1292 VDD.n1241 4.5005
R86580 VDD.n1393 VDD.n1241 4.5005
R86581 VDD.n1291 VDD.n1241 4.5005
R86582 VDD.n1394 VDD.n1241 4.5005
R86583 VDD.n1289 VDD.n1241 4.5005
R86584 VDD.n1395 VDD.n1241 4.5005
R86585 VDD.n1288 VDD.n1241 4.5005
R86586 VDD.n1396 VDD.n1241 4.5005
R86587 VDD.n1286 VDD.n1241 4.5005
R86588 VDD.n1397 VDD.n1241 4.5005
R86589 VDD.n1285 VDD.n1241 4.5005
R86590 VDD.n1398 VDD.n1241 4.5005
R86591 VDD.n1283 VDD.n1241 4.5005
R86592 VDD.n1399 VDD.n1241 4.5005
R86593 VDD.n1282 VDD.n1241 4.5005
R86594 VDD.n1400 VDD.n1241 4.5005
R86595 VDD.n1280 VDD.n1241 4.5005
R86596 VDD.n1401 VDD.n1241 4.5005
R86597 VDD.n1279 VDD.n1241 4.5005
R86598 VDD.n1402 VDD.n1241 4.5005
R86599 VDD.n1277 VDD.n1241 4.5005
R86600 VDD.n1403 VDD.n1241 4.5005
R86601 VDD.n1276 VDD.n1241 4.5005
R86602 VDD.n1404 VDD.n1241 4.5005
R86603 VDD.n1274 VDD.n1241 4.5005
R86604 VDD.n1405 VDD.n1241 4.5005
R86605 VDD.n1273 VDD.n1241 4.5005
R86606 VDD.n1406 VDD.n1241 4.5005
R86607 VDD.n1271 VDD.n1241 4.5005
R86608 VDD.n1407 VDD.n1241 4.5005
R86609 VDD.n1270 VDD.n1241 4.5005
R86610 VDD.n1408 VDD.n1241 4.5005
R86611 VDD.n1268 VDD.n1241 4.5005
R86612 VDD.n1409 VDD.n1241 4.5005
R86613 VDD.n1267 VDD.n1241 4.5005
R86614 VDD.n1410 VDD.n1241 4.5005
R86615 VDD.n1265 VDD.n1241 4.5005
R86616 VDD.n1411 VDD.n1241 4.5005
R86617 VDD.n1264 VDD.n1241 4.5005
R86618 VDD.n1412 VDD.n1241 4.5005
R86619 VDD.n1262 VDD.n1241 4.5005
R86620 VDD.n1413 VDD.n1241 4.5005
R86621 VDD.n1261 VDD.n1241 4.5005
R86622 VDD.n1414 VDD.n1241 4.5005
R86623 VDD.n1415 VDD.n1241 4.5005
R86624 VDD.n1674 VDD.n1241 4.5005
R86625 VDD.n1676 VDD.n1148 4.5005
R86626 VDD.n1341 VDD.n1148 4.5005
R86627 VDD.n1342 VDD.n1148 4.5005
R86628 VDD.n1340 VDD.n1148 4.5005
R86629 VDD.n1344 VDD.n1148 4.5005
R86630 VDD.n1339 VDD.n1148 4.5005
R86631 VDD.n1345 VDD.n1148 4.5005
R86632 VDD.n1338 VDD.n1148 4.5005
R86633 VDD.n1347 VDD.n1148 4.5005
R86634 VDD.n1337 VDD.n1148 4.5005
R86635 VDD.n1348 VDD.n1148 4.5005
R86636 VDD.n1336 VDD.n1148 4.5005
R86637 VDD.n1350 VDD.n1148 4.5005
R86638 VDD.n1335 VDD.n1148 4.5005
R86639 VDD.n1351 VDD.n1148 4.5005
R86640 VDD.n1334 VDD.n1148 4.5005
R86641 VDD.n1353 VDD.n1148 4.5005
R86642 VDD.n1333 VDD.n1148 4.5005
R86643 VDD.n1354 VDD.n1148 4.5005
R86644 VDD.n1332 VDD.n1148 4.5005
R86645 VDD.n1356 VDD.n1148 4.5005
R86646 VDD.n1331 VDD.n1148 4.5005
R86647 VDD.n1357 VDD.n1148 4.5005
R86648 VDD.n1330 VDD.n1148 4.5005
R86649 VDD.n1359 VDD.n1148 4.5005
R86650 VDD.n1329 VDD.n1148 4.5005
R86651 VDD.n1360 VDD.n1148 4.5005
R86652 VDD.n1328 VDD.n1148 4.5005
R86653 VDD.n1362 VDD.n1148 4.5005
R86654 VDD.n1327 VDD.n1148 4.5005
R86655 VDD.n1363 VDD.n1148 4.5005
R86656 VDD.n1326 VDD.n1148 4.5005
R86657 VDD.n1365 VDD.n1148 4.5005
R86658 VDD.n1325 VDD.n1148 4.5005
R86659 VDD.n1366 VDD.n1148 4.5005
R86660 VDD.n1324 VDD.n1148 4.5005
R86661 VDD.n1368 VDD.n1148 4.5005
R86662 VDD.n1323 VDD.n1148 4.5005
R86663 VDD.n1369 VDD.n1148 4.5005
R86664 VDD.n1322 VDD.n1148 4.5005
R86665 VDD.n1371 VDD.n1148 4.5005
R86666 VDD.n1321 VDD.n1148 4.5005
R86667 VDD.n1372 VDD.n1148 4.5005
R86668 VDD.n1320 VDD.n1148 4.5005
R86669 VDD.n1374 VDD.n1148 4.5005
R86670 VDD.n1319 VDD.n1148 4.5005
R86671 VDD.n1375 VDD.n1148 4.5005
R86672 VDD.n1318 VDD.n1148 4.5005
R86673 VDD.n1376 VDD.n1148 4.5005
R86674 VDD.n1316 VDD.n1148 4.5005
R86675 VDD.n1377 VDD.n1148 4.5005
R86676 VDD.n1315 VDD.n1148 4.5005
R86677 VDD.n1378 VDD.n1148 4.5005
R86678 VDD.n1313 VDD.n1148 4.5005
R86679 VDD.n1379 VDD.n1148 4.5005
R86680 VDD.n1312 VDD.n1148 4.5005
R86681 VDD.n1380 VDD.n1148 4.5005
R86682 VDD.n1310 VDD.n1148 4.5005
R86683 VDD.n1381 VDD.n1148 4.5005
R86684 VDD.n1309 VDD.n1148 4.5005
R86685 VDD.n1382 VDD.n1148 4.5005
R86686 VDD.n1307 VDD.n1148 4.5005
R86687 VDD.n1383 VDD.n1148 4.5005
R86688 VDD.n1306 VDD.n1148 4.5005
R86689 VDD.n1384 VDD.n1148 4.5005
R86690 VDD.n1304 VDD.n1148 4.5005
R86691 VDD.n1385 VDD.n1148 4.5005
R86692 VDD.n1303 VDD.n1148 4.5005
R86693 VDD.n1386 VDD.n1148 4.5005
R86694 VDD.n1301 VDD.n1148 4.5005
R86695 VDD.n1387 VDD.n1148 4.5005
R86696 VDD.n1300 VDD.n1148 4.5005
R86697 VDD.n1388 VDD.n1148 4.5005
R86698 VDD.n1298 VDD.n1148 4.5005
R86699 VDD.n1389 VDD.n1148 4.5005
R86700 VDD.n1297 VDD.n1148 4.5005
R86701 VDD.n1390 VDD.n1148 4.5005
R86702 VDD.n1295 VDD.n1148 4.5005
R86703 VDD.n1391 VDD.n1148 4.5005
R86704 VDD.n1294 VDD.n1148 4.5005
R86705 VDD.n1392 VDD.n1148 4.5005
R86706 VDD.n1292 VDD.n1148 4.5005
R86707 VDD.n1393 VDD.n1148 4.5005
R86708 VDD.n1291 VDD.n1148 4.5005
R86709 VDD.n1394 VDD.n1148 4.5005
R86710 VDD.n1289 VDD.n1148 4.5005
R86711 VDD.n1395 VDD.n1148 4.5005
R86712 VDD.n1288 VDD.n1148 4.5005
R86713 VDD.n1396 VDD.n1148 4.5005
R86714 VDD.n1286 VDD.n1148 4.5005
R86715 VDD.n1397 VDD.n1148 4.5005
R86716 VDD.n1285 VDD.n1148 4.5005
R86717 VDD.n1398 VDD.n1148 4.5005
R86718 VDD.n1283 VDD.n1148 4.5005
R86719 VDD.n1399 VDD.n1148 4.5005
R86720 VDD.n1282 VDD.n1148 4.5005
R86721 VDD.n1400 VDD.n1148 4.5005
R86722 VDD.n1280 VDD.n1148 4.5005
R86723 VDD.n1401 VDD.n1148 4.5005
R86724 VDD.n1279 VDD.n1148 4.5005
R86725 VDD.n1402 VDD.n1148 4.5005
R86726 VDD.n1277 VDD.n1148 4.5005
R86727 VDD.n1403 VDD.n1148 4.5005
R86728 VDD.n1276 VDD.n1148 4.5005
R86729 VDD.n1404 VDD.n1148 4.5005
R86730 VDD.n1274 VDD.n1148 4.5005
R86731 VDD.n1405 VDD.n1148 4.5005
R86732 VDD.n1273 VDD.n1148 4.5005
R86733 VDD.n1406 VDD.n1148 4.5005
R86734 VDD.n1271 VDD.n1148 4.5005
R86735 VDD.n1407 VDD.n1148 4.5005
R86736 VDD.n1270 VDD.n1148 4.5005
R86737 VDD.n1408 VDD.n1148 4.5005
R86738 VDD.n1268 VDD.n1148 4.5005
R86739 VDD.n1409 VDD.n1148 4.5005
R86740 VDD.n1267 VDD.n1148 4.5005
R86741 VDD.n1410 VDD.n1148 4.5005
R86742 VDD.n1265 VDD.n1148 4.5005
R86743 VDD.n1411 VDD.n1148 4.5005
R86744 VDD.n1264 VDD.n1148 4.5005
R86745 VDD.n1412 VDD.n1148 4.5005
R86746 VDD.n1262 VDD.n1148 4.5005
R86747 VDD.n1413 VDD.n1148 4.5005
R86748 VDD.n1261 VDD.n1148 4.5005
R86749 VDD.n1414 VDD.n1148 4.5005
R86750 VDD.n1415 VDD.n1148 4.5005
R86751 VDD.n1674 VDD.n1148 4.5005
R86752 VDD.n1676 VDD.n1242 4.5005
R86753 VDD.n1341 VDD.n1242 4.5005
R86754 VDD.n1342 VDD.n1242 4.5005
R86755 VDD.n1340 VDD.n1242 4.5005
R86756 VDD.n1344 VDD.n1242 4.5005
R86757 VDD.n1339 VDD.n1242 4.5005
R86758 VDD.n1345 VDD.n1242 4.5005
R86759 VDD.n1338 VDD.n1242 4.5005
R86760 VDD.n1347 VDD.n1242 4.5005
R86761 VDD.n1337 VDD.n1242 4.5005
R86762 VDD.n1348 VDD.n1242 4.5005
R86763 VDD.n1336 VDD.n1242 4.5005
R86764 VDD.n1350 VDD.n1242 4.5005
R86765 VDD.n1335 VDD.n1242 4.5005
R86766 VDD.n1351 VDD.n1242 4.5005
R86767 VDD.n1334 VDD.n1242 4.5005
R86768 VDD.n1353 VDD.n1242 4.5005
R86769 VDD.n1333 VDD.n1242 4.5005
R86770 VDD.n1354 VDD.n1242 4.5005
R86771 VDD.n1332 VDD.n1242 4.5005
R86772 VDD.n1356 VDD.n1242 4.5005
R86773 VDD.n1331 VDD.n1242 4.5005
R86774 VDD.n1357 VDD.n1242 4.5005
R86775 VDD.n1330 VDD.n1242 4.5005
R86776 VDD.n1359 VDD.n1242 4.5005
R86777 VDD.n1329 VDD.n1242 4.5005
R86778 VDD.n1360 VDD.n1242 4.5005
R86779 VDD.n1328 VDD.n1242 4.5005
R86780 VDD.n1362 VDD.n1242 4.5005
R86781 VDD.n1327 VDD.n1242 4.5005
R86782 VDD.n1363 VDD.n1242 4.5005
R86783 VDD.n1326 VDD.n1242 4.5005
R86784 VDD.n1365 VDD.n1242 4.5005
R86785 VDD.n1325 VDD.n1242 4.5005
R86786 VDD.n1366 VDD.n1242 4.5005
R86787 VDD.n1324 VDD.n1242 4.5005
R86788 VDD.n1368 VDD.n1242 4.5005
R86789 VDD.n1323 VDD.n1242 4.5005
R86790 VDD.n1369 VDD.n1242 4.5005
R86791 VDD.n1322 VDD.n1242 4.5005
R86792 VDD.n1371 VDD.n1242 4.5005
R86793 VDD.n1321 VDD.n1242 4.5005
R86794 VDD.n1372 VDD.n1242 4.5005
R86795 VDD.n1320 VDD.n1242 4.5005
R86796 VDD.n1374 VDD.n1242 4.5005
R86797 VDD.n1319 VDD.n1242 4.5005
R86798 VDD.n1375 VDD.n1242 4.5005
R86799 VDD.n1318 VDD.n1242 4.5005
R86800 VDD.n1376 VDD.n1242 4.5005
R86801 VDD.n1316 VDD.n1242 4.5005
R86802 VDD.n1377 VDD.n1242 4.5005
R86803 VDD.n1315 VDD.n1242 4.5005
R86804 VDD.n1378 VDD.n1242 4.5005
R86805 VDD.n1313 VDD.n1242 4.5005
R86806 VDD.n1379 VDD.n1242 4.5005
R86807 VDD.n1312 VDD.n1242 4.5005
R86808 VDD.n1380 VDD.n1242 4.5005
R86809 VDD.n1310 VDD.n1242 4.5005
R86810 VDD.n1381 VDD.n1242 4.5005
R86811 VDD.n1309 VDD.n1242 4.5005
R86812 VDD.n1382 VDD.n1242 4.5005
R86813 VDD.n1307 VDD.n1242 4.5005
R86814 VDD.n1383 VDD.n1242 4.5005
R86815 VDD.n1306 VDD.n1242 4.5005
R86816 VDD.n1384 VDD.n1242 4.5005
R86817 VDD.n1304 VDD.n1242 4.5005
R86818 VDD.n1385 VDD.n1242 4.5005
R86819 VDD.n1303 VDD.n1242 4.5005
R86820 VDD.n1386 VDD.n1242 4.5005
R86821 VDD.n1301 VDD.n1242 4.5005
R86822 VDD.n1387 VDD.n1242 4.5005
R86823 VDD.n1300 VDD.n1242 4.5005
R86824 VDD.n1388 VDD.n1242 4.5005
R86825 VDD.n1298 VDD.n1242 4.5005
R86826 VDD.n1389 VDD.n1242 4.5005
R86827 VDD.n1297 VDD.n1242 4.5005
R86828 VDD.n1390 VDD.n1242 4.5005
R86829 VDD.n1295 VDD.n1242 4.5005
R86830 VDD.n1391 VDD.n1242 4.5005
R86831 VDD.n1294 VDD.n1242 4.5005
R86832 VDD.n1392 VDD.n1242 4.5005
R86833 VDD.n1292 VDD.n1242 4.5005
R86834 VDD.n1393 VDD.n1242 4.5005
R86835 VDD.n1291 VDD.n1242 4.5005
R86836 VDD.n1394 VDD.n1242 4.5005
R86837 VDD.n1289 VDD.n1242 4.5005
R86838 VDD.n1395 VDD.n1242 4.5005
R86839 VDD.n1288 VDD.n1242 4.5005
R86840 VDD.n1396 VDD.n1242 4.5005
R86841 VDD.n1286 VDD.n1242 4.5005
R86842 VDD.n1397 VDD.n1242 4.5005
R86843 VDD.n1285 VDD.n1242 4.5005
R86844 VDD.n1398 VDD.n1242 4.5005
R86845 VDD.n1283 VDD.n1242 4.5005
R86846 VDD.n1399 VDD.n1242 4.5005
R86847 VDD.n1282 VDD.n1242 4.5005
R86848 VDD.n1400 VDD.n1242 4.5005
R86849 VDD.n1280 VDD.n1242 4.5005
R86850 VDD.n1401 VDD.n1242 4.5005
R86851 VDD.n1279 VDD.n1242 4.5005
R86852 VDD.n1402 VDD.n1242 4.5005
R86853 VDD.n1277 VDD.n1242 4.5005
R86854 VDD.n1403 VDD.n1242 4.5005
R86855 VDD.n1276 VDD.n1242 4.5005
R86856 VDD.n1404 VDD.n1242 4.5005
R86857 VDD.n1274 VDD.n1242 4.5005
R86858 VDD.n1405 VDD.n1242 4.5005
R86859 VDD.n1273 VDD.n1242 4.5005
R86860 VDD.n1406 VDD.n1242 4.5005
R86861 VDD.n1271 VDD.n1242 4.5005
R86862 VDD.n1407 VDD.n1242 4.5005
R86863 VDD.n1270 VDD.n1242 4.5005
R86864 VDD.n1408 VDD.n1242 4.5005
R86865 VDD.n1268 VDD.n1242 4.5005
R86866 VDD.n1409 VDD.n1242 4.5005
R86867 VDD.n1267 VDD.n1242 4.5005
R86868 VDD.n1410 VDD.n1242 4.5005
R86869 VDD.n1265 VDD.n1242 4.5005
R86870 VDD.n1411 VDD.n1242 4.5005
R86871 VDD.n1264 VDD.n1242 4.5005
R86872 VDD.n1412 VDD.n1242 4.5005
R86873 VDD.n1262 VDD.n1242 4.5005
R86874 VDD.n1413 VDD.n1242 4.5005
R86875 VDD.n1261 VDD.n1242 4.5005
R86876 VDD.n1414 VDD.n1242 4.5005
R86877 VDD.n1415 VDD.n1242 4.5005
R86878 VDD.n1674 VDD.n1242 4.5005
R86879 VDD.n1676 VDD.n1147 4.5005
R86880 VDD.n1341 VDD.n1147 4.5005
R86881 VDD.n1342 VDD.n1147 4.5005
R86882 VDD.n1340 VDD.n1147 4.5005
R86883 VDD.n1344 VDD.n1147 4.5005
R86884 VDD.n1339 VDD.n1147 4.5005
R86885 VDD.n1345 VDD.n1147 4.5005
R86886 VDD.n1338 VDD.n1147 4.5005
R86887 VDD.n1347 VDD.n1147 4.5005
R86888 VDD.n1337 VDD.n1147 4.5005
R86889 VDD.n1348 VDD.n1147 4.5005
R86890 VDD.n1336 VDD.n1147 4.5005
R86891 VDD.n1350 VDD.n1147 4.5005
R86892 VDD.n1335 VDD.n1147 4.5005
R86893 VDD.n1351 VDD.n1147 4.5005
R86894 VDD.n1334 VDD.n1147 4.5005
R86895 VDD.n1353 VDD.n1147 4.5005
R86896 VDD.n1333 VDD.n1147 4.5005
R86897 VDD.n1354 VDD.n1147 4.5005
R86898 VDD.n1332 VDD.n1147 4.5005
R86899 VDD.n1356 VDD.n1147 4.5005
R86900 VDD.n1331 VDD.n1147 4.5005
R86901 VDD.n1357 VDD.n1147 4.5005
R86902 VDD.n1330 VDD.n1147 4.5005
R86903 VDD.n1359 VDD.n1147 4.5005
R86904 VDD.n1329 VDD.n1147 4.5005
R86905 VDD.n1360 VDD.n1147 4.5005
R86906 VDD.n1328 VDD.n1147 4.5005
R86907 VDD.n1362 VDD.n1147 4.5005
R86908 VDD.n1327 VDD.n1147 4.5005
R86909 VDD.n1363 VDD.n1147 4.5005
R86910 VDD.n1326 VDD.n1147 4.5005
R86911 VDD.n1365 VDD.n1147 4.5005
R86912 VDD.n1325 VDD.n1147 4.5005
R86913 VDD.n1366 VDD.n1147 4.5005
R86914 VDD.n1324 VDD.n1147 4.5005
R86915 VDD.n1368 VDD.n1147 4.5005
R86916 VDD.n1323 VDD.n1147 4.5005
R86917 VDD.n1369 VDD.n1147 4.5005
R86918 VDD.n1322 VDD.n1147 4.5005
R86919 VDD.n1371 VDD.n1147 4.5005
R86920 VDD.n1321 VDD.n1147 4.5005
R86921 VDD.n1372 VDD.n1147 4.5005
R86922 VDD.n1320 VDD.n1147 4.5005
R86923 VDD.n1374 VDD.n1147 4.5005
R86924 VDD.n1319 VDD.n1147 4.5005
R86925 VDD.n1375 VDD.n1147 4.5005
R86926 VDD.n1318 VDD.n1147 4.5005
R86927 VDD.n1376 VDD.n1147 4.5005
R86928 VDD.n1316 VDD.n1147 4.5005
R86929 VDD.n1377 VDD.n1147 4.5005
R86930 VDD.n1315 VDD.n1147 4.5005
R86931 VDD.n1378 VDD.n1147 4.5005
R86932 VDD.n1313 VDD.n1147 4.5005
R86933 VDD.n1379 VDD.n1147 4.5005
R86934 VDD.n1312 VDD.n1147 4.5005
R86935 VDD.n1380 VDD.n1147 4.5005
R86936 VDD.n1310 VDD.n1147 4.5005
R86937 VDD.n1381 VDD.n1147 4.5005
R86938 VDD.n1309 VDD.n1147 4.5005
R86939 VDD.n1382 VDD.n1147 4.5005
R86940 VDD.n1307 VDD.n1147 4.5005
R86941 VDD.n1383 VDD.n1147 4.5005
R86942 VDD.n1306 VDD.n1147 4.5005
R86943 VDD.n1384 VDD.n1147 4.5005
R86944 VDD.n1304 VDD.n1147 4.5005
R86945 VDD.n1385 VDD.n1147 4.5005
R86946 VDD.n1303 VDD.n1147 4.5005
R86947 VDD.n1386 VDD.n1147 4.5005
R86948 VDD.n1301 VDD.n1147 4.5005
R86949 VDD.n1387 VDD.n1147 4.5005
R86950 VDD.n1300 VDD.n1147 4.5005
R86951 VDD.n1388 VDD.n1147 4.5005
R86952 VDD.n1298 VDD.n1147 4.5005
R86953 VDD.n1389 VDD.n1147 4.5005
R86954 VDD.n1297 VDD.n1147 4.5005
R86955 VDD.n1390 VDD.n1147 4.5005
R86956 VDD.n1295 VDD.n1147 4.5005
R86957 VDD.n1391 VDD.n1147 4.5005
R86958 VDD.n1294 VDD.n1147 4.5005
R86959 VDD.n1392 VDD.n1147 4.5005
R86960 VDD.n1292 VDD.n1147 4.5005
R86961 VDD.n1393 VDD.n1147 4.5005
R86962 VDD.n1291 VDD.n1147 4.5005
R86963 VDD.n1394 VDD.n1147 4.5005
R86964 VDD.n1289 VDD.n1147 4.5005
R86965 VDD.n1395 VDD.n1147 4.5005
R86966 VDD.n1288 VDD.n1147 4.5005
R86967 VDD.n1396 VDD.n1147 4.5005
R86968 VDD.n1286 VDD.n1147 4.5005
R86969 VDD.n1397 VDD.n1147 4.5005
R86970 VDD.n1285 VDD.n1147 4.5005
R86971 VDD.n1398 VDD.n1147 4.5005
R86972 VDD.n1283 VDD.n1147 4.5005
R86973 VDD.n1399 VDD.n1147 4.5005
R86974 VDD.n1282 VDD.n1147 4.5005
R86975 VDD.n1400 VDD.n1147 4.5005
R86976 VDD.n1280 VDD.n1147 4.5005
R86977 VDD.n1401 VDD.n1147 4.5005
R86978 VDD.n1279 VDD.n1147 4.5005
R86979 VDD.n1402 VDD.n1147 4.5005
R86980 VDD.n1277 VDD.n1147 4.5005
R86981 VDD.n1403 VDD.n1147 4.5005
R86982 VDD.n1276 VDD.n1147 4.5005
R86983 VDD.n1404 VDD.n1147 4.5005
R86984 VDD.n1274 VDD.n1147 4.5005
R86985 VDD.n1405 VDD.n1147 4.5005
R86986 VDD.n1273 VDD.n1147 4.5005
R86987 VDD.n1406 VDD.n1147 4.5005
R86988 VDD.n1271 VDD.n1147 4.5005
R86989 VDD.n1407 VDD.n1147 4.5005
R86990 VDD.n1270 VDD.n1147 4.5005
R86991 VDD.n1408 VDD.n1147 4.5005
R86992 VDD.n1268 VDD.n1147 4.5005
R86993 VDD.n1409 VDD.n1147 4.5005
R86994 VDD.n1267 VDD.n1147 4.5005
R86995 VDD.n1410 VDD.n1147 4.5005
R86996 VDD.n1265 VDD.n1147 4.5005
R86997 VDD.n1411 VDD.n1147 4.5005
R86998 VDD.n1264 VDD.n1147 4.5005
R86999 VDD.n1412 VDD.n1147 4.5005
R87000 VDD.n1262 VDD.n1147 4.5005
R87001 VDD.n1413 VDD.n1147 4.5005
R87002 VDD.n1261 VDD.n1147 4.5005
R87003 VDD.n1414 VDD.n1147 4.5005
R87004 VDD.n1415 VDD.n1147 4.5005
R87005 VDD.n1674 VDD.n1147 4.5005
R87006 VDD.n1676 VDD.n1243 4.5005
R87007 VDD.n1341 VDD.n1243 4.5005
R87008 VDD.n1342 VDD.n1243 4.5005
R87009 VDD.n1340 VDD.n1243 4.5005
R87010 VDD.n1344 VDD.n1243 4.5005
R87011 VDD.n1339 VDD.n1243 4.5005
R87012 VDD.n1345 VDD.n1243 4.5005
R87013 VDD.n1338 VDD.n1243 4.5005
R87014 VDD.n1347 VDD.n1243 4.5005
R87015 VDD.n1337 VDD.n1243 4.5005
R87016 VDD.n1348 VDD.n1243 4.5005
R87017 VDD.n1336 VDD.n1243 4.5005
R87018 VDD.n1350 VDD.n1243 4.5005
R87019 VDD.n1335 VDD.n1243 4.5005
R87020 VDD.n1351 VDD.n1243 4.5005
R87021 VDD.n1334 VDD.n1243 4.5005
R87022 VDD.n1353 VDD.n1243 4.5005
R87023 VDD.n1333 VDD.n1243 4.5005
R87024 VDD.n1354 VDD.n1243 4.5005
R87025 VDD.n1332 VDD.n1243 4.5005
R87026 VDD.n1356 VDD.n1243 4.5005
R87027 VDD.n1331 VDD.n1243 4.5005
R87028 VDD.n1357 VDD.n1243 4.5005
R87029 VDD.n1330 VDD.n1243 4.5005
R87030 VDD.n1359 VDD.n1243 4.5005
R87031 VDD.n1329 VDD.n1243 4.5005
R87032 VDD.n1360 VDD.n1243 4.5005
R87033 VDD.n1328 VDD.n1243 4.5005
R87034 VDD.n1362 VDD.n1243 4.5005
R87035 VDD.n1327 VDD.n1243 4.5005
R87036 VDD.n1363 VDD.n1243 4.5005
R87037 VDD.n1326 VDD.n1243 4.5005
R87038 VDD.n1365 VDD.n1243 4.5005
R87039 VDD.n1325 VDD.n1243 4.5005
R87040 VDD.n1366 VDD.n1243 4.5005
R87041 VDD.n1324 VDD.n1243 4.5005
R87042 VDD.n1368 VDD.n1243 4.5005
R87043 VDD.n1323 VDD.n1243 4.5005
R87044 VDD.n1369 VDD.n1243 4.5005
R87045 VDD.n1322 VDD.n1243 4.5005
R87046 VDD.n1371 VDD.n1243 4.5005
R87047 VDD.n1321 VDD.n1243 4.5005
R87048 VDD.n1372 VDD.n1243 4.5005
R87049 VDD.n1320 VDD.n1243 4.5005
R87050 VDD.n1374 VDD.n1243 4.5005
R87051 VDD.n1319 VDD.n1243 4.5005
R87052 VDD.n1375 VDD.n1243 4.5005
R87053 VDD.n1318 VDD.n1243 4.5005
R87054 VDD.n1376 VDD.n1243 4.5005
R87055 VDD.n1316 VDD.n1243 4.5005
R87056 VDD.n1377 VDD.n1243 4.5005
R87057 VDD.n1315 VDD.n1243 4.5005
R87058 VDD.n1378 VDD.n1243 4.5005
R87059 VDD.n1313 VDD.n1243 4.5005
R87060 VDD.n1379 VDD.n1243 4.5005
R87061 VDD.n1312 VDD.n1243 4.5005
R87062 VDD.n1380 VDD.n1243 4.5005
R87063 VDD.n1310 VDD.n1243 4.5005
R87064 VDD.n1381 VDD.n1243 4.5005
R87065 VDD.n1309 VDD.n1243 4.5005
R87066 VDD.n1382 VDD.n1243 4.5005
R87067 VDD.n1307 VDD.n1243 4.5005
R87068 VDD.n1383 VDD.n1243 4.5005
R87069 VDD.n1306 VDD.n1243 4.5005
R87070 VDD.n1384 VDD.n1243 4.5005
R87071 VDD.n1304 VDD.n1243 4.5005
R87072 VDD.n1385 VDD.n1243 4.5005
R87073 VDD.n1303 VDD.n1243 4.5005
R87074 VDD.n1386 VDD.n1243 4.5005
R87075 VDD.n1301 VDD.n1243 4.5005
R87076 VDD.n1387 VDD.n1243 4.5005
R87077 VDD.n1300 VDD.n1243 4.5005
R87078 VDD.n1388 VDD.n1243 4.5005
R87079 VDD.n1298 VDD.n1243 4.5005
R87080 VDD.n1389 VDD.n1243 4.5005
R87081 VDD.n1297 VDD.n1243 4.5005
R87082 VDD.n1390 VDD.n1243 4.5005
R87083 VDD.n1295 VDD.n1243 4.5005
R87084 VDD.n1391 VDD.n1243 4.5005
R87085 VDD.n1294 VDD.n1243 4.5005
R87086 VDD.n1392 VDD.n1243 4.5005
R87087 VDD.n1292 VDD.n1243 4.5005
R87088 VDD.n1393 VDD.n1243 4.5005
R87089 VDD.n1291 VDD.n1243 4.5005
R87090 VDD.n1394 VDD.n1243 4.5005
R87091 VDD.n1289 VDD.n1243 4.5005
R87092 VDD.n1395 VDD.n1243 4.5005
R87093 VDD.n1288 VDD.n1243 4.5005
R87094 VDD.n1396 VDD.n1243 4.5005
R87095 VDD.n1286 VDD.n1243 4.5005
R87096 VDD.n1397 VDD.n1243 4.5005
R87097 VDD.n1285 VDD.n1243 4.5005
R87098 VDD.n1398 VDD.n1243 4.5005
R87099 VDD.n1283 VDD.n1243 4.5005
R87100 VDD.n1399 VDD.n1243 4.5005
R87101 VDD.n1282 VDD.n1243 4.5005
R87102 VDD.n1400 VDD.n1243 4.5005
R87103 VDD.n1280 VDD.n1243 4.5005
R87104 VDD.n1401 VDD.n1243 4.5005
R87105 VDD.n1279 VDD.n1243 4.5005
R87106 VDD.n1402 VDD.n1243 4.5005
R87107 VDD.n1277 VDD.n1243 4.5005
R87108 VDD.n1403 VDD.n1243 4.5005
R87109 VDD.n1276 VDD.n1243 4.5005
R87110 VDD.n1404 VDD.n1243 4.5005
R87111 VDD.n1274 VDD.n1243 4.5005
R87112 VDD.n1405 VDD.n1243 4.5005
R87113 VDD.n1273 VDD.n1243 4.5005
R87114 VDD.n1406 VDD.n1243 4.5005
R87115 VDD.n1271 VDD.n1243 4.5005
R87116 VDD.n1407 VDD.n1243 4.5005
R87117 VDD.n1270 VDD.n1243 4.5005
R87118 VDD.n1408 VDD.n1243 4.5005
R87119 VDD.n1268 VDD.n1243 4.5005
R87120 VDD.n1409 VDD.n1243 4.5005
R87121 VDD.n1267 VDD.n1243 4.5005
R87122 VDD.n1410 VDD.n1243 4.5005
R87123 VDD.n1265 VDD.n1243 4.5005
R87124 VDD.n1411 VDD.n1243 4.5005
R87125 VDD.n1264 VDD.n1243 4.5005
R87126 VDD.n1412 VDD.n1243 4.5005
R87127 VDD.n1262 VDD.n1243 4.5005
R87128 VDD.n1413 VDD.n1243 4.5005
R87129 VDD.n1261 VDD.n1243 4.5005
R87130 VDD.n1414 VDD.n1243 4.5005
R87131 VDD.n1415 VDD.n1243 4.5005
R87132 VDD.n1674 VDD.n1243 4.5005
R87133 VDD.n1676 VDD.n1146 4.5005
R87134 VDD.n1341 VDD.n1146 4.5005
R87135 VDD.n1342 VDD.n1146 4.5005
R87136 VDD.n1340 VDD.n1146 4.5005
R87137 VDD.n1344 VDD.n1146 4.5005
R87138 VDD.n1339 VDD.n1146 4.5005
R87139 VDD.n1345 VDD.n1146 4.5005
R87140 VDD.n1338 VDD.n1146 4.5005
R87141 VDD.n1347 VDD.n1146 4.5005
R87142 VDD.n1337 VDD.n1146 4.5005
R87143 VDD.n1348 VDD.n1146 4.5005
R87144 VDD.n1336 VDD.n1146 4.5005
R87145 VDD.n1350 VDD.n1146 4.5005
R87146 VDD.n1335 VDD.n1146 4.5005
R87147 VDD.n1351 VDD.n1146 4.5005
R87148 VDD.n1334 VDD.n1146 4.5005
R87149 VDD.n1353 VDD.n1146 4.5005
R87150 VDD.n1333 VDD.n1146 4.5005
R87151 VDD.n1354 VDD.n1146 4.5005
R87152 VDD.n1332 VDD.n1146 4.5005
R87153 VDD.n1356 VDD.n1146 4.5005
R87154 VDD.n1331 VDD.n1146 4.5005
R87155 VDD.n1357 VDD.n1146 4.5005
R87156 VDD.n1330 VDD.n1146 4.5005
R87157 VDD.n1359 VDD.n1146 4.5005
R87158 VDD.n1329 VDD.n1146 4.5005
R87159 VDD.n1360 VDD.n1146 4.5005
R87160 VDD.n1328 VDD.n1146 4.5005
R87161 VDD.n1362 VDD.n1146 4.5005
R87162 VDD.n1327 VDD.n1146 4.5005
R87163 VDD.n1363 VDD.n1146 4.5005
R87164 VDD.n1326 VDD.n1146 4.5005
R87165 VDD.n1365 VDD.n1146 4.5005
R87166 VDD.n1325 VDD.n1146 4.5005
R87167 VDD.n1366 VDD.n1146 4.5005
R87168 VDD.n1324 VDD.n1146 4.5005
R87169 VDD.n1368 VDD.n1146 4.5005
R87170 VDD.n1323 VDD.n1146 4.5005
R87171 VDD.n1369 VDD.n1146 4.5005
R87172 VDD.n1322 VDD.n1146 4.5005
R87173 VDD.n1371 VDD.n1146 4.5005
R87174 VDD.n1321 VDD.n1146 4.5005
R87175 VDD.n1372 VDD.n1146 4.5005
R87176 VDD.n1320 VDD.n1146 4.5005
R87177 VDD.n1374 VDD.n1146 4.5005
R87178 VDD.n1319 VDD.n1146 4.5005
R87179 VDD.n1375 VDD.n1146 4.5005
R87180 VDD.n1318 VDD.n1146 4.5005
R87181 VDD.n1376 VDD.n1146 4.5005
R87182 VDD.n1316 VDD.n1146 4.5005
R87183 VDD.n1377 VDD.n1146 4.5005
R87184 VDD.n1315 VDD.n1146 4.5005
R87185 VDD.n1378 VDD.n1146 4.5005
R87186 VDD.n1313 VDD.n1146 4.5005
R87187 VDD.n1379 VDD.n1146 4.5005
R87188 VDD.n1312 VDD.n1146 4.5005
R87189 VDD.n1380 VDD.n1146 4.5005
R87190 VDD.n1310 VDD.n1146 4.5005
R87191 VDD.n1381 VDD.n1146 4.5005
R87192 VDD.n1309 VDD.n1146 4.5005
R87193 VDD.n1382 VDD.n1146 4.5005
R87194 VDD.n1307 VDD.n1146 4.5005
R87195 VDD.n1383 VDD.n1146 4.5005
R87196 VDD.n1306 VDD.n1146 4.5005
R87197 VDD.n1384 VDD.n1146 4.5005
R87198 VDD.n1304 VDD.n1146 4.5005
R87199 VDD.n1385 VDD.n1146 4.5005
R87200 VDD.n1303 VDD.n1146 4.5005
R87201 VDD.n1386 VDD.n1146 4.5005
R87202 VDD.n1301 VDD.n1146 4.5005
R87203 VDD.n1387 VDD.n1146 4.5005
R87204 VDD.n1300 VDD.n1146 4.5005
R87205 VDD.n1388 VDD.n1146 4.5005
R87206 VDD.n1298 VDD.n1146 4.5005
R87207 VDD.n1389 VDD.n1146 4.5005
R87208 VDD.n1297 VDD.n1146 4.5005
R87209 VDD.n1390 VDD.n1146 4.5005
R87210 VDD.n1295 VDD.n1146 4.5005
R87211 VDD.n1391 VDD.n1146 4.5005
R87212 VDD.n1294 VDD.n1146 4.5005
R87213 VDD.n1392 VDD.n1146 4.5005
R87214 VDD.n1292 VDD.n1146 4.5005
R87215 VDD.n1393 VDD.n1146 4.5005
R87216 VDD.n1291 VDD.n1146 4.5005
R87217 VDD.n1394 VDD.n1146 4.5005
R87218 VDD.n1289 VDD.n1146 4.5005
R87219 VDD.n1395 VDD.n1146 4.5005
R87220 VDD.n1288 VDD.n1146 4.5005
R87221 VDD.n1396 VDD.n1146 4.5005
R87222 VDD.n1286 VDD.n1146 4.5005
R87223 VDD.n1397 VDD.n1146 4.5005
R87224 VDD.n1285 VDD.n1146 4.5005
R87225 VDD.n1398 VDD.n1146 4.5005
R87226 VDD.n1283 VDD.n1146 4.5005
R87227 VDD.n1399 VDD.n1146 4.5005
R87228 VDD.n1282 VDD.n1146 4.5005
R87229 VDD.n1400 VDD.n1146 4.5005
R87230 VDD.n1280 VDD.n1146 4.5005
R87231 VDD.n1401 VDD.n1146 4.5005
R87232 VDD.n1279 VDD.n1146 4.5005
R87233 VDD.n1402 VDD.n1146 4.5005
R87234 VDD.n1277 VDD.n1146 4.5005
R87235 VDD.n1403 VDD.n1146 4.5005
R87236 VDD.n1276 VDD.n1146 4.5005
R87237 VDD.n1404 VDD.n1146 4.5005
R87238 VDD.n1274 VDD.n1146 4.5005
R87239 VDD.n1405 VDD.n1146 4.5005
R87240 VDD.n1273 VDD.n1146 4.5005
R87241 VDD.n1406 VDD.n1146 4.5005
R87242 VDD.n1271 VDD.n1146 4.5005
R87243 VDD.n1407 VDD.n1146 4.5005
R87244 VDD.n1270 VDD.n1146 4.5005
R87245 VDD.n1408 VDD.n1146 4.5005
R87246 VDD.n1268 VDD.n1146 4.5005
R87247 VDD.n1409 VDD.n1146 4.5005
R87248 VDD.n1267 VDD.n1146 4.5005
R87249 VDD.n1410 VDD.n1146 4.5005
R87250 VDD.n1265 VDD.n1146 4.5005
R87251 VDD.n1411 VDD.n1146 4.5005
R87252 VDD.n1264 VDD.n1146 4.5005
R87253 VDD.n1412 VDD.n1146 4.5005
R87254 VDD.n1262 VDD.n1146 4.5005
R87255 VDD.n1413 VDD.n1146 4.5005
R87256 VDD.n1261 VDD.n1146 4.5005
R87257 VDD.n1414 VDD.n1146 4.5005
R87258 VDD.n1415 VDD.n1146 4.5005
R87259 VDD.n1674 VDD.n1146 4.5005
R87260 VDD.n1676 VDD.n1244 4.5005
R87261 VDD.n1341 VDD.n1244 4.5005
R87262 VDD.n1342 VDD.n1244 4.5005
R87263 VDD.n1340 VDD.n1244 4.5005
R87264 VDD.n1344 VDD.n1244 4.5005
R87265 VDD.n1339 VDD.n1244 4.5005
R87266 VDD.n1345 VDD.n1244 4.5005
R87267 VDD.n1338 VDD.n1244 4.5005
R87268 VDD.n1347 VDD.n1244 4.5005
R87269 VDD.n1337 VDD.n1244 4.5005
R87270 VDD.n1348 VDD.n1244 4.5005
R87271 VDD.n1336 VDD.n1244 4.5005
R87272 VDD.n1350 VDD.n1244 4.5005
R87273 VDD.n1335 VDD.n1244 4.5005
R87274 VDD.n1351 VDD.n1244 4.5005
R87275 VDD.n1334 VDD.n1244 4.5005
R87276 VDD.n1353 VDD.n1244 4.5005
R87277 VDD.n1333 VDD.n1244 4.5005
R87278 VDD.n1354 VDD.n1244 4.5005
R87279 VDD.n1332 VDD.n1244 4.5005
R87280 VDD.n1356 VDD.n1244 4.5005
R87281 VDD.n1331 VDD.n1244 4.5005
R87282 VDD.n1357 VDD.n1244 4.5005
R87283 VDD.n1330 VDD.n1244 4.5005
R87284 VDD.n1359 VDD.n1244 4.5005
R87285 VDD.n1329 VDD.n1244 4.5005
R87286 VDD.n1360 VDD.n1244 4.5005
R87287 VDD.n1328 VDD.n1244 4.5005
R87288 VDD.n1362 VDD.n1244 4.5005
R87289 VDD.n1327 VDD.n1244 4.5005
R87290 VDD.n1363 VDD.n1244 4.5005
R87291 VDD.n1326 VDD.n1244 4.5005
R87292 VDD.n1365 VDD.n1244 4.5005
R87293 VDD.n1325 VDD.n1244 4.5005
R87294 VDD.n1366 VDD.n1244 4.5005
R87295 VDD.n1324 VDD.n1244 4.5005
R87296 VDD.n1368 VDD.n1244 4.5005
R87297 VDD.n1323 VDD.n1244 4.5005
R87298 VDD.n1369 VDD.n1244 4.5005
R87299 VDD.n1322 VDD.n1244 4.5005
R87300 VDD.n1371 VDD.n1244 4.5005
R87301 VDD.n1321 VDD.n1244 4.5005
R87302 VDD.n1372 VDD.n1244 4.5005
R87303 VDD.n1320 VDD.n1244 4.5005
R87304 VDD.n1374 VDD.n1244 4.5005
R87305 VDD.n1319 VDD.n1244 4.5005
R87306 VDD.n1375 VDD.n1244 4.5005
R87307 VDD.n1318 VDD.n1244 4.5005
R87308 VDD.n1376 VDD.n1244 4.5005
R87309 VDD.n1316 VDD.n1244 4.5005
R87310 VDD.n1377 VDD.n1244 4.5005
R87311 VDD.n1315 VDD.n1244 4.5005
R87312 VDD.n1378 VDD.n1244 4.5005
R87313 VDD.n1313 VDD.n1244 4.5005
R87314 VDD.n1379 VDD.n1244 4.5005
R87315 VDD.n1312 VDD.n1244 4.5005
R87316 VDD.n1380 VDD.n1244 4.5005
R87317 VDD.n1310 VDD.n1244 4.5005
R87318 VDD.n1381 VDD.n1244 4.5005
R87319 VDD.n1309 VDD.n1244 4.5005
R87320 VDD.n1382 VDD.n1244 4.5005
R87321 VDD.n1307 VDD.n1244 4.5005
R87322 VDD.n1383 VDD.n1244 4.5005
R87323 VDD.n1306 VDD.n1244 4.5005
R87324 VDD.n1384 VDD.n1244 4.5005
R87325 VDD.n1304 VDD.n1244 4.5005
R87326 VDD.n1385 VDD.n1244 4.5005
R87327 VDD.n1303 VDD.n1244 4.5005
R87328 VDD.n1386 VDD.n1244 4.5005
R87329 VDD.n1301 VDD.n1244 4.5005
R87330 VDD.n1387 VDD.n1244 4.5005
R87331 VDD.n1300 VDD.n1244 4.5005
R87332 VDD.n1388 VDD.n1244 4.5005
R87333 VDD.n1298 VDD.n1244 4.5005
R87334 VDD.n1389 VDD.n1244 4.5005
R87335 VDD.n1297 VDD.n1244 4.5005
R87336 VDD.n1390 VDD.n1244 4.5005
R87337 VDD.n1295 VDD.n1244 4.5005
R87338 VDD.n1391 VDD.n1244 4.5005
R87339 VDD.n1294 VDD.n1244 4.5005
R87340 VDD.n1392 VDD.n1244 4.5005
R87341 VDD.n1292 VDD.n1244 4.5005
R87342 VDD.n1393 VDD.n1244 4.5005
R87343 VDD.n1291 VDD.n1244 4.5005
R87344 VDD.n1394 VDD.n1244 4.5005
R87345 VDD.n1289 VDD.n1244 4.5005
R87346 VDD.n1395 VDD.n1244 4.5005
R87347 VDD.n1288 VDD.n1244 4.5005
R87348 VDD.n1396 VDD.n1244 4.5005
R87349 VDD.n1286 VDD.n1244 4.5005
R87350 VDD.n1397 VDD.n1244 4.5005
R87351 VDD.n1285 VDD.n1244 4.5005
R87352 VDD.n1398 VDD.n1244 4.5005
R87353 VDD.n1283 VDD.n1244 4.5005
R87354 VDD.n1399 VDD.n1244 4.5005
R87355 VDD.n1282 VDD.n1244 4.5005
R87356 VDD.n1400 VDD.n1244 4.5005
R87357 VDD.n1280 VDD.n1244 4.5005
R87358 VDD.n1401 VDD.n1244 4.5005
R87359 VDD.n1279 VDD.n1244 4.5005
R87360 VDD.n1402 VDD.n1244 4.5005
R87361 VDD.n1277 VDD.n1244 4.5005
R87362 VDD.n1403 VDD.n1244 4.5005
R87363 VDD.n1276 VDD.n1244 4.5005
R87364 VDD.n1404 VDD.n1244 4.5005
R87365 VDD.n1274 VDD.n1244 4.5005
R87366 VDD.n1405 VDD.n1244 4.5005
R87367 VDD.n1273 VDD.n1244 4.5005
R87368 VDD.n1406 VDD.n1244 4.5005
R87369 VDD.n1271 VDD.n1244 4.5005
R87370 VDD.n1407 VDD.n1244 4.5005
R87371 VDD.n1270 VDD.n1244 4.5005
R87372 VDD.n1408 VDD.n1244 4.5005
R87373 VDD.n1268 VDD.n1244 4.5005
R87374 VDD.n1409 VDD.n1244 4.5005
R87375 VDD.n1267 VDD.n1244 4.5005
R87376 VDD.n1410 VDD.n1244 4.5005
R87377 VDD.n1265 VDD.n1244 4.5005
R87378 VDD.n1411 VDD.n1244 4.5005
R87379 VDD.n1264 VDD.n1244 4.5005
R87380 VDD.n1412 VDD.n1244 4.5005
R87381 VDD.n1262 VDD.n1244 4.5005
R87382 VDD.n1413 VDD.n1244 4.5005
R87383 VDD.n1261 VDD.n1244 4.5005
R87384 VDD.n1414 VDD.n1244 4.5005
R87385 VDD.n1415 VDD.n1244 4.5005
R87386 VDD.n1674 VDD.n1244 4.5005
R87387 VDD.n1676 VDD.n1145 4.5005
R87388 VDD.n1341 VDD.n1145 4.5005
R87389 VDD.n1342 VDD.n1145 4.5005
R87390 VDD.n1340 VDD.n1145 4.5005
R87391 VDD.n1344 VDD.n1145 4.5005
R87392 VDD.n1339 VDD.n1145 4.5005
R87393 VDD.n1345 VDD.n1145 4.5005
R87394 VDD.n1338 VDD.n1145 4.5005
R87395 VDD.n1347 VDD.n1145 4.5005
R87396 VDD.n1337 VDD.n1145 4.5005
R87397 VDD.n1348 VDD.n1145 4.5005
R87398 VDD.n1336 VDD.n1145 4.5005
R87399 VDD.n1350 VDD.n1145 4.5005
R87400 VDD.n1335 VDD.n1145 4.5005
R87401 VDD.n1351 VDD.n1145 4.5005
R87402 VDD.n1334 VDD.n1145 4.5005
R87403 VDD.n1353 VDD.n1145 4.5005
R87404 VDD.n1333 VDD.n1145 4.5005
R87405 VDD.n1354 VDD.n1145 4.5005
R87406 VDD.n1332 VDD.n1145 4.5005
R87407 VDD.n1356 VDD.n1145 4.5005
R87408 VDD.n1331 VDD.n1145 4.5005
R87409 VDD.n1357 VDD.n1145 4.5005
R87410 VDD.n1330 VDD.n1145 4.5005
R87411 VDD.n1359 VDD.n1145 4.5005
R87412 VDD.n1329 VDD.n1145 4.5005
R87413 VDD.n1360 VDD.n1145 4.5005
R87414 VDD.n1328 VDD.n1145 4.5005
R87415 VDD.n1362 VDD.n1145 4.5005
R87416 VDD.n1327 VDD.n1145 4.5005
R87417 VDD.n1363 VDD.n1145 4.5005
R87418 VDD.n1326 VDD.n1145 4.5005
R87419 VDD.n1365 VDD.n1145 4.5005
R87420 VDD.n1325 VDD.n1145 4.5005
R87421 VDD.n1366 VDD.n1145 4.5005
R87422 VDD.n1324 VDD.n1145 4.5005
R87423 VDD.n1368 VDD.n1145 4.5005
R87424 VDD.n1323 VDD.n1145 4.5005
R87425 VDD.n1369 VDD.n1145 4.5005
R87426 VDD.n1322 VDD.n1145 4.5005
R87427 VDD.n1371 VDD.n1145 4.5005
R87428 VDD.n1321 VDD.n1145 4.5005
R87429 VDD.n1372 VDD.n1145 4.5005
R87430 VDD.n1320 VDD.n1145 4.5005
R87431 VDD.n1374 VDD.n1145 4.5005
R87432 VDD.n1319 VDD.n1145 4.5005
R87433 VDD.n1375 VDD.n1145 4.5005
R87434 VDD.n1318 VDD.n1145 4.5005
R87435 VDD.n1376 VDD.n1145 4.5005
R87436 VDD.n1316 VDD.n1145 4.5005
R87437 VDD.n1377 VDD.n1145 4.5005
R87438 VDD.n1315 VDD.n1145 4.5005
R87439 VDD.n1378 VDD.n1145 4.5005
R87440 VDD.n1313 VDD.n1145 4.5005
R87441 VDD.n1379 VDD.n1145 4.5005
R87442 VDD.n1312 VDD.n1145 4.5005
R87443 VDD.n1380 VDD.n1145 4.5005
R87444 VDD.n1310 VDD.n1145 4.5005
R87445 VDD.n1381 VDD.n1145 4.5005
R87446 VDD.n1309 VDD.n1145 4.5005
R87447 VDD.n1382 VDD.n1145 4.5005
R87448 VDD.n1307 VDD.n1145 4.5005
R87449 VDD.n1383 VDD.n1145 4.5005
R87450 VDD.n1306 VDD.n1145 4.5005
R87451 VDD.n1384 VDD.n1145 4.5005
R87452 VDD.n1304 VDD.n1145 4.5005
R87453 VDD.n1385 VDD.n1145 4.5005
R87454 VDD.n1303 VDD.n1145 4.5005
R87455 VDD.n1386 VDD.n1145 4.5005
R87456 VDD.n1301 VDD.n1145 4.5005
R87457 VDD.n1387 VDD.n1145 4.5005
R87458 VDD.n1300 VDD.n1145 4.5005
R87459 VDD.n1388 VDD.n1145 4.5005
R87460 VDD.n1298 VDD.n1145 4.5005
R87461 VDD.n1389 VDD.n1145 4.5005
R87462 VDD.n1297 VDD.n1145 4.5005
R87463 VDD.n1390 VDD.n1145 4.5005
R87464 VDD.n1295 VDD.n1145 4.5005
R87465 VDD.n1391 VDD.n1145 4.5005
R87466 VDD.n1294 VDD.n1145 4.5005
R87467 VDD.n1392 VDD.n1145 4.5005
R87468 VDD.n1292 VDD.n1145 4.5005
R87469 VDD.n1393 VDD.n1145 4.5005
R87470 VDD.n1291 VDD.n1145 4.5005
R87471 VDD.n1394 VDD.n1145 4.5005
R87472 VDD.n1289 VDD.n1145 4.5005
R87473 VDD.n1395 VDD.n1145 4.5005
R87474 VDD.n1288 VDD.n1145 4.5005
R87475 VDD.n1396 VDD.n1145 4.5005
R87476 VDD.n1286 VDD.n1145 4.5005
R87477 VDD.n1397 VDD.n1145 4.5005
R87478 VDD.n1285 VDD.n1145 4.5005
R87479 VDD.n1398 VDD.n1145 4.5005
R87480 VDD.n1283 VDD.n1145 4.5005
R87481 VDD.n1399 VDD.n1145 4.5005
R87482 VDD.n1282 VDD.n1145 4.5005
R87483 VDD.n1400 VDD.n1145 4.5005
R87484 VDD.n1280 VDD.n1145 4.5005
R87485 VDD.n1401 VDD.n1145 4.5005
R87486 VDD.n1279 VDD.n1145 4.5005
R87487 VDD.n1402 VDD.n1145 4.5005
R87488 VDD.n1277 VDD.n1145 4.5005
R87489 VDD.n1403 VDD.n1145 4.5005
R87490 VDD.n1276 VDD.n1145 4.5005
R87491 VDD.n1404 VDD.n1145 4.5005
R87492 VDD.n1274 VDD.n1145 4.5005
R87493 VDD.n1405 VDD.n1145 4.5005
R87494 VDD.n1273 VDD.n1145 4.5005
R87495 VDD.n1406 VDD.n1145 4.5005
R87496 VDD.n1271 VDD.n1145 4.5005
R87497 VDD.n1407 VDD.n1145 4.5005
R87498 VDD.n1270 VDD.n1145 4.5005
R87499 VDD.n1408 VDD.n1145 4.5005
R87500 VDD.n1268 VDD.n1145 4.5005
R87501 VDD.n1409 VDD.n1145 4.5005
R87502 VDD.n1267 VDD.n1145 4.5005
R87503 VDD.n1410 VDD.n1145 4.5005
R87504 VDD.n1265 VDD.n1145 4.5005
R87505 VDD.n1411 VDD.n1145 4.5005
R87506 VDD.n1264 VDD.n1145 4.5005
R87507 VDD.n1412 VDD.n1145 4.5005
R87508 VDD.n1262 VDD.n1145 4.5005
R87509 VDD.n1413 VDD.n1145 4.5005
R87510 VDD.n1261 VDD.n1145 4.5005
R87511 VDD.n1414 VDD.n1145 4.5005
R87512 VDD.n1415 VDD.n1145 4.5005
R87513 VDD.n1674 VDD.n1145 4.5005
R87514 VDD.n1676 VDD.n1245 4.5005
R87515 VDD.n1341 VDD.n1245 4.5005
R87516 VDD.n1342 VDD.n1245 4.5005
R87517 VDD.n1340 VDD.n1245 4.5005
R87518 VDD.n1344 VDD.n1245 4.5005
R87519 VDD.n1339 VDD.n1245 4.5005
R87520 VDD.n1345 VDD.n1245 4.5005
R87521 VDD.n1338 VDD.n1245 4.5005
R87522 VDD.n1347 VDD.n1245 4.5005
R87523 VDD.n1337 VDD.n1245 4.5005
R87524 VDD.n1348 VDD.n1245 4.5005
R87525 VDD.n1336 VDD.n1245 4.5005
R87526 VDD.n1350 VDD.n1245 4.5005
R87527 VDD.n1335 VDD.n1245 4.5005
R87528 VDD.n1351 VDD.n1245 4.5005
R87529 VDD.n1334 VDD.n1245 4.5005
R87530 VDD.n1353 VDD.n1245 4.5005
R87531 VDD.n1333 VDD.n1245 4.5005
R87532 VDD.n1354 VDD.n1245 4.5005
R87533 VDD.n1332 VDD.n1245 4.5005
R87534 VDD.n1356 VDD.n1245 4.5005
R87535 VDD.n1331 VDD.n1245 4.5005
R87536 VDD.n1357 VDD.n1245 4.5005
R87537 VDD.n1330 VDD.n1245 4.5005
R87538 VDD.n1359 VDD.n1245 4.5005
R87539 VDD.n1329 VDD.n1245 4.5005
R87540 VDD.n1360 VDD.n1245 4.5005
R87541 VDD.n1328 VDD.n1245 4.5005
R87542 VDD.n1362 VDD.n1245 4.5005
R87543 VDD.n1327 VDD.n1245 4.5005
R87544 VDD.n1363 VDD.n1245 4.5005
R87545 VDD.n1326 VDD.n1245 4.5005
R87546 VDD.n1365 VDD.n1245 4.5005
R87547 VDD.n1325 VDD.n1245 4.5005
R87548 VDD.n1366 VDD.n1245 4.5005
R87549 VDD.n1324 VDD.n1245 4.5005
R87550 VDD.n1368 VDD.n1245 4.5005
R87551 VDD.n1323 VDD.n1245 4.5005
R87552 VDD.n1369 VDD.n1245 4.5005
R87553 VDD.n1322 VDD.n1245 4.5005
R87554 VDD.n1371 VDD.n1245 4.5005
R87555 VDD.n1321 VDD.n1245 4.5005
R87556 VDD.n1372 VDD.n1245 4.5005
R87557 VDD.n1320 VDD.n1245 4.5005
R87558 VDD.n1374 VDD.n1245 4.5005
R87559 VDD.n1319 VDD.n1245 4.5005
R87560 VDD.n1375 VDD.n1245 4.5005
R87561 VDD.n1318 VDD.n1245 4.5005
R87562 VDD.n1376 VDD.n1245 4.5005
R87563 VDD.n1316 VDD.n1245 4.5005
R87564 VDD.n1377 VDD.n1245 4.5005
R87565 VDD.n1315 VDD.n1245 4.5005
R87566 VDD.n1378 VDD.n1245 4.5005
R87567 VDD.n1313 VDD.n1245 4.5005
R87568 VDD.n1379 VDD.n1245 4.5005
R87569 VDD.n1312 VDD.n1245 4.5005
R87570 VDD.n1380 VDD.n1245 4.5005
R87571 VDD.n1310 VDD.n1245 4.5005
R87572 VDD.n1381 VDD.n1245 4.5005
R87573 VDD.n1309 VDD.n1245 4.5005
R87574 VDD.n1382 VDD.n1245 4.5005
R87575 VDD.n1307 VDD.n1245 4.5005
R87576 VDD.n1383 VDD.n1245 4.5005
R87577 VDD.n1306 VDD.n1245 4.5005
R87578 VDD.n1384 VDD.n1245 4.5005
R87579 VDD.n1304 VDD.n1245 4.5005
R87580 VDD.n1385 VDD.n1245 4.5005
R87581 VDD.n1303 VDD.n1245 4.5005
R87582 VDD.n1386 VDD.n1245 4.5005
R87583 VDD.n1301 VDD.n1245 4.5005
R87584 VDD.n1387 VDD.n1245 4.5005
R87585 VDD.n1300 VDD.n1245 4.5005
R87586 VDD.n1388 VDD.n1245 4.5005
R87587 VDD.n1298 VDD.n1245 4.5005
R87588 VDD.n1389 VDD.n1245 4.5005
R87589 VDD.n1297 VDD.n1245 4.5005
R87590 VDD.n1390 VDD.n1245 4.5005
R87591 VDD.n1295 VDD.n1245 4.5005
R87592 VDD.n1391 VDD.n1245 4.5005
R87593 VDD.n1294 VDD.n1245 4.5005
R87594 VDD.n1392 VDD.n1245 4.5005
R87595 VDD.n1292 VDD.n1245 4.5005
R87596 VDD.n1393 VDD.n1245 4.5005
R87597 VDD.n1291 VDD.n1245 4.5005
R87598 VDD.n1394 VDD.n1245 4.5005
R87599 VDD.n1289 VDD.n1245 4.5005
R87600 VDD.n1395 VDD.n1245 4.5005
R87601 VDD.n1288 VDD.n1245 4.5005
R87602 VDD.n1396 VDD.n1245 4.5005
R87603 VDD.n1286 VDD.n1245 4.5005
R87604 VDD.n1397 VDD.n1245 4.5005
R87605 VDD.n1285 VDD.n1245 4.5005
R87606 VDD.n1398 VDD.n1245 4.5005
R87607 VDD.n1283 VDD.n1245 4.5005
R87608 VDD.n1399 VDD.n1245 4.5005
R87609 VDD.n1282 VDD.n1245 4.5005
R87610 VDD.n1400 VDD.n1245 4.5005
R87611 VDD.n1280 VDD.n1245 4.5005
R87612 VDD.n1401 VDD.n1245 4.5005
R87613 VDD.n1279 VDD.n1245 4.5005
R87614 VDD.n1402 VDD.n1245 4.5005
R87615 VDD.n1277 VDD.n1245 4.5005
R87616 VDD.n1403 VDD.n1245 4.5005
R87617 VDD.n1276 VDD.n1245 4.5005
R87618 VDD.n1404 VDD.n1245 4.5005
R87619 VDD.n1274 VDD.n1245 4.5005
R87620 VDD.n1405 VDD.n1245 4.5005
R87621 VDD.n1273 VDD.n1245 4.5005
R87622 VDD.n1406 VDD.n1245 4.5005
R87623 VDD.n1271 VDD.n1245 4.5005
R87624 VDD.n1407 VDD.n1245 4.5005
R87625 VDD.n1270 VDD.n1245 4.5005
R87626 VDD.n1408 VDD.n1245 4.5005
R87627 VDD.n1268 VDD.n1245 4.5005
R87628 VDD.n1409 VDD.n1245 4.5005
R87629 VDD.n1267 VDD.n1245 4.5005
R87630 VDD.n1410 VDD.n1245 4.5005
R87631 VDD.n1265 VDD.n1245 4.5005
R87632 VDD.n1411 VDD.n1245 4.5005
R87633 VDD.n1264 VDD.n1245 4.5005
R87634 VDD.n1412 VDD.n1245 4.5005
R87635 VDD.n1262 VDD.n1245 4.5005
R87636 VDD.n1413 VDD.n1245 4.5005
R87637 VDD.n1261 VDD.n1245 4.5005
R87638 VDD.n1414 VDD.n1245 4.5005
R87639 VDD.n1415 VDD.n1245 4.5005
R87640 VDD.n1674 VDD.n1245 4.5005
R87641 VDD.n1676 VDD.n1144 4.5005
R87642 VDD.n1341 VDD.n1144 4.5005
R87643 VDD.n1342 VDD.n1144 4.5005
R87644 VDD.n1340 VDD.n1144 4.5005
R87645 VDD.n1344 VDD.n1144 4.5005
R87646 VDD.n1339 VDD.n1144 4.5005
R87647 VDD.n1345 VDD.n1144 4.5005
R87648 VDD.n1338 VDD.n1144 4.5005
R87649 VDD.n1347 VDD.n1144 4.5005
R87650 VDD.n1337 VDD.n1144 4.5005
R87651 VDD.n1348 VDD.n1144 4.5005
R87652 VDD.n1336 VDD.n1144 4.5005
R87653 VDD.n1350 VDD.n1144 4.5005
R87654 VDD.n1335 VDD.n1144 4.5005
R87655 VDD.n1351 VDD.n1144 4.5005
R87656 VDD.n1334 VDD.n1144 4.5005
R87657 VDD.n1353 VDD.n1144 4.5005
R87658 VDD.n1333 VDD.n1144 4.5005
R87659 VDD.n1354 VDD.n1144 4.5005
R87660 VDD.n1332 VDD.n1144 4.5005
R87661 VDD.n1356 VDD.n1144 4.5005
R87662 VDD.n1331 VDD.n1144 4.5005
R87663 VDD.n1357 VDD.n1144 4.5005
R87664 VDD.n1330 VDD.n1144 4.5005
R87665 VDD.n1359 VDD.n1144 4.5005
R87666 VDD.n1329 VDD.n1144 4.5005
R87667 VDD.n1360 VDD.n1144 4.5005
R87668 VDD.n1328 VDD.n1144 4.5005
R87669 VDD.n1362 VDD.n1144 4.5005
R87670 VDD.n1327 VDD.n1144 4.5005
R87671 VDD.n1363 VDD.n1144 4.5005
R87672 VDD.n1326 VDD.n1144 4.5005
R87673 VDD.n1365 VDD.n1144 4.5005
R87674 VDD.n1325 VDD.n1144 4.5005
R87675 VDD.n1366 VDD.n1144 4.5005
R87676 VDD.n1324 VDD.n1144 4.5005
R87677 VDD.n1368 VDD.n1144 4.5005
R87678 VDD.n1323 VDD.n1144 4.5005
R87679 VDD.n1369 VDD.n1144 4.5005
R87680 VDD.n1322 VDD.n1144 4.5005
R87681 VDD.n1371 VDD.n1144 4.5005
R87682 VDD.n1321 VDD.n1144 4.5005
R87683 VDD.n1372 VDD.n1144 4.5005
R87684 VDD.n1320 VDD.n1144 4.5005
R87685 VDD.n1374 VDD.n1144 4.5005
R87686 VDD.n1319 VDD.n1144 4.5005
R87687 VDD.n1375 VDD.n1144 4.5005
R87688 VDD.n1318 VDD.n1144 4.5005
R87689 VDD.n1376 VDD.n1144 4.5005
R87690 VDD.n1316 VDD.n1144 4.5005
R87691 VDD.n1377 VDD.n1144 4.5005
R87692 VDD.n1315 VDD.n1144 4.5005
R87693 VDD.n1378 VDD.n1144 4.5005
R87694 VDD.n1313 VDD.n1144 4.5005
R87695 VDD.n1379 VDD.n1144 4.5005
R87696 VDD.n1312 VDD.n1144 4.5005
R87697 VDD.n1380 VDD.n1144 4.5005
R87698 VDD.n1310 VDD.n1144 4.5005
R87699 VDD.n1381 VDD.n1144 4.5005
R87700 VDD.n1309 VDD.n1144 4.5005
R87701 VDD.n1382 VDD.n1144 4.5005
R87702 VDD.n1307 VDD.n1144 4.5005
R87703 VDD.n1383 VDD.n1144 4.5005
R87704 VDD.n1306 VDD.n1144 4.5005
R87705 VDD.n1384 VDD.n1144 4.5005
R87706 VDD.n1304 VDD.n1144 4.5005
R87707 VDD.n1385 VDD.n1144 4.5005
R87708 VDD.n1303 VDD.n1144 4.5005
R87709 VDD.n1386 VDD.n1144 4.5005
R87710 VDD.n1301 VDD.n1144 4.5005
R87711 VDD.n1387 VDD.n1144 4.5005
R87712 VDD.n1300 VDD.n1144 4.5005
R87713 VDD.n1388 VDD.n1144 4.5005
R87714 VDD.n1298 VDD.n1144 4.5005
R87715 VDD.n1389 VDD.n1144 4.5005
R87716 VDD.n1297 VDD.n1144 4.5005
R87717 VDD.n1390 VDD.n1144 4.5005
R87718 VDD.n1295 VDD.n1144 4.5005
R87719 VDD.n1391 VDD.n1144 4.5005
R87720 VDD.n1294 VDD.n1144 4.5005
R87721 VDD.n1392 VDD.n1144 4.5005
R87722 VDD.n1292 VDD.n1144 4.5005
R87723 VDD.n1393 VDD.n1144 4.5005
R87724 VDD.n1291 VDD.n1144 4.5005
R87725 VDD.n1394 VDD.n1144 4.5005
R87726 VDD.n1289 VDD.n1144 4.5005
R87727 VDD.n1395 VDD.n1144 4.5005
R87728 VDD.n1288 VDD.n1144 4.5005
R87729 VDD.n1396 VDD.n1144 4.5005
R87730 VDD.n1286 VDD.n1144 4.5005
R87731 VDD.n1397 VDD.n1144 4.5005
R87732 VDD.n1285 VDD.n1144 4.5005
R87733 VDD.n1398 VDD.n1144 4.5005
R87734 VDD.n1283 VDD.n1144 4.5005
R87735 VDD.n1399 VDD.n1144 4.5005
R87736 VDD.n1282 VDD.n1144 4.5005
R87737 VDD.n1400 VDD.n1144 4.5005
R87738 VDD.n1280 VDD.n1144 4.5005
R87739 VDD.n1401 VDD.n1144 4.5005
R87740 VDD.n1279 VDD.n1144 4.5005
R87741 VDD.n1402 VDD.n1144 4.5005
R87742 VDD.n1277 VDD.n1144 4.5005
R87743 VDD.n1403 VDD.n1144 4.5005
R87744 VDD.n1276 VDD.n1144 4.5005
R87745 VDD.n1404 VDD.n1144 4.5005
R87746 VDD.n1274 VDD.n1144 4.5005
R87747 VDD.n1405 VDD.n1144 4.5005
R87748 VDD.n1273 VDD.n1144 4.5005
R87749 VDD.n1406 VDD.n1144 4.5005
R87750 VDD.n1271 VDD.n1144 4.5005
R87751 VDD.n1407 VDD.n1144 4.5005
R87752 VDD.n1270 VDD.n1144 4.5005
R87753 VDD.n1408 VDD.n1144 4.5005
R87754 VDD.n1268 VDD.n1144 4.5005
R87755 VDD.n1409 VDD.n1144 4.5005
R87756 VDD.n1267 VDD.n1144 4.5005
R87757 VDD.n1410 VDD.n1144 4.5005
R87758 VDD.n1265 VDD.n1144 4.5005
R87759 VDD.n1411 VDD.n1144 4.5005
R87760 VDD.n1264 VDD.n1144 4.5005
R87761 VDD.n1412 VDD.n1144 4.5005
R87762 VDD.n1262 VDD.n1144 4.5005
R87763 VDD.n1413 VDD.n1144 4.5005
R87764 VDD.n1261 VDD.n1144 4.5005
R87765 VDD.n1414 VDD.n1144 4.5005
R87766 VDD.n1415 VDD.n1144 4.5005
R87767 VDD.n1674 VDD.n1144 4.5005
R87768 VDD.n1676 VDD.n1246 4.5005
R87769 VDD.n1341 VDD.n1246 4.5005
R87770 VDD.n1342 VDD.n1246 4.5005
R87771 VDD.n1340 VDD.n1246 4.5005
R87772 VDD.n1344 VDD.n1246 4.5005
R87773 VDD.n1339 VDD.n1246 4.5005
R87774 VDD.n1345 VDD.n1246 4.5005
R87775 VDD.n1338 VDD.n1246 4.5005
R87776 VDD.n1347 VDD.n1246 4.5005
R87777 VDD.n1337 VDD.n1246 4.5005
R87778 VDD.n1348 VDD.n1246 4.5005
R87779 VDD.n1336 VDD.n1246 4.5005
R87780 VDD.n1350 VDD.n1246 4.5005
R87781 VDD.n1335 VDD.n1246 4.5005
R87782 VDD.n1351 VDD.n1246 4.5005
R87783 VDD.n1334 VDD.n1246 4.5005
R87784 VDD.n1353 VDD.n1246 4.5005
R87785 VDD.n1333 VDD.n1246 4.5005
R87786 VDD.n1354 VDD.n1246 4.5005
R87787 VDD.n1332 VDD.n1246 4.5005
R87788 VDD.n1356 VDD.n1246 4.5005
R87789 VDD.n1331 VDD.n1246 4.5005
R87790 VDD.n1357 VDD.n1246 4.5005
R87791 VDD.n1330 VDD.n1246 4.5005
R87792 VDD.n1359 VDD.n1246 4.5005
R87793 VDD.n1329 VDD.n1246 4.5005
R87794 VDD.n1360 VDD.n1246 4.5005
R87795 VDD.n1328 VDD.n1246 4.5005
R87796 VDD.n1362 VDD.n1246 4.5005
R87797 VDD.n1327 VDD.n1246 4.5005
R87798 VDD.n1363 VDD.n1246 4.5005
R87799 VDD.n1326 VDD.n1246 4.5005
R87800 VDD.n1365 VDD.n1246 4.5005
R87801 VDD.n1325 VDD.n1246 4.5005
R87802 VDD.n1366 VDD.n1246 4.5005
R87803 VDD.n1324 VDD.n1246 4.5005
R87804 VDD.n1368 VDD.n1246 4.5005
R87805 VDD.n1323 VDD.n1246 4.5005
R87806 VDD.n1369 VDD.n1246 4.5005
R87807 VDD.n1322 VDD.n1246 4.5005
R87808 VDD.n1371 VDD.n1246 4.5005
R87809 VDD.n1321 VDD.n1246 4.5005
R87810 VDD.n1372 VDD.n1246 4.5005
R87811 VDD.n1320 VDD.n1246 4.5005
R87812 VDD.n1374 VDD.n1246 4.5005
R87813 VDD.n1319 VDD.n1246 4.5005
R87814 VDD.n1375 VDD.n1246 4.5005
R87815 VDD.n1318 VDD.n1246 4.5005
R87816 VDD.n1376 VDD.n1246 4.5005
R87817 VDD.n1316 VDD.n1246 4.5005
R87818 VDD.n1377 VDD.n1246 4.5005
R87819 VDD.n1315 VDD.n1246 4.5005
R87820 VDD.n1378 VDD.n1246 4.5005
R87821 VDD.n1313 VDD.n1246 4.5005
R87822 VDD.n1379 VDD.n1246 4.5005
R87823 VDD.n1312 VDD.n1246 4.5005
R87824 VDD.n1380 VDD.n1246 4.5005
R87825 VDD.n1310 VDD.n1246 4.5005
R87826 VDD.n1381 VDD.n1246 4.5005
R87827 VDD.n1309 VDD.n1246 4.5005
R87828 VDD.n1382 VDD.n1246 4.5005
R87829 VDD.n1307 VDD.n1246 4.5005
R87830 VDD.n1383 VDD.n1246 4.5005
R87831 VDD.n1306 VDD.n1246 4.5005
R87832 VDD.n1384 VDD.n1246 4.5005
R87833 VDD.n1304 VDD.n1246 4.5005
R87834 VDD.n1385 VDD.n1246 4.5005
R87835 VDD.n1303 VDD.n1246 4.5005
R87836 VDD.n1386 VDD.n1246 4.5005
R87837 VDD.n1301 VDD.n1246 4.5005
R87838 VDD.n1387 VDD.n1246 4.5005
R87839 VDD.n1300 VDD.n1246 4.5005
R87840 VDD.n1388 VDD.n1246 4.5005
R87841 VDD.n1298 VDD.n1246 4.5005
R87842 VDD.n1389 VDD.n1246 4.5005
R87843 VDD.n1297 VDD.n1246 4.5005
R87844 VDD.n1390 VDD.n1246 4.5005
R87845 VDD.n1295 VDD.n1246 4.5005
R87846 VDD.n1391 VDD.n1246 4.5005
R87847 VDD.n1294 VDD.n1246 4.5005
R87848 VDD.n1392 VDD.n1246 4.5005
R87849 VDD.n1292 VDD.n1246 4.5005
R87850 VDD.n1393 VDD.n1246 4.5005
R87851 VDD.n1291 VDD.n1246 4.5005
R87852 VDD.n1394 VDD.n1246 4.5005
R87853 VDD.n1289 VDD.n1246 4.5005
R87854 VDD.n1395 VDD.n1246 4.5005
R87855 VDD.n1288 VDD.n1246 4.5005
R87856 VDD.n1396 VDD.n1246 4.5005
R87857 VDD.n1286 VDD.n1246 4.5005
R87858 VDD.n1397 VDD.n1246 4.5005
R87859 VDD.n1285 VDD.n1246 4.5005
R87860 VDD.n1398 VDD.n1246 4.5005
R87861 VDD.n1283 VDD.n1246 4.5005
R87862 VDD.n1399 VDD.n1246 4.5005
R87863 VDD.n1282 VDD.n1246 4.5005
R87864 VDD.n1400 VDD.n1246 4.5005
R87865 VDD.n1280 VDD.n1246 4.5005
R87866 VDD.n1401 VDD.n1246 4.5005
R87867 VDD.n1279 VDD.n1246 4.5005
R87868 VDD.n1402 VDD.n1246 4.5005
R87869 VDD.n1277 VDD.n1246 4.5005
R87870 VDD.n1403 VDD.n1246 4.5005
R87871 VDD.n1276 VDD.n1246 4.5005
R87872 VDD.n1404 VDD.n1246 4.5005
R87873 VDD.n1274 VDD.n1246 4.5005
R87874 VDD.n1405 VDD.n1246 4.5005
R87875 VDD.n1273 VDD.n1246 4.5005
R87876 VDD.n1406 VDD.n1246 4.5005
R87877 VDD.n1271 VDD.n1246 4.5005
R87878 VDD.n1407 VDD.n1246 4.5005
R87879 VDD.n1270 VDD.n1246 4.5005
R87880 VDD.n1408 VDD.n1246 4.5005
R87881 VDD.n1268 VDD.n1246 4.5005
R87882 VDD.n1409 VDD.n1246 4.5005
R87883 VDD.n1267 VDD.n1246 4.5005
R87884 VDD.n1410 VDD.n1246 4.5005
R87885 VDD.n1265 VDD.n1246 4.5005
R87886 VDD.n1411 VDD.n1246 4.5005
R87887 VDD.n1264 VDD.n1246 4.5005
R87888 VDD.n1412 VDD.n1246 4.5005
R87889 VDD.n1262 VDD.n1246 4.5005
R87890 VDD.n1413 VDD.n1246 4.5005
R87891 VDD.n1261 VDD.n1246 4.5005
R87892 VDD.n1414 VDD.n1246 4.5005
R87893 VDD.n1415 VDD.n1246 4.5005
R87894 VDD.n1674 VDD.n1246 4.5005
R87895 VDD.n1676 VDD.n1143 4.5005
R87896 VDD.n1341 VDD.n1143 4.5005
R87897 VDD.n1342 VDD.n1143 4.5005
R87898 VDD.n1340 VDD.n1143 4.5005
R87899 VDD.n1344 VDD.n1143 4.5005
R87900 VDD.n1339 VDD.n1143 4.5005
R87901 VDD.n1345 VDD.n1143 4.5005
R87902 VDD.n1338 VDD.n1143 4.5005
R87903 VDD.n1347 VDD.n1143 4.5005
R87904 VDD.n1337 VDD.n1143 4.5005
R87905 VDD.n1348 VDD.n1143 4.5005
R87906 VDD.n1336 VDD.n1143 4.5005
R87907 VDD.n1350 VDD.n1143 4.5005
R87908 VDD.n1335 VDD.n1143 4.5005
R87909 VDD.n1351 VDD.n1143 4.5005
R87910 VDD.n1334 VDD.n1143 4.5005
R87911 VDD.n1353 VDD.n1143 4.5005
R87912 VDD.n1333 VDD.n1143 4.5005
R87913 VDD.n1354 VDD.n1143 4.5005
R87914 VDD.n1332 VDD.n1143 4.5005
R87915 VDD.n1356 VDD.n1143 4.5005
R87916 VDD.n1331 VDD.n1143 4.5005
R87917 VDD.n1357 VDD.n1143 4.5005
R87918 VDD.n1330 VDD.n1143 4.5005
R87919 VDD.n1359 VDD.n1143 4.5005
R87920 VDD.n1329 VDD.n1143 4.5005
R87921 VDD.n1360 VDD.n1143 4.5005
R87922 VDD.n1328 VDD.n1143 4.5005
R87923 VDD.n1362 VDD.n1143 4.5005
R87924 VDD.n1327 VDD.n1143 4.5005
R87925 VDD.n1363 VDD.n1143 4.5005
R87926 VDD.n1326 VDD.n1143 4.5005
R87927 VDD.n1365 VDD.n1143 4.5005
R87928 VDD.n1325 VDD.n1143 4.5005
R87929 VDD.n1366 VDD.n1143 4.5005
R87930 VDD.n1324 VDD.n1143 4.5005
R87931 VDD.n1368 VDD.n1143 4.5005
R87932 VDD.n1323 VDD.n1143 4.5005
R87933 VDD.n1369 VDD.n1143 4.5005
R87934 VDD.n1322 VDD.n1143 4.5005
R87935 VDD.n1371 VDD.n1143 4.5005
R87936 VDD.n1321 VDD.n1143 4.5005
R87937 VDD.n1372 VDD.n1143 4.5005
R87938 VDD.n1320 VDD.n1143 4.5005
R87939 VDD.n1374 VDD.n1143 4.5005
R87940 VDD.n1319 VDD.n1143 4.5005
R87941 VDD.n1375 VDD.n1143 4.5005
R87942 VDD.n1318 VDD.n1143 4.5005
R87943 VDD.n1376 VDD.n1143 4.5005
R87944 VDD.n1316 VDD.n1143 4.5005
R87945 VDD.n1377 VDD.n1143 4.5005
R87946 VDD.n1315 VDD.n1143 4.5005
R87947 VDD.n1378 VDD.n1143 4.5005
R87948 VDD.n1313 VDD.n1143 4.5005
R87949 VDD.n1379 VDD.n1143 4.5005
R87950 VDD.n1312 VDD.n1143 4.5005
R87951 VDD.n1380 VDD.n1143 4.5005
R87952 VDD.n1310 VDD.n1143 4.5005
R87953 VDD.n1381 VDD.n1143 4.5005
R87954 VDD.n1309 VDD.n1143 4.5005
R87955 VDD.n1382 VDD.n1143 4.5005
R87956 VDD.n1307 VDD.n1143 4.5005
R87957 VDD.n1383 VDD.n1143 4.5005
R87958 VDD.n1306 VDD.n1143 4.5005
R87959 VDD.n1384 VDD.n1143 4.5005
R87960 VDD.n1304 VDD.n1143 4.5005
R87961 VDD.n1385 VDD.n1143 4.5005
R87962 VDD.n1303 VDD.n1143 4.5005
R87963 VDD.n1386 VDD.n1143 4.5005
R87964 VDD.n1301 VDD.n1143 4.5005
R87965 VDD.n1387 VDD.n1143 4.5005
R87966 VDD.n1300 VDD.n1143 4.5005
R87967 VDD.n1388 VDD.n1143 4.5005
R87968 VDD.n1298 VDD.n1143 4.5005
R87969 VDD.n1389 VDD.n1143 4.5005
R87970 VDD.n1297 VDD.n1143 4.5005
R87971 VDD.n1390 VDD.n1143 4.5005
R87972 VDD.n1295 VDD.n1143 4.5005
R87973 VDD.n1391 VDD.n1143 4.5005
R87974 VDD.n1294 VDD.n1143 4.5005
R87975 VDD.n1392 VDD.n1143 4.5005
R87976 VDD.n1292 VDD.n1143 4.5005
R87977 VDD.n1393 VDD.n1143 4.5005
R87978 VDD.n1291 VDD.n1143 4.5005
R87979 VDD.n1394 VDD.n1143 4.5005
R87980 VDD.n1289 VDD.n1143 4.5005
R87981 VDD.n1395 VDD.n1143 4.5005
R87982 VDD.n1288 VDD.n1143 4.5005
R87983 VDD.n1396 VDD.n1143 4.5005
R87984 VDD.n1286 VDD.n1143 4.5005
R87985 VDD.n1397 VDD.n1143 4.5005
R87986 VDD.n1285 VDD.n1143 4.5005
R87987 VDD.n1398 VDD.n1143 4.5005
R87988 VDD.n1283 VDD.n1143 4.5005
R87989 VDD.n1399 VDD.n1143 4.5005
R87990 VDD.n1282 VDD.n1143 4.5005
R87991 VDD.n1400 VDD.n1143 4.5005
R87992 VDD.n1280 VDD.n1143 4.5005
R87993 VDD.n1401 VDD.n1143 4.5005
R87994 VDD.n1279 VDD.n1143 4.5005
R87995 VDD.n1402 VDD.n1143 4.5005
R87996 VDD.n1277 VDD.n1143 4.5005
R87997 VDD.n1403 VDD.n1143 4.5005
R87998 VDD.n1276 VDD.n1143 4.5005
R87999 VDD.n1404 VDD.n1143 4.5005
R88000 VDD.n1274 VDD.n1143 4.5005
R88001 VDD.n1405 VDD.n1143 4.5005
R88002 VDD.n1273 VDD.n1143 4.5005
R88003 VDD.n1406 VDD.n1143 4.5005
R88004 VDD.n1271 VDD.n1143 4.5005
R88005 VDD.n1407 VDD.n1143 4.5005
R88006 VDD.n1270 VDD.n1143 4.5005
R88007 VDD.n1408 VDD.n1143 4.5005
R88008 VDD.n1268 VDD.n1143 4.5005
R88009 VDD.n1409 VDD.n1143 4.5005
R88010 VDD.n1267 VDD.n1143 4.5005
R88011 VDD.n1410 VDD.n1143 4.5005
R88012 VDD.n1265 VDD.n1143 4.5005
R88013 VDD.n1411 VDD.n1143 4.5005
R88014 VDD.n1264 VDD.n1143 4.5005
R88015 VDD.n1412 VDD.n1143 4.5005
R88016 VDD.n1262 VDD.n1143 4.5005
R88017 VDD.n1413 VDD.n1143 4.5005
R88018 VDD.n1261 VDD.n1143 4.5005
R88019 VDD.n1414 VDD.n1143 4.5005
R88020 VDD.n1415 VDD.n1143 4.5005
R88021 VDD.n1674 VDD.n1143 4.5005
R88022 VDD.n1676 VDD.n1247 4.5005
R88023 VDD.n1341 VDD.n1247 4.5005
R88024 VDD.n1342 VDD.n1247 4.5005
R88025 VDD.n1340 VDD.n1247 4.5005
R88026 VDD.n1344 VDD.n1247 4.5005
R88027 VDD.n1339 VDD.n1247 4.5005
R88028 VDD.n1345 VDD.n1247 4.5005
R88029 VDD.n1338 VDD.n1247 4.5005
R88030 VDD.n1347 VDD.n1247 4.5005
R88031 VDD.n1337 VDD.n1247 4.5005
R88032 VDD.n1348 VDD.n1247 4.5005
R88033 VDD.n1336 VDD.n1247 4.5005
R88034 VDD.n1350 VDD.n1247 4.5005
R88035 VDD.n1335 VDD.n1247 4.5005
R88036 VDD.n1351 VDD.n1247 4.5005
R88037 VDD.n1334 VDD.n1247 4.5005
R88038 VDD.n1353 VDD.n1247 4.5005
R88039 VDD.n1333 VDD.n1247 4.5005
R88040 VDD.n1354 VDD.n1247 4.5005
R88041 VDD.n1332 VDD.n1247 4.5005
R88042 VDD.n1356 VDD.n1247 4.5005
R88043 VDD.n1331 VDD.n1247 4.5005
R88044 VDD.n1357 VDD.n1247 4.5005
R88045 VDD.n1330 VDD.n1247 4.5005
R88046 VDD.n1359 VDD.n1247 4.5005
R88047 VDD.n1329 VDD.n1247 4.5005
R88048 VDD.n1360 VDD.n1247 4.5005
R88049 VDD.n1328 VDD.n1247 4.5005
R88050 VDD.n1362 VDD.n1247 4.5005
R88051 VDD.n1327 VDD.n1247 4.5005
R88052 VDD.n1363 VDD.n1247 4.5005
R88053 VDD.n1326 VDD.n1247 4.5005
R88054 VDD.n1365 VDD.n1247 4.5005
R88055 VDD.n1325 VDD.n1247 4.5005
R88056 VDD.n1366 VDD.n1247 4.5005
R88057 VDD.n1324 VDD.n1247 4.5005
R88058 VDD.n1368 VDD.n1247 4.5005
R88059 VDD.n1323 VDD.n1247 4.5005
R88060 VDD.n1369 VDD.n1247 4.5005
R88061 VDD.n1322 VDD.n1247 4.5005
R88062 VDD.n1371 VDD.n1247 4.5005
R88063 VDD.n1321 VDD.n1247 4.5005
R88064 VDD.n1372 VDD.n1247 4.5005
R88065 VDD.n1320 VDD.n1247 4.5005
R88066 VDD.n1374 VDD.n1247 4.5005
R88067 VDD.n1319 VDD.n1247 4.5005
R88068 VDD.n1375 VDD.n1247 4.5005
R88069 VDD.n1318 VDD.n1247 4.5005
R88070 VDD.n1376 VDD.n1247 4.5005
R88071 VDD.n1316 VDD.n1247 4.5005
R88072 VDD.n1377 VDD.n1247 4.5005
R88073 VDD.n1315 VDD.n1247 4.5005
R88074 VDD.n1378 VDD.n1247 4.5005
R88075 VDD.n1313 VDD.n1247 4.5005
R88076 VDD.n1379 VDD.n1247 4.5005
R88077 VDD.n1312 VDD.n1247 4.5005
R88078 VDD.n1380 VDD.n1247 4.5005
R88079 VDD.n1310 VDD.n1247 4.5005
R88080 VDD.n1381 VDD.n1247 4.5005
R88081 VDD.n1309 VDD.n1247 4.5005
R88082 VDD.n1382 VDD.n1247 4.5005
R88083 VDD.n1307 VDD.n1247 4.5005
R88084 VDD.n1383 VDD.n1247 4.5005
R88085 VDD.n1306 VDD.n1247 4.5005
R88086 VDD.n1384 VDD.n1247 4.5005
R88087 VDD.n1304 VDD.n1247 4.5005
R88088 VDD.n1385 VDD.n1247 4.5005
R88089 VDD.n1303 VDD.n1247 4.5005
R88090 VDD.n1386 VDD.n1247 4.5005
R88091 VDD.n1301 VDD.n1247 4.5005
R88092 VDD.n1387 VDD.n1247 4.5005
R88093 VDD.n1300 VDD.n1247 4.5005
R88094 VDD.n1388 VDD.n1247 4.5005
R88095 VDD.n1298 VDD.n1247 4.5005
R88096 VDD.n1389 VDD.n1247 4.5005
R88097 VDD.n1297 VDD.n1247 4.5005
R88098 VDD.n1390 VDD.n1247 4.5005
R88099 VDD.n1295 VDD.n1247 4.5005
R88100 VDD.n1391 VDD.n1247 4.5005
R88101 VDD.n1294 VDD.n1247 4.5005
R88102 VDD.n1392 VDD.n1247 4.5005
R88103 VDD.n1292 VDD.n1247 4.5005
R88104 VDD.n1393 VDD.n1247 4.5005
R88105 VDD.n1291 VDD.n1247 4.5005
R88106 VDD.n1394 VDD.n1247 4.5005
R88107 VDD.n1289 VDD.n1247 4.5005
R88108 VDD.n1395 VDD.n1247 4.5005
R88109 VDD.n1288 VDD.n1247 4.5005
R88110 VDD.n1396 VDD.n1247 4.5005
R88111 VDD.n1286 VDD.n1247 4.5005
R88112 VDD.n1397 VDD.n1247 4.5005
R88113 VDD.n1285 VDD.n1247 4.5005
R88114 VDD.n1398 VDD.n1247 4.5005
R88115 VDD.n1283 VDD.n1247 4.5005
R88116 VDD.n1399 VDD.n1247 4.5005
R88117 VDD.n1282 VDD.n1247 4.5005
R88118 VDD.n1400 VDD.n1247 4.5005
R88119 VDD.n1280 VDD.n1247 4.5005
R88120 VDD.n1401 VDD.n1247 4.5005
R88121 VDD.n1279 VDD.n1247 4.5005
R88122 VDD.n1402 VDD.n1247 4.5005
R88123 VDD.n1277 VDD.n1247 4.5005
R88124 VDD.n1403 VDD.n1247 4.5005
R88125 VDD.n1276 VDD.n1247 4.5005
R88126 VDD.n1404 VDD.n1247 4.5005
R88127 VDD.n1274 VDD.n1247 4.5005
R88128 VDD.n1405 VDD.n1247 4.5005
R88129 VDD.n1273 VDD.n1247 4.5005
R88130 VDD.n1406 VDD.n1247 4.5005
R88131 VDD.n1271 VDD.n1247 4.5005
R88132 VDD.n1407 VDD.n1247 4.5005
R88133 VDD.n1270 VDD.n1247 4.5005
R88134 VDD.n1408 VDD.n1247 4.5005
R88135 VDD.n1268 VDD.n1247 4.5005
R88136 VDD.n1409 VDD.n1247 4.5005
R88137 VDD.n1267 VDD.n1247 4.5005
R88138 VDD.n1410 VDD.n1247 4.5005
R88139 VDD.n1265 VDD.n1247 4.5005
R88140 VDD.n1411 VDD.n1247 4.5005
R88141 VDD.n1264 VDD.n1247 4.5005
R88142 VDD.n1412 VDD.n1247 4.5005
R88143 VDD.n1262 VDD.n1247 4.5005
R88144 VDD.n1413 VDD.n1247 4.5005
R88145 VDD.n1261 VDD.n1247 4.5005
R88146 VDD.n1414 VDD.n1247 4.5005
R88147 VDD.n1415 VDD.n1247 4.5005
R88148 VDD.n1674 VDD.n1247 4.5005
R88149 VDD.n1676 VDD.n1142 4.5005
R88150 VDD.n1341 VDD.n1142 4.5005
R88151 VDD.n1342 VDD.n1142 4.5005
R88152 VDD.n1340 VDD.n1142 4.5005
R88153 VDD.n1344 VDD.n1142 4.5005
R88154 VDD.n1339 VDD.n1142 4.5005
R88155 VDD.n1345 VDD.n1142 4.5005
R88156 VDD.n1338 VDD.n1142 4.5005
R88157 VDD.n1347 VDD.n1142 4.5005
R88158 VDD.n1337 VDD.n1142 4.5005
R88159 VDD.n1348 VDD.n1142 4.5005
R88160 VDD.n1336 VDD.n1142 4.5005
R88161 VDD.n1350 VDD.n1142 4.5005
R88162 VDD.n1335 VDD.n1142 4.5005
R88163 VDD.n1351 VDD.n1142 4.5005
R88164 VDD.n1334 VDD.n1142 4.5005
R88165 VDD.n1353 VDD.n1142 4.5005
R88166 VDD.n1333 VDD.n1142 4.5005
R88167 VDD.n1354 VDD.n1142 4.5005
R88168 VDD.n1332 VDD.n1142 4.5005
R88169 VDD.n1356 VDD.n1142 4.5005
R88170 VDD.n1331 VDD.n1142 4.5005
R88171 VDD.n1357 VDD.n1142 4.5005
R88172 VDD.n1330 VDD.n1142 4.5005
R88173 VDD.n1359 VDD.n1142 4.5005
R88174 VDD.n1329 VDD.n1142 4.5005
R88175 VDD.n1360 VDD.n1142 4.5005
R88176 VDD.n1328 VDD.n1142 4.5005
R88177 VDD.n1362 VDD.n1142 4.5005
R88178 VDD.n1327 VDD.n1142 4.5005
R88179 VDD.n1363 VDD.n1142 4.5005
R88180 VDD.n1326 VDD.n1142 4.5005
R88181 VDD.n1365 VDD.n1142 4.5005
R88182 VDD.n1325 VDD.n1142 4.5005
R88183 VDD.n1366 VDD.n1142 4.5005
R88184 VDD.n1324 VDD.n1142 4.5005
R88185 VDD.n1368 VDD.n1142 4.5005
R88186 VDD.n1323 VDD.n1142 4.5005
R88187 VDD.n1369 VDD.n1142 4.5005
R88188 VDD.n1322 VDD.n1142 4.5005
R88189 VDD.n1371 VDD.n1142 4.5005
R88190 VDD.n1321 VDD.n1142 4.5005
R88191 VDD.n1372 VDD.n1142 4.5005
R88192 VDD.n1320 VDD.n1142 4.5005
R88193 VDD.n1374 VDD.n1142 4.5005
R88194 VDD.n1319 VDD.n1142 4.5005
R88195 VDD.n1375 VDD.n1142 4.5005
R88196 VDD.n1318 VDD.n1142 4.5005
R88197 VDD.n1376 VDD.n1142 4.5005
R88198 VDD.n1316 VDD.n1142 4.5005
R88199 VDD.n1377 VDD.n1142 4.5005
R88200 VDD.n1315 VDD.n1142 4.5005
R88201 VDD.n1378 VDD.n1142 4.5005
R88202 VDD.n1313 VDD.n1142 4.5005
R88203 VDD.n1379 VDD.n1142 4.5005
R88204 VDD.n1312 VDD.n1142 4.5005
R88205 VDD.n1380 VDD.n1142 4.5005
R88206 VDD.n1310 VDD.n1142 4.5005
R88207 VDD.n1381 VDD.n1142 4.5005
R88208 VDD.n1309 VDD.n1142 4.5005
R88209 VDD.n1382 VDD.n1142 4.5005
R88210 VDD.n1307 VDD.n1142 4.5005
R88211 VDD.n1383 VDD.n1142 4.5005
R88212 VDD.n1306 VDD.n1142 4.5005
R88213 VDD.n1384 VDD.n1142 4.5005
R88214 VDD.n1304 VDD.n1142 4.5005
R88215 VDD.n1385 VDD.n1142 4.5005
R88216 VDD.n1303 VDD.n1142 4.5005
R88217 VDD.n1386 VDD.n1142 4.5005
R88218 VDD.n1301 VDD.n1142 4.5005
R88219 VDD.n1387 VDD.n1142 4.5005
R88220 VDD.n1300 VDD.n1142 4.5005
R88221 VDD.n1388 VDD.n1142 4.5005
R88222 VDD.n1298 VDD.n1142 4.5005
R88223 VDD.n1389 VDD.n1142 4.5005
R88224 VDD.n1297 VDD.n1142 4.5005
R88225 VDD.n1390 VDD.n1142 4.5005
R88226 VDD.n1295 VDD.n1142 4.5005
R88227 VDD.n1391 VDD.n1142 4.5005
R88228 VDD.n1294 VDD.n1142 4.5005
R88229 VDD.n1392 VDD.n1142 4.5005
R88230 VDD.n1292 VDD.n1142 4.5005
R88231 VDD.n1393 VDD.n1142 4.5005
R88232 VDD.n1291 VDD.n1142 4.5005
R88233 VDD.n1394 VDD.n1142 4.5005
R88234 VDD.n1289 VDD.n1142 4.5005
R88235 VDD.n1395 VDD.n1142 4.5005
R88236 VDD.n1288 VDD.n1142 4.5005
R88237 VDD.n1396 VDD.n1142 4.5005
R88238 VDD.n1286 VDD.n1142 4.5005
R88239 VDD.n1397 VDD.n1142 4.5005
R88240 VDD.n1285 VDD.n1142 4.5005
R88241 VDD.n1398 VDD.n1142 4.5005
R88242 VDD.n1283 VDD.n1142 4.5005
R88243 VDD.n1399 VDD.n1142 4.5005
R88244 VDD.n1282 VDD.n1142 4.5005
R88245 VDD.n1400 VDD.n1142 4.5005
R88246 VDD.n1280 VDD.n1142 4.5005
R88247 VDD.n1401 VDD.n1142 4.5005
R88248 VDD.n1279 VDD.n1142 4.5005
R88249 VDD.n1402 VDD.n1142 4.5005
R88250 VDD.n1277 VDD.n1142 4.5005
R88251 VDD.n1403 VDD.n1142 4.5005
R88252 VDD.n1276 VDD.n1142 4.5005
R88253 VDD.n1404 VDD.n1142 4.5005
R88254 VDD.n1274 VDD.n1142 4.5005
R88255 VDD.n1405 VDD.n1142 4.5005
R88256 VDD.n1273 VDD.n1142 4.5005
R88257 VDD.n1406 VDD.n1142 4.5005
R88258 VDD.n1271 VDD.n1142 4.5005
R88259 VDD.n1407 VDD.n1142 4.5005
R88260 VDD.n1270 VDD.n1142 4.5005
R88261 VDD.n1408 VDD.n1142 4.5005
R88262 VDD.n1268 VDD.n1142 4.5005
R88263 VDD.n1409 VDD.n1142 4.5005
R88264 VDD.n1267 VDD.n1142 4.5005
R88265 VDD.n1410 VDD.n1142 4.5005
R88266 VDD.n1265 VDD.n1142 4.5005
R88267 VDD.n1411 VDD.n1142 4.5005
R88268 VDD.n1264 VDD.n1142 4.5005
R88269 VDD.n1412 VDD.n1142 4.5005
R88270 VDD.n1262 VDD.n1142 4.5005
R88271 VDD.n1413 VDD.n1142 4.5005
R88272 VDD.n1261 VDD.n1142 4.5005
R88273 VDD.n1414 VDD.n1142 4.5005
R88274 VDD.n1415 VDD.n1142 4.5005
R88275 VDD.n1674 VDD.n1142 4.5005
R88276 VDD.n1676 VDD.n1248 4.5005
R88277 VDD.n1341 VDD.n1248 4.5005
R88278 VDD.n1342 VDD.n1248 4.5005
R88279 VDD.n1340 VDD.n1248 4.5005
R88280 VDD.n1344 VDD.n1248 4.5005
R88281 VDD.n1339 VDD.n1248 4.5005
R88282 VDD.n1345 VDD.n1248 4.5005
R88283 VDD.n1338 VDD.n1248 4.5005
R88284 VDD.n1347 VDD.n1248 4.5005
R88285 VDD.n1337 VDD.n1248 4.5005
R88286 VDD.n1348 VDD.n1248 4.5005
R88287 VDD.n1336 VDD.n1248 4.5005
R88288 VDD.n1350 VDD.n1248 4.5005
R88289 VDD.n1335 VDD.n1248 4.5005
R88290 VDD.n1351 VDD.n1248 4.5005
R88291 VDD.n1334 VDD.n1248 4.5005
R88292 VDD.n1353 VDD.n1248 4.5005
R88293 VDD.n1333 VDD.n1248 4.5005
R88294 VDD.n1354 VDD.n1248 4.5005
R88295 VDD.n1332 VDD.n1248 4.5005
R88296 VDD.n1356 VDD.n1248 4.5005
R88297 VDD.n1331 VDD.n1248 4.5005
R88298 VDD.n1357 VDD.n1248 4.5005
R88299 VDD.n1330 VDD.n1248 4.5005
R88300 VDD.n1359 VDD.n1248 4.5005
R88301 VDD.n1329 VDD.n1248 4.5005
R88302 VDD.n1360 VDD.n1248 4.5005
R88303 VDD.n1328 VDD.n1248 4.5005
R88304 VDD.n1362 VDD.n1248 4.5005
R88305 VDD.n1327 VDD.n1248 4.5005
R88306 VDD.n1363 VDD.n1248 4.5005
R88307 VDD.n1326 VDD.n1248 4.5005
R88308 VDD.n1365 VDD.n1248 4.5005
R88309 VDD.n1325 VDD.n1248 4.5005
R88310 VDD.n1366 VDD.n1248 4.5005
R88311 VDD.n1324 VDD.n1248 4.5005
R88312 VDD.n1368 VDD.n1248 4.5005
R88313 VDD.n1323 VDD.n1248 4.5005
R88314 VDD.n1369 VDD.n1248 4.5005
R88315 VDD.n1322 VDD.n1248 4.5005
R88316 VDD.n1371 VDD.n1248 4.5005
R88317 VDD.n1321 VDD.n1248 4.5005
R88318 VDD.n1372 VDD.n1248 4.5005
R88319 VDD.n1320 VDD.n1248 4.5005
R88320 VDD.n1374 VDD.n1248 4.5005
R88321 VDD.n1319 VDD.n1248 4.5005
R88322 VDD.n1375 VDD.n1248 4.5005
R88323 VDD.n1318 VDD.n1248 4.5005
R88324 VDD.n1376 VDD.n1248 4.5005
R88325 VDD.n1316 VDD.n1248 4.5005
R88326 VDD.n1377 VDD.n1248 4.5005
R88327 VDD.n1315 VDD.n1248 4.5005
R88328 VDD.n1378 VDD.n1248 4.5005
R88329 VDD.n1313 VDD.n1248 4.5005
R88330 VDD.n1379 VDD.n1248 4.5005
R88331 VDD.n1312 VDD.n1248 4.5005
R88332 VDD.n1380 VDD.n1248 4.5005
R88333 VDD.n1310 VDD.n1248 4.5005
R88334 VDD.n1381 VDD.n1248 4.5005
R88335 VDD.n1309 VDD.n1248 4.5005
R88336 VDD.n1382 VDD.n1248 4.5005
R88337 VDD.n1307 VDD.n1248 4.5005
R88338 VDD.n1383 VDD.n1248 4.5005
R88339 VDD.n1306 VDD.n1248 4.5005
R88340 VDD.n1384 VDD.n1248 4.5005
R88341 VDD.n1304 VDD.n1248 4.5005
R88342 VDD.n1385 VDD.n1248 4.5005
R88343 VDD.n1303 VDD.n1248 4.5005
R88344 VDD.n1386 VDD.n1248 4.5005
R88345 VDD.n1301 VDD.n1248 4.5005
R88346 VDD.n1387 VDD.n1248 4.5005
R88347 VDD.n1300 VDD.n1248 4.5005
R88348 VDD.n1388 VDD.n1248 4.5005
R88349 VDD.n1298 VDD.n1248 4.5005
R88350 VDD.n1389 VDD.n1248 4.5005
R88351 VDD.n1297 VDD.n1248 4.5005
R88352 VDD.n1390 VDD.n1248 4.5005
R88353 VDD.n1295 VDD.n1248 4.5005
R88354 VDD.n1391 VDD.n1248 4.5005
R88355 VDD.n1294 VDD.n1248 4.5005
R88356 VDD.n1392 VDD.n1248 4.5005
R88357 VDD.n1292 VDD.n1248 4.5005
R88358 VDD.n1393 VDD.n1248 4.5005
R88359 VDD.n1291 VDD.n1248 4.5005
R88360 VDD.n1394 VDD.n1248 4.5005
R88361 VDD.n1289 VDD.n1248 4.5005
R88362 VDD.n1395 VDD.n1248 4.5005
R88363 VDD.n1288 VDD.n1248 4.5005
R88364 VDD.n1396 VDD.n1248 4.5005
R88365 VDD.n1286 VDD.n1248 4.5005
R88366 VDD.n1397 VDD.n1248 4.5005
R88367 VDD.n1285 VDD.n1248 4.5005
R88368 VDD.n1398 VDD.n1248 4.5005
R88369 VDD.n1283 VDD.n1248 4.5005
R88370 VDD.n1399 VDD.n1248 4.5005
R88371 VDD.n1282 VDD.n1248 4.5005
R88372 VDD.n1400 VDD.n1248 4.5005
R88373 VDD.n1280 VDD.n1248 4.5005
R88374 VDD.n1401 VDD.n1248 4.5005
R88375 VDD.n1279 VDD.n1248 4.5005
R88376 VDD.n1402 VDD.n1248 4.5005
R88377 VDD.n1277 VDD.n1248 4.5005
R88378 VDD.n1403 VDD.n1248 4.5005
R88379 VDD.n1276 VDD.n1248 4.5005
R88380 VDD.n1404 VDD.n1248 4.5005
R88381 VDD.n1274 VDD.n1248 4.5005
R88382 VDD.n1405 VDD.n1248 4.5005
R88383 VDD.n1273 VDD.n1248 4.5005
R88384 VDD.n1406 VDD.n1248 4.5005
R88385 VDD.n1271 VDD.n1248 4.5005
R88386 VDD.n1407 VDD.n1248 4.5005
R88387 VDD.n1270 VDD.n1248 4.5005
R88388 VDD.n1408 VDD.n1248 4.5005
R88389 VDD.n1268 VDD.n1248 4.5005
R88390 VDD.n1409 VDD.n1248 4.5005
R88391 VDD.n1267 VDD.n1248 4.5005
R88392 VDD.n1410 VDD.n1248 4.5005
R88393 VDD.n1265 VDD.n1248 4.5005
R88394 VDD.n1411 VDD.n1248 4.5005
R88395 VDD.n1264 VDD.n1248 4.5005
R88396 VDD.n1412 VDD.n1248 4.5005
R88397 VDD.n1262 VDD.n1248 4.5005
R88398 VDD.n1413 VDD.n1248 4.5005
R88399 VDD.n1261 VDD.n1248 4.5005
R88400 VDD.n1414 VDD.n1248 4.5005
R88401 VDD.n1415 VDD.n1248 4.5005
R88402 VDD.n1674 VDD.n1248 4.5005
R88403 VDD.n1676 VDD.n1141 4.5005
R88404 VDD.n1341 VDD.n1141 4.5005
R88405 VDD.n1342 VDD.n1141 4.5005
R88406 VDD.n1340 VDD.n1141 4.5005
R88407 VDD.n1344 VDD.n1141 4.5005
R88408 VDD.n1339 VDD.n1141 4.5005
R88409 VDD.n1345 VDD.n1141 4.5005
R88410 VDD.n1338 VDD.n1141 4.5005
R88411 VDD.n1347 VDD.n1141 4.5005
R88412 VDD.n1337 VDD.n1141 4.5005
R88413 VDD.n1348 VDD.n1141 4.5005
R88414 VDD.n1336 VDD.n1141 4.5005
R88415 VDD.n1350 VDD.n1141 4.5005
R88416 VDD.n1335 VDD.n1141 4.5005
R88417 VDD.n1351 VDD.n1141 4.5005
R88418 VDD.n1334 VDD.n1141 4.5005
R88419 VDD.n1353 VDD.n1141 4.5005
R88420 VDD.n1333 VDD.n1141 4.5005
R88421 VDD.n1354 VDD.n1141 4.5005
R88422 VDD.n1332 VDD.n1141 4.5005
R88423 VDD.n1356 VDD.n1141 4.5005
R88424 VDD.n1331 VDD.n1141 4.5005
R88425 VDD.n1357 VDD.n1141 4.5005
R88426 VDD.n1330 VDD.n1141 4.5005
R88427 VDD.n1359 VDD.n1141 4.5005
R88428 VDD.n1329 VDD.n1141 4.5005
R88429 VDD.n1360 VDD.n1141 4.5005
R88430 VDD.n1328 VDD.n1141 4.5005
R88431 VDD.n1362 VDD.n1141 4.5005
R88432 VDD.n1327 VDD.n1141 4.5005
R88433 VDD.n1363 VDD.n1141 4.5005
R88434 VDD.n1326 VDD.n1141 4.5005
R88435 VDD.n1365 VDD.n1141 4.5005
R88436 VDD.n1325 VDD.n1141 4.5005
R88437 VDD.n1366 VDD.n1141 4.5005
R88438 VDD.n1324 VDD.n1141 4.5005
R88439 VDD.n1368 VDD.n1141 4.5005
R88440 VDD.n1323 VDD.n1141 4.5005
R88441 VDD.n1369 VDD.n1141 4.5005
R88442 VDD.n1322 VDD.n1141 4.5005
R88443 VDD.n1371 VDD.n1141 4.5005
R88444 VDD.n1321 VDD.n1141 4.5005
R88445 VDD.n1372 VDD.n1141 4.5005
R88446 VDD.n1320 VDD.n1141 4.5005
R88447 VDD.n1374 VDD.n1141 4.5005
R88448 VDD.n1319 VDD.n1141 4.5005
R88449 VDD.n1375 VDD.n1141 4.5005
R88450 VDD.n1318 VDD.n1141 4.5005
R88451 VDD.n1376 VDD.n1141 4.5005
R88452 VDD.n1316 VDD.n1141 4.5005
R88453 VDD.n1377 VDD.n1141 4.5005
R88454 VDD.n1315 VDD.n1141 4.5005
R88455 VDD.n1378 VDD.n1141 4.5005
R88456 VDD.n1313 VDD.n1141 4.5005
R88457 VDD.n1379 VDD.n1141 4.5005
R88458 VDD.n1312 VDD.n1141 4.5005
R88459 VDD.n1380 VDD.n1141 4.5005
R88460 VDD.n1310 VDD.n1141 4.5005
R88461 VDD.n1381 VDD.n1141 4.5005
R88462 VDD.n1309 VDD.n1141 4.5005
R88463 VDD.n1382 VDD.n1141 4.5005
R88464 VDD.n1307 VDD.n1141 4.5005
R88465 VDD.n1383 VDD.n1141 4.5005
R88466 VDD.n1306 VDD.n1141 4.5005
R88467 VDD.n1384 VDD.n1141 4.5005
R88468 VDD.n1304 VDD.n1141 4.5005
R88469 VDD.n1385 VDD.n1141 4.5005
R88470 VDD.n1303 VDD.n1141 4.5005
R88471 VDD.n1386 VDD.n1141 4.5005
R88472 VDD.n1301 VDD.n1141 4.5005
R88473 VDD.n1387 VDD.n1141 4.5005
R88474 VDD.n1300 VDD.n1141 4.5005
R88475 VDD.n1388 VDD.n1141 4.5005
R88476 VDD.n1298 VDD.n1141 4.5005
R88477 VDD.n1389 VDD.n1141 4.5005
R88478 VDD.n1297 VDD.n1141 4.5005
R88479 VDD.n1390 VDD.n1141 4.5005
R88480 VDD.n1295 VDD.n1141 4.5005
R88481 VDD.n1391 VDD.n1141 4.5005
R88482 VDD.n1294 VDD.n1141 4.5005
R88483 VDD.n1392 VDD.n1141 4.5005
R88484 VDD.n1292 VDD.n1141 4.5005
R88485 VDD.n1393 VDD.n1141 4.5005
R88486 VDD.n1291 VDD.n1141 4.5005
R88487 VDD.n1394 VDD.n1141 4.5005
R88488 VDD.n1289 VDD.n1141 4.5005
R88489 VDD.n1395 VDD.n1141 4.5005
R88490 VDD.n1288 VDD.n1141 4.5005
R88491 VDD.n1396 VDD.n1141 4.5005
R88492 VDD.n1286 VDD.n1141 4.5005
R88493 VDD.n1397 VDD.n1141 4.5005
R88494 VDD.n1285 VDD.n1141 4.5005
R88495 VDD.n1398 VDD.n1141 4.5005
R88496 VDD.n1283 VDD.n1141 4.5005
R88497 VDD.n1399 VDD.n1141 4.5005
R88498 VDD.n1282 VDD.n1141 4.5005
R88499 VDD.n1400 VDD.n1141 4.5005
R88500 VDD.n1280 VDD.n1141 4.5005
R88501 VDD.n1401 VDD.n1141 4.5005
R88502 VDD.n1279 VDD.n1141 4.5005
R88503 VDD.n1402 VDD.n1141 4.5005
R88504 VDD.n1277 VDD.n1141 4.5005
R88505 VDD.n1403 VDD.n1141 4.5005
R88506 VDD.n1276 VDD.n1141 4.5005
R88507 VDD.n1404 VDD.n1141 4.5005
R88508 VDD.n1274 VDD.n1141 4.5005
R88509 VDD.n1405 VDD.n1141 4.5005
R88510 VDD.n1273 VDD.n1141 4.5005
R88511 VDD.n1406 VDD.n1141 4.5005
R88512 VDD.n1271 VDD.n1141 4.5005
R88513 VDD.n1407 VDD.n1141 4.5005
R88514 VDD.n1270 VDD.n1141 4.5005
R88515 VDD.n1408 VDD.n1141 4.5005
R88516 VDD.n1268 VDD.n1141 4.5005
R88517 VDD.n1409 VDD.n1141 4.5005
R88518 VDD.n1267 VDD.n1141 4.5005
R88519 VDD.n1410 VDD.n1141 4.5005
R88520 VDD.n1265 VDD.n1141 4.5005
R88521 VDD.n1411 VDD.n1141 4.5005
R88522 VDD.n1264 VDD.n1141 4.5005
R88523 VDD.n1412 VDD.n1141 4.5005
R88524 VDD.n1262 VDD.n1141 4.5005
R88525 VDD.n1413 VDD.n1141 4.5005
R88526 VDD.n1261 VDD.n1141 4.5005
R88527 VDD.n1414 VDD.n1141 4.5005
R88528 VDD.n1415 VDD.n1141 4.5005
R88529 VDD.n1674 VDD.n1141 4.5005
R88530 VDD.n1676 VDD.n1249 4.5005
R88531 VDD.n1341 VDD.n1249 4.5005
R88532 VDD.n1342 VDD.n1249 4.5005
R88533 VDD.n1340 VDD.n1249 4.5005
R88534 VDD.n1344 VDD.n1249 4.5005
R88535 VDD.n1339 VDD.n1249 4.5005
R88536 VDD.n1345 VDD.n1249 4.5005
R88537 VDD.n1338 VDD.n1249 4.5005
R88538 VDD.n1347 VDD.n1249 4.5005
R88539 VDD.n1337 VDD.n1249 4.5005
R88540 VDD.n1348 VDD.n1249 4.5005
R88541 VDD.n1336 VDD.n1249 4.5005
R88542 VDD.n1350 VDD.n1249 4.5005
R88543 VDD.n1335 VDD.n1249 4.5005
R88544 VDD.n1351 VDD.n1249 4.5005
R88545 VDD.n1334 VDD.n1249 4.5005
R88546 VDD.n1353 VDD.n1249 4.5005
R88547 VDD.n1333 VDD.n1249 4.5005
R88548 VDD.n1354 VDD.n1249 4.5005
R88549 VDD.n1332 VDD.n1249 4.5005
R88550 VDD.n1356 VDD.n1249 4.5005
R88551 VDD.n1331 VDD.n1249 4.5005
R88552 VDD.n1357 VDD.n1249 4.5005
R88553 VDD.n1330 VDD.n1249 4.5005
R88554 VDD.n1359 VDD.n1249 4.5005
R88555 VDD.n1329 VDD.n1249 4.5005
R88556 VDD.n1360 VDD.n1249 4.5005
R88557 VDD.n1328 VDD.n1249 4.5005
R88558 VDD.n1362 VDD.n1249 4.5005
R88559 VDD.n1327 VDD.n1249 4.5005
R88560 VDD.n1363 VDD.n1249 4.5005
R88561 VDD.n1326 VDD.n1249 4.5005
R88562 VDD.n1365 VDD.n1249 4.5005
R88563 VDD.n1325 VDD.n1249 4.5005
R88564 VDD.n1366 VDD.n1249 4.5005
R88565 VDD.n1324 VDD.n1249 4.5005
R88566 VDD.n1368 VDD.n1249 4.5005
R88567 VDD.n1323 VDD.n1249 4.5005
R88568 VDD.n1369 VDD.n1249 4.5005
R88569 VDD.n1322 VDD.n1249 4.5005
R88570 VDD.n1371 VDD.n1249 4.5005
R88571 VDD.n1321 VDD.n1249 4.5005
R88572 VDD.n1372 VDD.n1249 4.5005
R88573 VDD.n1320 VDD.n1249 4.5005
R88574 VDD.n1374 VDD.n1249 4.5005
R88575 VDD.n1319 VDD.n1249 4.5005
R88576 VDD.n1375 VDD.n1249 4.5005
R88577 VDD.n1318 VDD.n1249 4.5005
R88578 VDD.n1376 VDD.n1249 4.5005
R88579 VDD.n1316 VDD.n1249 4.5005
R88580 VDD.n1377 VDD.n1249 4.5005
R88581 VDD.n1315 VDD.n1249 4.5005
R88582 VDD.n1378 VDD.n1249 4.5005
R88583 VDD.n1313 VDD.n1249 4.5005
R88584 VDD.n1379 VDD.n1249 4.5005
R88585 VDD.n1312 VDD.n1249 4.5005
R88586 VDD.n1380 VDD.n1249 4.5005
R88587 VDD.n1310 VDD.n1249 4.5005
R88588 VDD.n1381 VDD.n1249 4.5005
R88589 VDD.n1309 VDD.n1249 4.5005
R88590 VDD.n1382 VDD.n1249 4.5005
R88591 VDD.n1307 VDD.n1249 4.5005
R88592 VDD.n1383 VDD.n1249 4.5005
R88593 VDD.n1306 VDD.n1249 4.5005
R88594 VDD.n1384 VDD.n1249 4.5005
R88595 VDD.n1304 VDD.n1249 4.5005
R88596 VDD.n1385 VDD.n1249 4.5005
R88597 VDD.n1303 VDD.n1249 4.5005
R88598 VDD.n1386 VDD.n1249 4.5005
R88599 VDD.n1301 VDD.n1249 4.5005
R88600 VDD.n1387 VDD.n1249 4.5005
R88601 VDD.n1300 VDD.n1249 4.5005
R88602 VDD.n1388 VDD.n1249 4.5005
R88603 VDD.n1298 VDD.n1249 4.5005
R88604 VDD.n1389 VDD.n1249 4.5005
R88605 VDD.n1297 VDD.n1249 4.5005
R88606 VDD.n1390 VDD.n1249 4.5005
R88607 VDD.n1295 VDD.n1249 4.5005
R88608 VDD.n1391 VDD.n1249 4.5005
R88609 VDD.n1294 VDD.n1249 4.5005
R88610 VDD.n1392 VDD.n1249 4.5005
R88611 VDD.n1292 VDD.n1249 4.5005
R88612 VDD.n1393 VDD.n1249 4.5005
R88613 VDD.n1291 VDD.n1249 4.5005
R88614 VDD.n1394 VDD.n1249 4.5005
R88615 VDD.n1289 VDD.n1249 4.5005
R88616 VDD.n1395 VDD.n1249 4.5005
R88617 VDD.n1288 VDD.n1249 4.5005
R88618 VDD.n1396 VDD.n1249 4.5005
R88619 VDD.n1286 VDD.n1249 4.5005
R88620 VDD.n1397 VDD.n1249 4.5005
R88621 VDD.n1285 VDD.n1249 4.5005
R88622 VDD.n1398 VDD.n1249 4.5005
R88623 VDD.n1283 VDD.n1249 4.5005
R88624 VDD.n1399 VDD.n1249 4.5005
R88625 VDD.n1282 VDD.n1249 4.5005
R88626 VDD.n1400 VDD.n1249 4.5005
R88627 VDD.n1280 VDD.n1249 4.5005
R88628 VDD.n1401 VDD.n1249 4.5005
R88629 VDD.n1279 VDD.n1249 4.5005
R88630 VDD.n1402 VDD.n1249 4.5005
R88631 VDD.n1277 VDD.n1249 4.5005
R88632 VDD.n1403 VDD.n1249 4.5005
R88633 VDD.n1276 VDD.n1249 4.5005
R88634 VDD.n1404 VDD.n1249 4.5005
R88635 VDD.n1274 VDD.n1249 4.5005
R88636 VDD.n1405 VDD.n1249 4.5005
R88637 VDD.n1273 VDD.n1249 4.5005
R88638 VDD.n1406 VDD.n1249 4.5005
R88639 VDD.n1271 VDD.n1249 4.5005
R88640 VDD.n1407 VDD.n1249 4.5005
R88641 VDD.n1270 VDD.n1249 4.5005
R88642 VDD.n1408 VDD.n1249 4.5005
R88643 VDD.n1268 VDD.n1249 4.5005
R88644 VDD.n1409 VDD.n1249 4.5005
R88645 VDD.n1267 VDD.n1249 4.5005
R88646 VDD.n1410 VDD.n1249 4.5005
R88647 VDD.n1265 VDD.n1249 4.5005
R88648 VDD.n1411 VDD.n1249 4.5005
R88649 VDD.n1264 VDD.n1249 4.5005
R88650 VDD.n1412 VDD.n1249 4.5005
R88651 VDD.n1262 VDD.n1249 4.5005
R88652 VDD.n1413 VDD.n1249 4.5005
R88653 VDD.n1261 VDD.n1249 4.5005
R88654 VDD.n1414 VDD.n1249 4.5005
R88655 VDD.n1415 VDD.n1249 4.5005
R88656 VDD.n1674 VDD.n1249 4.5005
R88657 VDD.n1676 VDD.n1140 4.5005
R88658 VDD.n1341 VDD.n1140 4.5005
R88659 VDD.n1342 VDD.n1140 4.5005
R88660 VDD.n1340 VDD.n1140 4.5005
R88661 VDD.n1344 VDD.n1140 4.5005
R88662 VDD.n1339 VDD.n1140 4.5005
R88663 VDD.n1345 VDD.n1140 4.5005
R88664 VDD.n1338 VDD.n1140 4.5005
R88665 VDD.n1347 VDD.n1140 4.5005
R88666 VDD.n1337 VDD.n1140 4.5005
R88667 VDD.n1348 VDD.n1140 4.5005
R88668 VDD.n1336 VDD.n1140 4.5005
R88669 VDD.n1350 VDD.n1140 4.5005
R88670 VDD.n1335 VDD.n1140 4.5005
R88671 VDD.n1351 VDD.n1140 4.5005
R88672 VDD.n1334 VDD.n1140 4.5005
R88673 VDD.n1353 VDD.n1140 4.5005
R88674 VDD.n1333 VDD.n1140 4.5005
R88675 VDD.n1354 VDD.n1140 4.5005
R88676 VDD.n1332 VDD.n1140 4.5005
R88677 VDD.n1356 VDD.n1140 4.5005
R88678 VDD.n1331 VDD.n1140 4.5005
R88679 VDD.n1357 VDD.n1140 4.5005
R88680 VDD.n1330 VDD.n1140 4.5005
R88681 VDD.n1359 VDD.n1140 4.5005
R88682 VDD.n1329 VDD.n1140 4.5005
R88683 VDD.n1360 VDD.n1140 4.5005
R88684 VDD.n1328 VDD.n1140 4.5005
R88685 VDD.n1362 VDD.n1140 4.5005
R88686 VDD.n1327 VDD.n1140 4.5005
R88687 VDD.n1363 VDD.n1140 4.5005
R88688 VDD.n1326 VDD.n1140 4.5005
R88689 VDD.n1365 VDD.n1140 4.5005
R88690 VDD.n1325 VDD.n1140 4.5005
R88691 VDD.n1366 VDD.n1140 4.5005
R88692 VDD.n1324 VDD.n1140 4.5005
R88693 VDD.n1368 VDD.n1140 4.5005
R88694 VDD.n1323 VDD.n1140 4.5005
R88695 VDD.n1369 VDD.n1140 4.5005
R88696 VDD.n1322 VDD.n1140 4.5005
R88697 VDD.n1371 VDD.n1140 4.5005
R88698 VDD.n1321 VDD.n1140 4.5005
R88699 VDD.n1372 VDD.n1140 4.5005
R88700 VDD.n1320 VDD.n1140 4.5005
R88701 VDD.n1374 VDD.n1140 4.5005
R88702 VDD.n1319 VDD.n1140 4.5005
R88703 VDD.n1375 VDD.n1140 4.5005
R88704 VDD.n1318 VDD.n1140 4.5005
R88705 VDD.n1376 VDD.n1140 4.5005
R88706 VDD.n1316 VDD.n1140 4.5005
R88707 VDD.n1377 VDD.n1140 4.5005
R88708 VDD.n1315 VDD.n1140 4.5005
R88709 VDD.n1378 VDD.n1140 4.5005
R88710 VDD.n1313 VDD.n1140 4.5005
R88711 VDD.n1379 VDD.n1140 4.5005
R88712 VDD.n1312 VDD.n1140 4.5005
R88713 VDD.n1380 VDD.n1140 4.5005
R88714 VDD.n1310 VDD.n1140 4.5005
R88715 VDD.n1381 VDD.n1140 4.5005
R88716 VDD.n1309 VDD.n1140 4.5005
R88717 VDD.n1382 VDD.n1140 4.5005
R88718 VDD.n1307 VDD.n1140 4.5005
R88719 VDD.n1383 VDD.n1140 4.5005
R88720 VDD.n1306 VDD.n1140 4.5005
R88721 VDD.n1384 VDD.n1140 4.5005
R88722 VDD.n1304 VDD.n1140 4.5005
R88723 VDD.n1385 VDD.n1140 4.5005
R88724 VDD.n1303 VDD.n1140 4.5005
R88725 VDD.n1386 VDD.n1140 4.5005
R88726 VDD.n1301 VDD.n1140 4.5005
R88727 VDD.n1387 VDD.n1140 4.5005
R88728 VDD.n1300 VDD.n1140 4.5005
R88729 VDD.n1388 VDD.n1140 4.5005
R88730 VDD.n1298 VDD.n1140 4.5005
R88731 VDD.n1389 VDD.n1140 4.5005
R88732 VDD.n1297 VDD.n1140 4.5005
R88733 VDD.n1390 VDD.n1140 4.5005
R88734 VDD.n1295 VDD.n1140 4.5005
R88735 VDD.n1391 VDD.n1140 4.5005
R88736 VDD.n1294 VDD.n1140 4.5005
R88737 VDD.n1392 VDD.n1140 4.5005
R88738 VDD.n1292 VDD.n1140 4.5005
R88739 VDD.n1393 VDD.n1140 4.5005
R88740 VDD.n1291 VDD.n1140 4.5005
R88741 VDD.n1394 VDD.n1140 4.5005
R88742 VDD.n1289 VDD.n1140 4.5005
R88743 VDD.n1395 VDD.n1140 4.5005
R88744 VDD.n1288 VDD.n1140 4.5005
R88745 VDD.n1396 VDD.n1140 4.5005
R88746 VDD.n1286 VDD.n1140 4.5005
R88747 VDD.n1397 VDD.n1140 4.5005
R88748 VDD.n1285 VDD.n1140 4.5005
R88749 VDD.n1398 VDD.n1140 4.5005
R88750 VDD.n1283 VDD.n1140 4.5005
R88751 VDD.n1399 VDD.n1140 4.5005
R88752 VDD.n1282 VDD.n1140 4.5005
R88753 VDD.n1400 VDD.n1140 4.5005
R88754 VDD.n1280 VDD.n1140 4.5005
R88755 VDD.n1401 VDD.n1140 4.5005
R88756 VDD.n1279 VDD.n1140 4.5005
R88757 VDD.n1402 VDD.n1140 4.5005
R88758 VDD.n1277 VDD.n1140 4.5005
R88759 VDD.n1403 VDD.n1140 4.5005
R88760 VDD.n1276 VDD.n1140 4.5005
R88761 VDD.n1404 VDD.n1140 4.5005
R88762 VDD.n1274 VDD.n1140 4.5005
R88763 VDD.n1405 VDD.n1140 4.5005
R88764 VDD.n1273 VDD.n1140 4.5005
R88765 VDD.n1406 VDD.n1140 4.5005
R88766 VDD.n1271 VDD.n1140 4.5005
R88767 VDD.n1407 VDD.n1140 4.5005
R88768 VDD.n1270 VDD.n1140 4.5005
R88769 VDD.n1408 VDD.n1140 4.5005
R88770 VDD.n1268 VDD.n1140 4.5005
R88771 VDD.n1409 VDD.n1140 4.5005
R88772 VDD.n1267 VDD.n1140 4.5005
R88773 VDD.n1410 VDD.n1140 4.5005
R88774 VDD.n1265 VDD.n1140 4.5005
R88775 VDD.n1411 VDD.n1140 4.5005
R88776 VDD.n1264 VDD.n1140 4.5005
R88777 VDD.n1412 VDD.n1140 4.5005
R88778 VDD.n1262 VDD.n1140 4.5005
R88779 VDD.n1413 VDD.n1140 4.5005
R88780 VDD.n1261 VDD.n1140 4.5005
R88781 VDD.n1414 VDD.n1140 4.5005
R88782 VDD.n1415 VDD.n1140 4.5005
R88783 VDD.n1674 VDD.n1140 4.5005
R88784 VDD.n1676 VDD.n1250 4.5005
R88785 VDD.n1341 VDD.n1250 4.5005
R88786 VDD.n1342 VDD.n1250 4.5005
R88787 VDD.n1340 VDD.n1250 4.5005
R88788 VDD.n1344 VDD.n1250 4.5005
R88789 VDD.n1339 VDD.n1250 4.5005
R88790 VDD.n1345 VDD.n1250 4.5005
R88791 VDD.n1338 VDD.n1250 4.5005
R88792 VDD.n1347 VDD.n1250 4.5005
R88793 VDD.n1337 VDD.n1250 4.5005
R88794 VDD.n1348 VDD.n1250 4.5005
R88795 VDD.n1336 VDD.n1250 4.5005
R88796 VDD.n1350 VDD.n1250 4.5005
R88797 VDD.n1335 VDD.n1250 4.5005
R88798 VDD.n1351 VDD.n1250 4.5005
R88799 VDD.n1334 VDD.n1250 4.5005
R88800 VDD.n1353 VDD.n1250 4.5005
R88801 VDD.n1333 VDD.n1250 4.5005
R88802 VDD.n1354 VDD.n1250 4.5005
R88803 VDD.n1332 VDD.n1250 4.5005
R88804 VDD.n1356 VDD.n1250 4.5005
R88805 VDD.n1331 VDD.n1250 4.5005
R88806 VDD.n1357 VDD.n1250 4.5005
R88807 VDD.n1330 VDD.n1250 4.5005
R88808 VDD.n1359 VDD.n1250 4.5005
R88809 VDD.n1329 VDD.n1250 4.5005
R88810 VDD.n1360 VDD.n1250 4.5005
R88811 VDD.n1328 VDD.n1250 4.5005
R88812 VDD.n1362 VDD.n1250 4.5005
R88813 VDD.n1327 VDD.n1250 4.5005
R88814 VDD.n1363 VDD.n1250 4.5005
R88815 VDD.n1326 VDD.n1250 4.5005
R88816 VDD.n1365 VDD.n1250 4.5005
R88817 VDD.n1325 VDD.n1250 4.5005
R88818 VDD.n1366 VDD.n1250 4.5005
R88819 VDD.n1324 VDD.n1250 4.5005
R88820 VDD.n1368 VDD.n1250 4.5005
R88821 VDD.n1323 VDD.n1250 4.5005
R88822 VDD.n1369 VDD.n1250 4.5005
R88823 VDD.n1322 VDD.n1250 4.5005
R88824 VDD.n1371 VDD.n1250 4.5005
R88825 VDD.n1321 VDD.n1250 4.5005
R88826 VDD.n1372 VDD.n1250 4.5005
R88827 VDD.n1320 VDD.n1250 4.5005
R88828 VDD.n1374 VDD.n1250 4.5005
R88829 VDD.n1319 VDD.n1250 4.5005
R88830 VDD.n1375 VDD.n1250 4.5005
R88831 VDD.n1318 VDD.n1250 4.5005
R88832 VDD.n1376 VDD.n1250 4.5005
R88833 VDD.n1316 VDD.n1250 4.5005
R88834 VDD.n1377 VDD.n1250 4.5005
R88835 VDD.n1315 VDD.n1250 4.5005
R88836 VDD.n1378 VDD.n1250 4.5005
R88837 VDD.n1313 VDD.n1250 4.5005
R88838 VDD.n1379 VDD.n1250 4.5005
R88839 VDD.n1312 VDD.n1250 4.5005
R88840 VDD.n1380 VDD.n1250 4.5005
R88841 VDD.n1310 VDD.n1250 4.5005
R88842 VDD.n1381 VDD.n1250 4.5005
R88843 VDD.n1309 VDD.n1250 4.5005
R88844 VDD.n1382 VDD.n1250 4.5005
R88845 VDD.n1307 VDD.n1250 4.5005
R88846 VDD.n1383 VDD.n1250 4.5005
R88847 VDD.n1306 VDD.n1250 4.5005
R88848 VDD.n1384 VDD.n1250 4.5005
R88849 VDD.n1304 VDD.n1250 4.5005
R88850 VDD.n1385 VDD.n1250 4.5005
R88851 VDD.n1303 VDD.n1250 4.5005
R88852 VDD.n1386 VDD.n1250 4.5005
R88853 VDD.n1301 VDD.n1250 4.5005
R88854 VDD.n1387 VDD.n1250 4.5005
R88855 VDD.n1300 VDD.n1250 4.5005
R88856 VDD.n1388 VDD.n1250 4.5005
R88857 VDD.n1298 VDD.n1250 4.5005
R88858 VDD.n1389 VDD.n1250 4.5005
R88859 VDD.n1297 VDD.n1250 4.5005
R88860 VDD.n1390 VDD.n1250 4.5005
R88861 VDD.n1295 VDD.n1250 4.5005
R88862 VDD.n1391 VDD.n1250 4.5005
R88863 VDD.n1294 VDD.n1250 4.5005
R88864 VDD.n1392 VDD.n1250 4.5005
R88865 VDD.n1292 VDD.n1250 4.5005
R88866 VDD.n1393 VDD.n1250 4.5005
R88867 VDD.n1291 VDD.n1250 4.5005
R88868 VDD.n1394 VDD.n1250 4.5005
R88869 VDD.n1289 VDD.n1250 4.5005
R88870 VDD.n1395 VDD.n1250 4.5005
R88871 VDD.n1288 VDD.n1250 4.5005
R88872 VDD.n1396 VDD.n1250 4.5005
R88873 VDD.n1286 VDD.n1250 4.5005
R88874 VDD.n1397 VDD.n1250 4.5005
R88875 VDD.n1285 VDD.n1250 4.5005
R88876 VDD.n1398 VDD.n1250 4.5005
R88877 VDD.n1283 VDD.n1250 4.5005
R88878 VDD.n1399 VDD.n1250 4.5005
R88879 VDD.n1282 VDD.n1250 4.5005
R88880 VDD.n1400 VDD.n1250 4.5005
R88881 VDD.n1280 VDD.n1250 4.5005
R88882 VDD.n1401 VDD.n1250 4.5005
R88883 VDD.n1279 VDD.n1250 4.5005
R88884 VDD.n1402 VDD.n1250 4.5005
R88885 VDD.n1277 VDD.n1250 4.5005
R88886 VDD.n1403 VDD.n1250 4.5005
R88887 VDD.n1276 VDD.n1250 4.5005
R88888 VDD.n1404 VDD.n1250 4.5005
R88889 VDD.n1274 VDD.n1250 4.5005
R88890 VDD.n1405 VDD.n1250 4.5005
R88891 VDD.n1273 VDD.n1250 4.5005
R88892 VDD.n1406 VDD.n1250 4.5005
R88893 VDD.n1271 VDD.n1250 4.5005
R88894 VDD.n1407 VDD.n1250 4.5005
R88895 VDD.n1270 VDD.n1250 4.5005
R88896 VDD.n1408 VDD.n1250 4.5005
R88897 VDD.n1268 VDD.n1250 4.5005
R88898 VDD.n1409 VDD.n1250 4.5005
R88899 VDD.n1267 VDD.n1250 4.5005
R88900 VDD.n1410 VDD.n1250 4.5005
R88901 VDD.n1265 VDD.n1250 4.5005
R88902 VDD.n1411 VDD.n1250 4.5005
R88903 VDD.n1264 VDD.n1250 4.5005
R88904 VDD.n1412 VDD.n1250 4.5005
R88905 VDD.n1262 VDD.n1250 4.5005
R88906 VDD.n1413 VDD.n1250 4.5005
R88907 VDD.n1261 VDD.n1250 4.5005
R88908 VDD.n1414 VDD.n1250 4.5005
R88909 VDD.n1415 VDD.n1250 4.5005
R88910 VDD.n1674 VDD.n1250 4.5005
R88911 VDD.n1676 VDD.n1139 4.5005
R88912 VDD.n1341 VDD.n1139 4.5005
R88913 VDD.n1342 VDD.n1139 4.5005
R88914 VDD.n1340 VDD.n1139 4.5005
R88915 VDD.n1344 VDD.n1139 4.5005
R88916 VDD.n1339 VDD.n1139 4.5005
R88917 VDD.n1345 VDD.n1139 4.5005
R88918 VDD.n1338 VDD.n1139 4.5005
R88919 VDD.n1347 VDD.n1139 4.5005
R88920 VDD.n1337 VDD.n1139 4.5005
R88921 VDD.n1348 VDD.n1139 4.5005
R88922 VDD.n1336 VDD.n1139 4.5005
R88923 VDD.n1350 VDD.n1139 4.5005
R88924 VDD.n1335 VDD.n1139 4.5005
R88925 VDD.n1351 VDD.n1139 4.5005
R88926 VDD.n1334 VDD.n1139 4.5005
R88927 VDD.n1353 VDD.n1139 4.5005
R88928 VDD.n1333 VDD.n1139 4.5005
R88929 VDD.n1354 VDD.n1139 4.5005
R88930 VDD.n1332 VDD.n1139 4.5005
R88931 VDD.n1356 VDD.n1139 4.5005
R88932 VDD.n1331 VDD.n1139 4.5005
R88933 VDD.n1357 VDD.n1139 4.5005
R88934 VDD.n1330 VDD.n1139 4.5005
R88935 VDD.n1359 VDD.n1139 4.5005
R88936 VDD.n1329 VDD.n1139 4.5005
R88937 VDD.n1360 VDD.n1139 4.5005
R88938 VDD.n1328 VDD.n1139 4.5005
R88939 VDD.n1362 VDD.n1139 4.5005
R88940 VDD.n1327 VDD.n1139 4.5005
R88941 VDD.n1363 VDD.n1139 4.5005
R88942 VDD.n1326 VDD.n1139 4.5005
R88943 VDD.n1365 VDD.n1139 4.5005
R88944 VDD.n1325 VDD.n1139 4.5005
R88945 VDD.n1366 VDD.n1139 4.5005
R88946 VDD.n1324 VDD.n1139 4.5005
R88947 VDD.n1368 VDD.n1139 4.5005
R88948 VDD.n1323 VDD.n1139 4.5005
R88949 VDD.n1369 VDD.n1139 4.5005
R88950 VDD.n1322 VDD.n1139 4.5005
R88951 VDD.n1371 VDD.n1139 4.5005
R88952 VDD.n1321 VDD.n1139 4.5005
R88953 VDD.n1372 VDD.n1139 4.5005
R88954 VDD.n1320 VDD.n1139 4.5005
R88955 VDD.n1374 VDD.n1139 4.5005
R88956 VDD.n1319 VDD.n1139 4.5005
R88957 VDD.n1375 VDD.n1139 4.5005
R88958 VDD.n1318 VDD.n1139 4.5005
R88959 VDD.n1376 VDD.n1139 4.5005
R88960 VDD.n1316 VDD.n1139 4.5005
R88961 VDD.n1377 VDD.n1139 4.5005
R88962 VDD.n1315 VDD.n1139 4.5005
R88963 VDD.n1378 VDD.n1139 4.5005
R88964 VDD.n1313 VDD.n1139 4.5005
R88965 VDD.n1379 VDD.n1139 4.5005
R88966 VDD.n1312 VDD.n1139 4.5005
R88967 VDD.n1380 VDD.n1139 4.5005
R88968 VDD.n1310 VDD.n1139 4.5005
R88969 VDD.n1381 VDD.n1139 4.5005
R88970 VDD.n1309 VDD.n1139 4.5005
R88971 VDD.n1382 VDD.n1139 4.5005
R88972 VDD.n1307 VDD.n1139 4.5005
R88973 VDD.n1383 VDD.n1139 4.5005
R88974 VDD.n1306 VDD.n1139 4.5005
R88975 VDD.n1384 VDD.n1139 4.5005
R88976 VDD.n1304 VDD.n1139 4.5005
R88977 VDD.n1385 VDD.n1139 4.5005
R88978 VDD.n1303 VDD.n1139 4.5005
R88979 VDD.n1386 VDD.n1139 4.5005
R88980 VDD.n1301 VDD.n1139 4.5005
R88981 VDD.n1387 VDD.n1139 4.5005
R88982 VDD.n1300 VDD.n1139 4.5005
R88983 VDD.n1388 VDD.n1139 4.5005
R88984 VDD.n1298 VDD.n1139 4.5005
R88985 VDD.n1389 VDD.n1139 4.5005
R88986 VDD.n1297 VDD.n1139 4.5005
R88987 VDD.n1390 VDD.n1139 4.5005
R88988 VDD.n1295 VDD.n1139 4.5005
R88989 VDD.n1391 VDD.n1139 4.5005
R88990 VDD.n1294 VDD.n1139 4.5005
R88991 VDD.n1392 VDD.n1139 4.5005
R88992 VDD.n1292 VDD.n1139 4.5005
R88993 VDD.n1393 VDD.n1139 4.5005
R88994 VDD.n1291 VDD.n1139 4.5005
R88995 VDD.n1394 VDD.n1139 4.5005
R88996 VDD.n1289 VDD.n1139 4.5005
R88997 VDD.n1395 VDD.n1139 4.5005
R88998 VDD.n1288 VDD.n1139 4.5005
R88999 VDD.n1396 VDD.n1139 4.5005
R89000 VDD.n1286 VDD.n1139 4.5005
R89001 VDD.n1397 VDD.n1139 4.5005
R89002 VDD.n1285 VDD.n1139 4.5005
R89003 VDD.n1398 VDD.n1139 4.5005
R89004 VDD.n1283 VDD.n1139 4.5005
R89005 VDD.n1399 VDD.n1139 4.5005
R89006 VDD.n1282 VDD.n1139 4.5005
R89007 VDD.n1400 VDD.n1139 4.5005
R89008 VDD.n1280 VDD.n1139 4.5005
R89009 VDD.n1401 VDD.n1139 4.5005
R89010 VDD.n1279 VDD.n1139 4.5005
R89011 VDD.n1402 VDD.n1139 4.5005
R89012 VDD.n1277 VDD.n1139 4.5005
R89013 VDD.n1403 VDD.n1139 4.5005
R89014 VDD.n1276 VDD.n1139 4.5005
R89015 VDD.n1404 VDD.n1139 4.5005
R89016 VDD.n1274 VDD.n1139 4.5005
R89017 VDD.n1405 VDD.n1139 4.5005
R89018 VDD.n1273 VDD.n1139 4.5005
R89019 VDD.n1406 VDD.n1139 4.5005
R89020 VDD.n1271 VDD.n1139 4.5005
R89021 VDD.n1407 VDD.n1139 4.5005
R89022 VDD.n1270 VDD.n1139 4.5005
R89023 VDD.n1408 VDD.n1139 4.5005
R89024 VDD.n1268 VDD.n1139 4.5005
R89025 VDD.n1409 VDD.n1139 4.5005
R89026 VDD.n1267 VDD.n1139 4.5005
R89027 VDD.n1410 VDD.n1139 4.5005
R89028 VDD.n1265 VDD.n1139 4.5005
R89029 VDD.n1411 VDD.n1139 4.5005
R89030 VDD.n1264 VDD.n1139 4.5005
R89031 VDD.n1412 VDD.n1139 4.5005
R89032 VDD.n1262 VDD.n1139 4.5005
R89033 VDD.n1413 VDD.n1139 4.5005
R89034 VDD.n1261 VDD.n1139 4.5005
R89035 VDD.n1414 VDD.n1139 4.5005
R89036 VDD.n1415 VDD.n1139 4.5005
R89037 VDD.n1674 VDD.n1139 4.5005
R89038 VDD.n1676 VDD.n1251 4.5005
R89039 VDD.n1341 VDD.n1251 4.5005
R89040 VDD.n1342 VDD.n1251 4.5005
R89041 VDD.n1340 VDD.n1251 4.5005
R89042 VDD.n1344 VDD.n1251 4.5005
R89043 VDD.n1339 VDD.n1251 4.5005
R89044 VDD.n1345 VDD.n1251 4.5005
R89045 VDD.n1338 VDD.n1251 4.5005
R89046 VDD.n1347 VDD.n1251 4.5005
R89047 VDD.n1337 VDD.n1251 4.5005
R89048 VDD.n1348 VDD.n1251 4.5005
R89049 VDD.n1336 VDD.n1251 4.5005
R89050 VDD.n1350 VDD.n1251 4.5005
R89051 VDD.n1335 VDD.n1251 4.5005
R89052 VDD.n1351 VDD.n1251 4.5005
R89053 VDD.n1334 VDD.n1251 4.5005
R89054 VDD.n1353 VDD.n1251 4.5005
R89055 VDD.n1333 VDD.n1251 4.5005
R89056 VDD.n1354 VDD.n1251 4.5005
R89057 VDD.n1332 VDD.n1251 4.5005
R89058 VDD.n1356 VDD.n1251 4.5005
R89059 VDD.n1331 VDD.n1251 4.5005
R89060 VDD.n1357 VDD.n1251 4.5005
R89061 VDD.n1330 VDD.n1251 4.5005
R89062 VDD.n1359 VDD.n1251 4.5005
R89063 VDD.n1329 VDD.n1251 4.5005
R89064 VDD.n1360 VDD.n1251 4.5005
R89065 VDD.n1328 VDD.n1251 4.5005
R89066 VDD.n1362 VDD.n1251 4.5005
R89067 VDD.n1327 VDD.n1251 4.5005
R89068 VDD.n1363 VDD.n1251 4.5005
R89069 VDD.n1326 VDD.n1251 4.5005
R89070 VDD.n1365 VDD.n1251 4.5005
R89071 VDD.n1325 VDD.n1251 4.5005
R89072 VDD.n1366 VDD.n1251 4.5005
R89073 VDD.n1324 VDD.n1251 4.5005
R89074 VDD.n1368 VDD.n1251 4.5005
R89075 VDD.n1323 VDD.n1251 4.5005
R89076 VDD.n1369 VDD.n1251 4.5005
R89077 VDD.n1322 VDD.n1251 4.5005
R89078 VDD.n1371 VDD.n1251 4.5005
R89079 VDD.n1321 VDD.n1251 4.5005
R89080 VDD.n1372 VDD.n1251 4.5005
R89081 VDD.n1320 VDD.n1251 4.5005
R89082 VDD.n1374 VDD.n1251 4.5005
R89083 VDD.n1319 VDD.n1251 4.5005
R89084 VDD.n1375 VDD.n1251 4.5005
R89085 VDD.n1318 VDD.n1251 4.5005
R89086 VDD.n1376 VDD.n1251 4.5005
R89087 VDD.n1316 VDD.n1251 4.5005
R89088 VDD.n1377 VDD.n1251 4.5005
R89089 VDD.n1315 VDD.n1251 4.5005
R89090 VDD.n1378 VDD.n1251 4.5005
R89091 VDD.n1313 VDD.n1251 4.5005
R89092 VDD.n1379 VDD.n1251 4.5005
R89093 VDD.n1312 VDD.n1251 4.5005
R89094 VDD.n1380 VDD.n1251 4.5005
R89095 VDD.n1310 VDD.n1251 4.5005
R89096 VDD.n1381 VDD.n1251 4.5005
R89097 VDD.n1309 VDD.n1251 4.5005
R89098 VDD.n1382 VDD.n1251 4.5005
R89099 VDD.n1307 VDD.n1251 4.5005
R89100 VDD.n1383 VDD.n1251 4.5005
R89101 VDD.n1306 VDD.n1251 4.5005
R89102 VDD.n1384 VDD.n1251 4.5005
R89103 VDD.n1304 VDD.n1251 4.5005
R89104 VDD.n1385 VDD.n1251 4.5005
R89105 VDD.n1303 VDD.n1251 4.5005
R89106 VDD.n1386 VDD.n1251 4.5005
R89107 VDD.n1301 VDD.n1251 4.5005
R89108 VDD.n1387 VDD.n1251 4.5005
R89109 VDD.n1300 VDD.n1251 4.5005
R89110 VDD.n1388 VDD.n1251 4.5005
R89111 VDD.n1298 VDD.n1251 4.5005
R89112 VDD.n1389 VDD.n1251 4.5005
R89113 VDD.n1297 VDD.n1251 4.5005
R89114 VDD.n1390 VDD.n1251 4.5005
R89115 VDD.n1295 VDD.n1251 4.5005
R89116 VDD.n1391 VDD.n1251 4.5005
R89117 VDD.n1294 VDD.n1251 4.5005
R89118 VDD.n1392 VDD.n1251 4.5005
R89119 VDD.n1292 VDD.n1251 4.5005
R89120 VDD.n1393 VDD.n1251 4.5005
R89121 VDD.n1291 VDD.n1251 4.5005
R89122 VDD.n1394 VDD.n1251 4.5005
R89123 VDD.n1289 VDD.n1251 4.5005
R89124 VDD.n1395 VDD.n1251 4.5005
R89125 VDD.n1288 VDD.n1251 4.5005
R89126 VDD.n1396 VDD.n1251 4.5005
R89127 VDD.n1286 VDD.n1251 4.5005
R89128 VDD.n1397 VDD.n1251 4.5005
R89129 VDD.n1285 VDD.n1251 4.5005
R89130 VDD.n1398 VDD.n1251 4.5005
R89131 VDD.n1283 VDD.n1251 4.5005
R89132 VDD.n1399 VDD.n1251 4.5005
R89133 VDD.n1282 VDD.n1251 4.5005
R89134 VDD.n1400 VDD.n1251 4.5005
R89135 VDD.n1280 VDD.n1251 4.5005
R89136 VDD.n1401 VDD.n1251 4.5005
R89137 VDD.n1279 VDD.n1251 4.5005
R89138 VDD.n1402 VDD.n1251 4.5005
R89139 VDD.n1277 VDD.n1251 4.5005
R89140 VDD.n1403 VDD.n1251 4.5005
R89141 VDD.n1276 VDD.n1251 4.5005
R89142 VDD.n1404 VDD.n1251 4.5005
R89143 VDD.n1274 VDD.n1251 4.5005
R89144 VDD.n1405 VDD.n1251 4.5005
R89145 VDD.n1273 VDD.n1251 4.5005
R89146 VDD.n1406 VDD.n1251 4.5005
R89147 VDD.n1271 VDD.n1251 4.5005
R89148 VDD.n1407 VDD.n1251 4.5005
R89149 VDD.n1270 VDD.n1251 4.5005
R89150 VDD.n1408 VDD.n1251 4.5005
R89151 VDD.n1268 VDD.n1251 4.5005
R89152 VDD.n1409 VDD.n1251 4.5005
R89153 VDD.n1267 VDD.n1251 4.5005
R89154 VDD.n1410 VDD.n1251 4.5005
R89155 VDD.n1265 VDD.n1251 4.5005
R89156 VDD.n1411 VDD.n1251 4.5005
R89157 VDD.n1264 VDD.n1251 4.5005
R89158 VDD.n1412 VDD.n1251 4.5005
R89159 VDD.n1262 VDD.n1251 4.5005
R89160 VDD.n1413 VDD.n1251 4.5005
R89161 VDD.n1261 VDD.n1251 4.5005
R89162 VDD.n1414 VDD.n1251 4.5005
R89163 VDD.n1415 VDD.n1251 4.5005
R89164 VDD.n1674 VDD.n1251 4.5005
R89165 VDD.n1676 VDD.n1138 4.5005
R89166 VDD.n1341 VDD.n1138 4.5005
R89167 VDD.n1342 VDD.n1138 4.5005
R89168 VDD.n1340 VDD.n1138 4.5005
R89169 VDD.n1344 VDD.n1138 4.5005
R89170 VDD.n1339 VDD.n1138 4.5005
R89171 VDD.n1345 VDD.n1138 4.5005
R89172 VDD.n1338 VDD.n1138 4.5005
R89173 VDD.n1347 VDD.n1138 4.5005
R89174 VDD.n1337 VDD.n1138 4.5005
R89175 VDD.n1348 VDD.n1138 4.5005
R89176 VDD.n1336 VDD.n1138 4.5005
R89177 VDD.n1350 VDD.n1138 4.5005
R89178 VDD.n1335 VDD.n1138 4.5005
R89179 VDD.n1351 VDD.n1138 4.5005
R89180 VDD.n1334 VDD.n1138 4.5005
R89181 VDD.n1353 VDD.n1138 4.5005
R89182 VDD.n1333 VDD.n1138 4.5005
R89183 VDD.n1354 VDD.n1138 4.5005
R89184 VDD.n1332 VDD.n1138 4.5005
R89185 VDD.n1356 VDD.n1138 4.5005
R89186 VDD.n1331 VDD.n1138 4.5005
R89187 VDD.n1357 VDD.n1138 4.5005
R89188 VDD.n1330 VDD.n1138 4.5005
R89189 VDD.n1359 VDD.n1138 4.5005
R89190 VDD.n1329 VDD.n1138 4.5005
R89191 VDD.n1360 VDD.n1138 4.5005
R89192 VDD.n1328 VDD.n1138 4.5005
R89193 VDD.n1362 VDD.n1138 4.5005
R89194 VDD.n1327 VDD.n1138 4.5005
R89195 VDD.n1363 VDD.n1138 4.5005
R89196 VDD.n1326 VDD.n1138 4.5005
R89197 VDD.n1365 VDD.n1138 4.5005
R89198 VDD.n1325 VDD.n1138 4.5005
R89199 VDD.n1366 VDD.n1138 4.5005
R89200 VDD.n1324 VDD.n1138 4.5005
R89201 VDD.n1368 VDD.n1138 4.5005
R89202 VDD.n1323 VDD.n1138 4.5005
R89203 VDD.n1369 VDD.n1138 4.5005
R89204 VDD.n1322 VDD.n1138 4.5005
R89205 VDD.n1371 VDD.n1138 4.5005
R89206 VDD.n1321 VDD.n1138 4.5005
R89207 VDD.n1372 VDD.n1138 4.5005
R89208 VDD.n1320 VDD.n1138 4.5005
R89209 VDD.n1374 VDD.n1138 4.5005
R89210 VDD.n1319 VDD.n1138 4.5005
R89211 VDD.n1375 VDD.n1138 4.5005
R89212 VDD.n1318 VDD.n1138 4.5005
R89213 VDD.n1376 VDD.n1138 4.5005
R89214 VDD.n1316 VDD.n1138 4.5005
R89215 VDD.n1377 VDD.n1138 4.5005
R89216 VDD.n1315 VDD.n1138 4.5005
R89217 VDD.n1378 VDD.n1138 4.5005
R89218 VDD.n1313 VDD.n1138 4.5005
R89219 VDD.n1379 VDD.n1138 4.5005
R89220 VDD.n1312 VDD.n1138 4.5005
R89221 VDD.n1380 VDD.n1138 4.5005
R89222 VDD.n1310 VDD.n1138 4.5005
R89223 VDD.n1381 VDD.n1138 4.5005
R89224 VDD.n1309 VDD.n1138 4.5005
R89225 VDD.n1382 VDD.n1138 4.5005
R89226 VDD.n1307 VDD.n1138 4.5005
R89227 VDD.n1383 VDD.n1138 4.5005
R89228 VDD.n1306 VDD.n1138 4.5005
R89229 VDD.n1384 VDD.n1138 4.5005
R89230 VDD.n1304 VDD.n1138 4.5005
R89231 VDD.n1385 VDD.n1138 4.5005
R89232 VDD.n1303 VDD.n1138 4.5005
R89233 VDD.n1386 VDD.n1138 4.5005
R89234 VDD.n1301 VDD.n1138 4.5005
R89235 VDD.n1387 VDD.n1138 4.5005
R89236 VDD.n1300 VDD.n1138 4.5005
R89237 VDD.n1388 VDD.n1138 4.5005
R89238 VDD.n1298 VDD.n1138 4.5005
R89239 VDD.n1389 VDD.n1138 4.5005
R89240 VDD.n1297 VDD.n1138 4.5005
R89241 VDD.n1390 VDD.n1138 4.5005
R89242 VDD.n1295 VDD.n1138 4.5005
R89243 VDD.n1391 VDD.n1138 4.5005
R89244 VDD.n1294 VDD.n1138 4.5005
R89245 VDD.n1392 VDD.n1138 4.5005
R89246 VDD.n1292 VDD.n1138 4.5005
R89247 VDD.n1393 VDD.n1138 4.5005
R89248 VDD.n1291 VDD.n1138 4.5005
R89249 VDD.n1394 VDD.n1138 4.5005
R89250 VDD.n1289 VDD.n1138 4.5005
R89251 VDD.n1395 VDD.n1138 4.5005
R89252 VDD.n1288 VDD.n1138 4.5005
R89253 VDD.n1396 VDD.n1138 4.5005
R89254 VDD.n1286 VDD.n1138 4.5005
R89255 VDD.n1397 VDD.n1138 4.5005
R89256 VDD.n1285 VDD.n1138 4.5005
R89257 VDD.n1398 VDD.n1138 4.5005
R89258 VDD.n1283 VDD.n1138 4.5005
R89259 VDD.n1399 VDD.n1138 4.5005
R89260 VDD.n1282 VDD.n1138 4.5005
R89261 VDD.n1400 VDD.n1138 4.5005
R89262 VDD.n1280 VDD.n1138 4.5005
R89263 VDD.n1401 VDD.n1138 4.5005
R89264 VDD.n1279 VDD.n1138 4.5005
R89265 VDD.n1402 VDD.n1138 4.5005
R89266 VDD.n1277 VDD.n1138 4.5005
R89267 VDD.n1403 VDD.n1138 4.5005
R89268 VDD.n1276 VDD.n1138 4.5005
R89269 VDD.n1404 VDD.n1138 4.5005
R89270 VDD.n1274 VDD.n1138 4.5005
R89271 VDD.n1405 VDD.n1138 4.5005
R89272 VDD.n1273 VDD.n1138 4.5005
R89273 VDD.n1406 VDD.n1138 4.5005
R89274 VDD.n1271 VDD.n1138 4.5005
R89275 VDD.n1407 VDD.n1138 4.5005
R89276 VDD.n1270 VDD.n1138 4.5005
R89277 VDD.n1408 VDD.n1138 4.5005
R89278 VDD.n1268 VDD.n1138 4.5005
R89279 VDD.n1409 VDD.n1138 4.5005
R89280 VDD.n1267 VDD.n1138 4.5005
R89281 VDD.n1410 VDD.n1138 4.5005
R89282 VDD.n1265 VDD.n1138 4.5005
R89283 VDD.n1411 VDD.n1138 4.5005
R89284 VDD.n1264 VDD.n1138 4.5005
R89285 VDD.n1412 VDD.n1138 4.5005
R89286 VDD.n1262 VDD.n1138 4.5005
R89287 VDD.n1413 VDD.n1138 4.5005
R89288 VDD.n1261 VDD.n1138 4.5005
R89289 VDD.n1414 VDD.n1138 4.5005
R89290 VDD.n1415 VDD.n1138 4.5005
R89291 VDD.n1674 VDD.n1138 4.5005
R89292 VDD.n1676 VDD.n1252 4.5005
R89293 VDD.n1341 VDD.n1252 4.5005
R89294 VDD.n1342 VDD.n1252 4.5005
R89295 VDD.n1340 VDD.n1252 4.5005
R89296 VDD.n1344 VDD.n1252 4.5005
R89297 VDD.n1339 VDD.n1252 4.5005
R89298 VDD.n1345 VDD.n1252 4.5005
R89299 VDD.n1338 VDD.n1252 4.5005
R89300 VDD.n1347 VDD.n1252 4.5005
R89301 VDD.n1337 VDD.n1252 4.5005
R89302 VDD.n1348 VDD.n1252 4.5005
R89303 VDD.n1336 VDD.n1252 4.5005
R89304 VDD.n1350 VDD.n1252 4.5005
R89305 VDD.n1335 VDD.n1252 4.5005
R89306 VDD.n1351 VDD.n1252 4.5005
R89307 VDD.n1334 VDD.n1252 4.5005
R89308 VDD.n1353 VDD.n1252 4.5005
R89309 VDD.n1333 VDD.n1252 4.5005
R89310 VDD.n1354 VDD.n1252 4.5005
R89311 VDD.n1332 VDD.n1252 4.5005
R89312 VDD.n1356 VDD.n1252 4.5005
R89313 VDD.n1331 VDD.n1252 4.5005
R89314 VDD.n1357 VDD.n1252 4.5005
R89315 VDD.n1330 VDD.n1252 4.5005
R89316 VDD.n1359 VDD.n1252 4.5005
R89317 VDD.n1329 VDD.n1252 4.5005
R89318 VDD.n1360 VDD.n1252 4.5005
R89319 VDD.n1328 VDD.n1252 4.5005
R89320 VDD.n1362 VDD.n1252 4.5005
R89321 VDD.n1327 VDD.n1252 4.5005
R89322 VDD.n1363 VDD.n1252 4.5005
R89323 VDD.n1326 VDD.n1252 4.5005
R89324 VDD.n1365 VDD.n1252 4.5005
R89325 VDD.n1325 VDD.n1252 4.5005
R89326 VDD.n1366 VDD.n1252 4.5005
R89327 VDD.n1324 VDD.n1252 4.5005
R89328 VDD.n1368 VDD.n1252 4.5005
R89329 VDD.n1323 VDD.n1252 4.5005
R89330 VDD.n1369 VDD.n1252 4.5005
R89331 VDD.n1322 VDD.n1252 4.5005
R89332 VDD.n1371 VDD.n1252 4.5005
R89333 VDD.n1321 VDD.n1252 4.5005
R89334 VDD.n1372 VDD.n1252 4.5005
R89335 VDD.n1320 VDD.n1252 4.5005
R89336 VDD.n1374 VDD.n1252 4.5005
R89337 VDD.n1319 VDD.n1252 4.5005
R89338 VDD.n1375 VDD.n1252 4.5005
R89339 VDD.n1318 VDD.n1252 4.5005
R89340 VDD.n1376 VDD.n1252 4.5005
R89341 VDD.n1316 VDD.n1252 4.5005
R89342 VDD.n1377 VDD.n1252 4.5005
R89343 VDD.n1315 VDD.n1252 4.5005
R89344 VDD.n1378 VDD.n1252 4.5005
R89345 VDD.n1313 VDD.n1252 4.5005
R89346 VDD.n1379 VDD.n1252 4.5005
R89347 VDD.n1312 VDD.n1252 4.5005
R89348 VDD.n1380 VDD.n1252 4.5005
R89349 VDD.n1310 VDD.n1252 4.5005
R89350 VDD.n1381 VDD.n1252 4.5005
R89351 VDD.n1309 VDD.n1252 4.5005
R89352 VDD.n1382 VDD.n1252 4.5005
R89353 VDD.n1307 VDD.n1252 4.5005
R89354 VDD.n1383 VDD.n1252 4.5005
R89355 VDD.n1306 VDD.n1252 4.5005
R89356 VDD.n1384 VDD.n1252 4.5005
R89357 VDD.n1304 VDD.n1252 4.5005
R89358 VDD.n1385 VDD.n1252 4.5005
R89359 VDD.n1303 VDD.n1252 4.5005
R89360 VDD.n1386 VDD.n1252 4.5005
R89361 VDD.n1301 VDD.n1252 4.5005
R89362 VDD.n1387 VDD.n1252 4.5005
R89363 VDD.n1300 VDD.n1252 4.5005
R89364 VDD.n1388 VDD.n1252 4.5005
R89365 VDD.n1298 VDD.n1252 4.5005
R89366 VDD.n1389 VDD.n1252 4.5005
R89367 VDD.n1297 VDD.n1252 4.5005
R89368 VDD.n1390 VDD.n1252 4.5005
R89369 VDD.n1295 VDD.n1252 4.5005
R89370 VDD.n1391 VDD.n1252 4.5005
R89371 VDD.n1294 VDD.n1252 4.5005
R89372 VDD.n1392 VDD.n1252 4.5005
R89373 VDD.n1292 VDD.n1252 4.5005
R89374 VDD.n1393 VDD.n1252 4.5005
R89375 VDD.n1291 VDD.n1252 4.5005
R89376 VDD.n1394 VDD.n1252 4.5005
R89377 VDD.n1289 VDD.n1252 4.5005
R89378 VDD.n1395 VDD.n1252 4.5005
R89379 VDD.n1288 VDD.n1252 4.5005
R89380 VDD.n1396 VDD.n1252 4.5005
R89381 VDD.n1286 VDD.n1252 4.5005
R89382 VDD.n1397 VDD.n1252 4.5005
R89383 VDD.n1285 VDD.n1252 4.5005
R89384 VDD.n1398 VDD.n1252 4.5005
R89385 VDD.n1283 VDD.n1252 4.5005
R89386 VDD.n1399 VDD.n1252 4.5005
R89387 VDD.n1282 VDD.n1252 4.5005
R89388 VDD.n1400 VDD.n1252 4.5005
R89389 VDD.n1280 VDD.n1252 4.5005
R89390 VDD.n1401 VDD.n1252 4.5005
R89391 VDD.n1279 VDD.n1252 4.5005
R89392 VDD.n1402 VDD.n1252 4.5005
R89393 VDD.n1277 VDD.n1252 4.5005
R89394 VDD.n1403 VDD.n1252 4.5005
R89395 VDD.n1276 VDD.n1252 4.5005
R89396 VDD.n1404 VDD.n1252 4.5005
R89397 VDD.n1274 VDD.n1252 4.5005
R89398 VDD.n1405 VDD.n1252 4.5005
R89399 VDD.n1273 VDD.n1252 4.5005
R89400 VDD.n1406 VDD.n1252 4.5005
R89401 VDD.n1271 VDD.n1252 4.5005
R89402 VDD.n1407 VDD.n1252 4.5005
R89403 VDD.n1270 VDD.n1252 4.5005
R89404 VDD.n1408 VDD.n1252 4.5005
R89405 VDD.n1268 VDD.n1252 4.5005
R89406 VDD.n1409 VDD.n1252 4.5005
R89407 VDD.n1267 VDD.n1252 4.5005
R89408 VDD.n1410 VDD.n1252 4.5005
R89409 VDD.n1265 VDD.n1252 4.5005
R89410 VDD.n1411 VDD.n1252 4.5005
R89411 VDD.n1264 VDD.n1252 4.5005
R89412 VDD.n1412 VDD.n1252 4.5005
R89413 VDD.n1262 VDD.n1252 4.5005
R89414 VDD.n1413 VDD.n1252 4.5005
R89415 VDD.n1261 VDD.n1252 4.5005
R89416 VDD.n1414 VDD.n1252 4.5005
R89417 VDD.n1415 VDD.n1252 4.5005
R89418 VDD.n1674 VDD.n1252 4.5005
R89419 VDD.n1676 VDD.n1137 4.5005
R89420 VDD.n1341 VDD.n1137 4.5005
R89421 VDD.n1342 VDD.n1137 4.5005
R89422 VDD.n1340 VDD.n1137 4.5005
R89423 VDD.n1344 VDD.n1137 4.5005
R89424 VDD.n1339 VDD.n1137 4.5005
R89425 VDD.n1345 VDD.n1137 4.5005
R89426 VDD.n1338 VDD.n1137 4.5005
R89427 VDD.n1347 VDD.n1137 4.5005
R89428 VDD.n1337 VDD.n1137 4.5005
R89429 VDD.n1348 VDD.n1137 4.5005
R89430 VDD.n1336 VDD.n1137 4.5005
R89431 VDD.n1350 VDD.n1137 4.5005
R89432 VDD.n1335 VDD.n1137 4.5005
R89433 VDD.n1351 VDD.n1137 4.5005
R89434 VDD.n1334 VDD.n1137 4.5005
R89435 VDD.n1353 VDD.n1137 4.5005
R89436 VDD.n1333 VDD.n1137 4.5005
R89437 VDD.n1354 VDD.n1137 4.5005
R89438 VDD.n1332 VDD.n1137 4.5005
R89439 VDD.n1356 VDD.n1137 4.5005
R89440 VDD.n1331 VDD.n1137 4.5005
R89441 VDD.n1357 VDD.n1137 4.5005
R89442 VDD.n1330 VDD.n1137 4.5005
R89443 VDD.n1359 VDD.n1137 4.5005
R89444 VDD.n1329 VDD.n1137 4.5005
R89445 VDD.n1360 VDD.n1137 4.5005
R89446 VDD.n1328 VDD.n1137 4.5005
R89447 VDD.n1362 VDD.n1137 4.5005
R89448 VDD.n1327 VDD.n1137 4.5005
R89449 VDD.n1363 VDD.n1137 4.5005
R89450 VDD.n1326 VDD.n1137 4.5005
R89451 VDD.n1365 VDD.n1137 4.5005
R89452 VDD.n1325 VDD.n1137 4.5005
R89453 VDD.n1366 VDD.n1137 4.5005
R89454 VDD.n1324 VDD.n1137 4.5005
R89455 VDD.n1368 VDD.n1137 4.5005
R89456 VDD.n1323 VDD.n1137 4.5005
R89457 VDD.n1369 VDD.n1137 4.5005
R89458 VDD.n1322 VDD.n1137 4.5005
R89459 VDD.n1371 VDD.n1137 4.5005
R89460 VDD.n1321 VDD.n1137 4.5005
R89461 VDD.n1372 VDD.n1137 4.5005
R89462 VDD.n1320 VDD.n1137 4.5005
R89463 VDD.n1374 VDD.n1137 4.5005
R89464 VDD.n1319 VDD.n1137 4.5005
R89465 VDD.n1375 VDD.n1137 4.5005
R89466 VDD.n1318 VDD.n1137 4.5005
R89467 VDD.n1376 VDD.n1137 4.5005
R89468 VDD.n1316 VDD.n1137 4.5005
R89469 VDD.n1377 VDD.n1137 4.5005
R89470 VDD.n1315 VDD.n1137 4.5005
R89471 VDD.n1378 VDD.n1137 4.5005
R89472 VDD.n1313 VDD.n1137 4.5005
R89473 VDD.n1379 VDD.n1137 4.5005
R89474 VDD.n1312 VDD.n1137 4.5005
R89475 VDD.n1380 VDD.n1137 4.5005
R89476 VDD.n1310 VDD.n1137 4.5005
R89477 VDD.n1381 VDD.n1137 4.5005
R89478 VDD.n1309 VDD.n1137 4.5005
R89479 VDD.n1382 VDD.n1137 4.5005
R89480 VDD.n1307 VDD.n1137 4.5005
R89481 VDD.n1383 VDD.n1137 4.5005
R89482 VDD.n1306 VDD.n1137 4.5005
R89483 VDD.n1384 VDD.n1137 4.5005
R89484 VDD.n1304 VDD.n1137 4.5005
R89485 VDD.n1385 VDD.n1137 4.5005
R89486 VDD.n1303 VDD.n1137 4.5005
R89487 VDD.n1386 VDD.n1137 4.5005
R89488 VDD.n1301 VDD.n1137 4.5005
R89489 VDD.n1387 VDD.n1137 4.5005
R89490 VDD.n1300 VDD.n1137 4.5005
R89491 VDD.n1388 VDD.n1137 4.5005
R89492 VDD.n1298 VDD.n1137 4.5005
R89493 VDD.n1389 VDD.n1137 4.5005
R89494 VDD.n1297 VDD.n1137 4.5005
R89495 VDD.n1390 VDD.n1137 4.5005
R89496 VDD.n1295 VDD.n1137 4.5005
R89497 VDD.n1391 VDD.n1137 4.5005
R89498 VDD.n1294 VDD.n1137 4.5005
R89499 VDD.n1392 VDD.n1137 4.5005
R89500 VDD.n1292 VDD.n1137 4.5005
R89501 VDD.n1393 VDD.n1137 4.5005
R89502 VDD.n1291 VDD.n1137 4.5005
R89503 VDD.n1394 VDD.n1137 4.5005
R89504 VDD.n1289 VDD.n1137 4.5005
R89505 VDD.n1395 VDD.n1137 4.5005
R89506 VDD.n1288 VDD.n1137 4.5005
R89507 VDD.n1396 VDD.n1137 4.5005
R89508 VDD.n1286 VDD.n1137 4.5005
R89509 VDD.n1397 VDD.n1137 4.5005
R89510 VDD.n1285 VDD.n1137 4.5005
R89511 VDD.n1398 VDD.n1137 4.5005
R89512 VDD.n1283 VDD.n1137 4.5005
R89513 VDD.n1399 VDD.n1137 4.5005
R89514 VDD.n1282 VDD.n1137 4.5005
R89515 VDD.n1400 VDD.n1137 4.5005
R89516 VDD.n1280 VDD.n1137 4.5005
R89517 VDD.n1401 VDD.n1137 4.5005
R89518 VDD.n1279 VDD.n1137 4.5005
R89519 VDD.n1402 VDD.n1137 4.5005
R89520 VDD.n1277 VDD.n1137 4.5005
R89521 VDD.n1403 VDD.n1137 4.5005
R89522 VDD.n1276 VDD.n1137 4.5005
R89523 VDD.n1404 VDD.n1137 4.5005
R89524 VDD.n1274 VDD.n1137 4.5005
R89525 VDD.n1405 VDD.n1137 4.5005
R89526 VDD.n1273 VDD.n1137 4.5005
R89527 VDD.n1406 VDD.n1137 4.5005
R89528 VDD.n1271 VDD.n1137 4.5005
R89529 VDD.n1407 VDD.n1137 4.5005
R89530 VDD.n1270 VDD.n1137 4.5005
R89531 VDD.n1408 VDD.n1137 4.5005
R89532 VDD.n1268 VDD.n1137 4.5005
R89533 VDD.n1409 VDD.n1137 4.5005
R89534 VDD.n1267 VDD.n1137 4.5005
R89535 VDD.n1410 VDD.n1137 4.5005
R89536 VDD.n1265 VDD.n1137 4.5005
R89537 VDD.n1411 VDD.n1137 4.5005
R89538 VDD.n1264 VDD.n1137 4.5005
R89539 VDD.n1412 VDD.n1137 4.5005
R89540 VDD.n1262 VDD.n1137 4.5005
R89541 VDD.n1413 VDD.n1137 4.5005
R89542 VDD.n1261 VDD.n1137 4.5005
R89543 VDD.n1414 VDD.n1137 4.5005
R89544 VDD.n1415 VDD.n1137 4.5005
R89545 VDD.n1674 VDD.n1137 4.5005
R89546 VDD.n1676 VDD.n1253 4.5005
R89547 VDD.n1341 VDD.n1253 4.5005
R89548 VDD.n1342 VDD.n1253 4.5005
R89549 VDD.n1340 VDD.n1253 4.5005
R89550 VDD.n1344 VDD.n1253 4.5005
R89551 VDD.n1339 VDD.n1253 4.5005
R89552 VDD.n1345 VDD.n1253 4.5005
R89553 VDD.n1338 VDD.n1253 4.5005
R89554 VDD.n1347 VDD.n1253 4.5005
R89555 VDD.n1337 VDD.n1253 4.5005
R89556 VDD.n1348 VDD.n1253 4.5005
R89557 VDD.n1336 VDD.n1253 4.5005
R89558 VDD.n1350 VDD.n1253 4.5005
R89559 VDD.n1335 VDD.n1253 4.5005
R89560 VDD.n1351 VDD.n1253 4.5005
R89561 VDD.n1334 VDD.n1253 4.5005
R89562 VDD.n1353 VDD.n1253 4.5005
R89563 VDD.n1333 VDD.n1253 4.5005
R89564 VDD.n1354 VDD.n1253 4.5005
R89565 VDD.n1332 VDD.n1253 4.5005
R89566 VDD.n1356 VDD.n1253 4.5005
R89567 VDD.n1331 VDD.n1253 4.5005
R89568 VDD.n1357 VDD.n1253 4.5005
R89569 VDD.n1330 VDD.n1253 4.5005
R89570 VDD.n1359 VDD.n1253 4.5005
R89571 VDD.n1329 VDD.n1253 4.5005
R89572 VDD.n1360 VDD.n1253 4.5005
R89573 VDD.n1328 VDD.n1253 4.5005
R89574 VDD.n1362 VDD.n1253 4.5005
R89575 VDD.n1327 VDD.n1253 4.5005
R89576 VDD.n1363 VDD.n1253 4.5005
R89577 VDD.n1326 VDD.n1253 4.5005
R89578 VDD.n1365 VDD.n1253 4.5005
R89579 VDD.n1325 VDD.n1253 4.5005
R89580 VDD.n1366 VDD.n1253 4.5005
R89581 VDD.n1324 VDD.n1253 4.5005
R89582 VDD.n1368 VDD.n1253 4.5005
R89583 VDD.n1323 VDD.n1253 4.5005
R89584 VDD.n1369 VDD.n1253 4.5005
R89585 VDD.n1322 VDD.n1253 4.5005
R89586 VDD.n1371 VDD.n1253 4.5005
R89587 VDD.n1321 VDD.n1253 4.5005
R89588 VDD.n1372 VDD.n1253 4.5005
R89589 VDD.n1320 VDD.n1253 4.5005
R89590 VDD.n1374 VDD.n1253 4.5005
R89591 VDD.n1319 VDD.n1253 4.5005
R89592 VDD.n1375 VDD.n1253 4.5005
R89593 VDD.n1318 VDD.n1253 4.5005
R89594 VDD.n1376 VDD.n1253 4.5005
R89595 VDD.n1316 VDD.n1253 4.5005
R89596 VDD.n1377 VDD.n1253 4.5005
R89597 VDD.n1315 VDD.n1253 4.5005
R89598 VDD.n1378 VDD.n1253 4.5005
R89599 VDD.n1313 VDD.n1253 4.5005
R89600 VDD.n1379 VDD.n1253 4.5005
R89601 VDD.n1312 VDD.n1253 4.5005
R89602 VDD.n1380 VDD.n1253 4.5005
R89603 VDD.n1310 VDD.n1253 4.5005
R89604 VDD.n1381 VDD.n1253 4.5005
R89605 VDD.n1309 VDD.n1253 4.5005
R89606 VDD.n1382 VDD.n1253 4.5005
R89607 VDD.n1307 VDD.n1253 4.5005
R89608 VDD.n1383 VDD.n1253 4.5005
R89609 VDD.n1306 VDD.n1253 4.5005
R89610 VDD.n1384 VDD.n1253 4.5005
R89611 VDD.n1304 VDD.n1253 4.5005
R89612 VDD.n1385 VDD.n1253 4.5005
R89613 VDD.n1303 VDD.n1253 4.5005
R89614 VDD.n1386 VDD.n1253 4.5005
R89615 VDD.n1301 VDD.n1253 4.5005
R89616 VDD.n1387 VDD.n1253 4.5005
R89617 VDD.n1300 VDD.n1253 4.5005
R89618 VDD.n1388 VDD.n1253 4.5005
R89619 VDD.n1298 VDD.n1253 4.5005
R89620 VDD.n1389 VDD.n1253 4.5005
R89621 VDD.n1297 VDD.n1253 4.5005
R89622 VDD.n1390 VDD.n1253 4.5005
R89623 VDD.n1295 VDD.n1253 4.5005
R89624 VDD.n1391 VDD.n1253 4.5005
R89625 VDD.n1294 VDD.n1253 4.5005
R89626 VDD.n1392 VDD.n1253 4.5005
R89627 VDD.n1292 VDD.n1253 4.5005
R89628 VDD.n1393 VDD.n1253 4.5005
R89629 VDD.n1291 VDD.n1253 4.5005
R89630 VDD.n1394 VDD.n1253 4.5005
R89631 VDD.n1289 VDD.n1253 4.5005
R89632 VDD.n1395 VDD.n1253 4.5005
R89633 VDD.n1288 VDD.n1253 4.5005
R89634 VDD.n1396 VDD.n1253 4.5005
R89635 VDD.n1286 VDD.n1253 4.5005
R89636 VDD.n1397 VDD.n1253 4.5005
R89637 VDD.n1285 VDD.n1253 4.5005
R89638 VDD.n1398 VDD.n1253 4.5005
R89639 VDD.n1283 VDD.n1253 4.5005
R89640 VDD.n1399 VDD.n1253 4.5005
R89641 VDD.n1282 VDD.n1253 4.5005
R89642 VDD.n1400 VDD.n1253 4.5005
R89643 VDD.n1280 VDD.n1253 4.5005
R89644 VDD.n1401 VDD.n1253 4.5005
R89645 VDD.n1279 VDD.n1253 4.5005
R89646 VDD.n1402 VDD.n1253 4.5005
R89647 VDD.n1277 VDD.n1253 4.5005
R89648 VDD.n1403 VDD.n1253 4.5005
R89649 VDD.n1276 VDD.n1253 4.5005
R89650 VDD.n1404 VDD.n1253 4.5005
R89651 VDD.n1274 VDD.n1253 4.5005
R89652 VDD.n1405 VDD.n1253 4.5005
R89653 VDD.n1273 VDD.n1253 4.5005
R89654 VDD.n1406 VDD.n1253 4.5005
R89655 VDD.n1271 VDD.n1253 4.5005
R89656 VDD.n1407 VDD.n1253 4.5005
R89657 VDD.n1270 VDD.n1253 4.5005
R89658 VDD.n1408 VDD.n1253 4.5005
R89659 VDD.n1268 VDD.n1253 4.5005
R89660 VDD.n1409 VDD.n1253 4.5005
R89661 VDD.n1267 VDD.n1253 4.5005
R89662 VDD.n1410 VDD.n1253 4.5005
R89663 VDD.n1265 VDD.n1253 4.5005
R89664 VDD.n1411 VDD.n1253 4.5005
R89665 VDD.n1264 VDD.n1253 4.5005
R89666 VDD.n1412 VDD.n1253 4.5005
R89667 VDD.n1262 VDD.n1253 4.5005
R89668 VDD.n1413 VDD.n1253 4.5005
R89669 VDD.n1261 VDD.n1253 4.5005
R89670 VDD.n1414 VDD.n1253 4.5005
R89671 VDD.n1415 VDD.n1253 4.5005
R89672 VDD.n1674 VDD.n1253 4.5005
R89673 VDD.n1676 VDD.n1136 4.5005
R89674 VDD.n1341 VDD.n1136 4.5005
R89675 VDD.n1342 VDD.n1136 4.5005
R89676 VDD.n1340 VDD.n1136 4.5005
R89677 VDD.n1344 VDD.n1136 4.5005
R89678 VDD.n1339 VDD.n1136 4.5005
R89679 VDD.n1345 VDD.n1136 4.5005
R89680 VDD.n1338 VDD.n1136 4.5005
R89681 VDD.n1347 VDD.n1136 4.5005
R89682 VDD.n1337 VDD.n1136 4.5005
R89683 VDD.n1348 VDD.n1136 4.5005
R89684 VDD.n1336 VDD.n1136 4.5005
R89685 VDD.n1350 VDD.n1136 4.5005
R89686 VDD.n1335 VDD.n1136 4.5005
R89687 VDD.n1351 VDD.n1136 4.5005
R89688 VDD.n1334 VDD.n1136 4.5005
R89689 VDD.n1353 VDD.n1136 4.5005
R89690 VDD.n1333 VDD.n1136 4.5005
R89691 VDD.n1354 VDD.n1136 4.5005
R89692 VDD.n1332 VDD.n1136 4.5005
R89693 VDD.n1356 VDD.n1136 4.5005
R89694 VDD.n1331 VDD.n1136 4.5005
R89695 VDD.n1357 VDD.n1136 4.5005
R89696 VDD.n1330 VDD.n1136 4.5005
R89697 VDD.n1359 VDD.n1136 4.5005
R89698 VDD.n1329 VDD.n1136 4.5005
R89699 VDD.n1360 VDD.n1136 4.5005
R89700 VDD.n1328 VDD.n1136 4.5005
R89701 VDD.n1362 VDD.n1136 4.5005
R89702 VDD.n1327 VDD.n1136 4.5005
R89703 VDD.n1363 VDD.n1136 4.5005
R89704 VDD.n1326 VDD.n1136 4.5005
R89705 VDD.n1365 VDD.n1136 4.5005
R89706 VDD.n1325 VDD.n1136 4.5005
R89707 VDD.n1366 VDD.n1136 4.5005
R89708 VDD.n1324 VDD.n1136 4.5005
R89709 VDD.n1368 VDD.n1136 4.5005
R89710 VDD.n1323 VDD.n1136 4.5005
R89711 VDD.n1369 VDD.n1136 4.5005
R89712 VDD.n1322 VDD.n1136 4.5005
R89713 VDD.n1371 VDD.n1136 4.5005
R89714 VDD.n1321 VDD.n1136 4.5005
R89715 VDD.n1372 VDD.n1136 4.5005
R89716 VDD.n1320 VDD.n1136 4.5005
R89717 VDD.n1374 VDD.n1136 4.5005
R89718 VDD.n1319 VDD.n1136 4.5005
R89719 VDD.n1375 VDD.n1136 4.5005
R89720 VDD.n1318 VDD.n1136 4.5005
R89721 VDD.n1376 VDD.n1136 4.5005
R89722 VDD.n1316 VDD.n1136 4.5005
R89723 VDD.n1377 VDD.n1136 4.5005
R89724 VDD.n1315 VDD.n1136 4.5005
R89725 VDD.n1378 VDD.n1136 4.5005
R89726 VDD.n1313 VDD.n1136 4.5005
R89727 VDD.n1379 VDD.n1136 4.5005
R89728 VDD.n1312 VDD.n1136 4.5005
R89729 VDD.n1380 VDD.n1136 4.5005
R89730 VDD.n1310 VDD.n1136 4.5005
R89731 VDD.n1381 VDD.n1136 4.5005
R89732 VDD.n1309 VDD.n1136 4.5005
R89733 VDD.n1382 VDD.n1136 4.5005
R89734 VDD.n1307 VDD.n1136 4.5005
R89735 VDD.n1383 VDD.n1136 4.5005
R89736 VDD.n1306 VDD.n1136 4.5005
R89737 VDD.n1384 VDD.n1136 4.5005
R89738 VDD.n1304 VDD.n1136 4.5005
R89739 VDD.n1385 VDD.n1136 4.5005
R89740 VDD.n1303 VDD.n1136 4.5005
R89741 VDD.n1386 VDD.n1136 4.5005
R89742 VDD.n1301 VDD.n1136 4.5005
R89743 VDD.n1387 VDD.n1136 4.5005
R89744 VDD.n1300 VDD.n1136 4.5005
R89745 VDD.n1388 VDD.n1136 4.5005
R89746 VDD.n1298 VDD.n1136 4.5005
R89747 VDD.n1389 VDD.n1136 4.5005
R89748 VDD.n1297 VDD.n1136 4.5005
R89749 VDD.n1390 VDD.n1136 4.5005
R89750 VDD.n1295 VDD.n1136 4.5005
R89751 VDD.n1391 VDD.n1136 4.5005
R89752 VDD.n1294 VDD.n1136 4.5005
R89753 VDD.n1392 VDD.n1136 4.5005
R89754 VDD.n1292 VDD.n1136 4.5005
R89755 VDD.n1393 VDD.n1136 4.5005
R89756 VDD.n1291 VDD.n1136 4.5005
R89757 VDD.n1394 VDD.n1136 4.5005
R89758 VDD.n1289 VDD.n1136 4.5005
R89759 VDD.n1395 VDD.n1136 4.5005
R89760 VDD.n1288 VDD.n1136 4.5005
R89761 VDD.n1396 VDD.n1136 4.5005
R89762 VDD.n1286 VDD.n1136 4.5005
R89763 VDD.n1397 VDD.n1136 4.5005
R89764 VDD.n1285 VDD.n1136 4.5005
R89765 VDD.n1398 VDD.n1136 4.5005
R89766 VDD.n1283 VDD.n1136 4.5005
R89767 VDD.n1399 VDD.n1136 4.5005
R89768 VDD.n1282 VDD.n1136 4.5005
R89769 VDD.n1400 VDD.n1136 4.5005
R89770 VDD.n1280 VDD.n1136 4.5005
R89771 VDD.n1401 VDD.n1136 4.5005
R89772 VDD.n1279 VDD.n1136 4.5005
R89773 VDD.n1402 VDD.n1136 4.5005
R89774 VDD.n1277 VDD.n1136 4.5005
R89775 VDD.n1403 VDD.n1136 4.5005
R89776 VDD.n1276 VDD.n1136 4.5005
R89777 VDD.n1404 VDD.n1136 4.5005
R89778 VDD.n1274 VDD.n1136 4.5005
R89779 VDD.n1405 VDD.n1136 4.5005
R89780 VDD.n1273 VDD.n1136 4.5005
R89781 VDD.n1406 VDD.n1136 4.5005
R89782 VDD.n1271 VDD.n1136 4.5005
R89783 VDD.n1407 VDD.n1136 4.5005
R89784 VDD.n1270 VDD.n1136 4.5005
R89785 VDD.n1408 VDD.n1136 4.5005
R89786 VDD.n1268 VDD.n1136 4.5005
R89787 VDD.n1409 VDD.n1136 4.5005
R89788 VDD.n1267 VDD.n1136 4.5005
R89789 VDD.n1410 VDD.n1136 4.5005
R89790 VDD.n1265 VDD.n1136 4.5005
R89791 VDD.n1411 VDD.n1136 4.5005
R89792 VDD.n1264 VDD.n1136 4.5005
R89793 VDD.n1412 VDD.n1136 4.5005
R89794 VDD.n1262 VDD.n1136 4.5005
R89795 VDD.n1413 VDD.n1136 4.5005
R89796 VDD.n1261 VDD.n1136 4.5005
R89797 VDD.n1414 VDD.n1136 4.5005
R89798 VDD.n1415 VDD.n1136 4.5005
R89799 VDD.n1674 VDD.n1136 4.5005
R89800 VDD.n1676 VDD.n1254 4.5005
R89801 VDD.n1341 VDD.n1254 4.5005
R89802 VDD.n1342 VDD.n1254 4.5005
R89803 VDD.n1340 VDD.n1254 4.5005
R89804 VDD.n1344 VDD.n1254 4.5005
R89805 VDD.n1339 VDD.n1254 4.5005
R89806 VDD.n1345 VDD.n1254 4.5005
R89807 VDD.n1338 VDD.n1254 4.5005
R89808 VDD.n1347 VDD.n1254 4.5005
R89809 VDD.n1337 VDD.n1254 4.5005
R89810 VDD.n1348 VDD.n1254 4.5005
R89811 VDD.n1336 VDD.n1254 4.5005
R89812 VDD.n1350 VDD.n1254 4.5005
R89813 VDD.n1335 VDD.n1254 4.5005
R89814 VDD.n1351 VDD.n1254 4.5005
R89815 VDD.n1334 VDD.n1254 4.5005
R89816 VDD.n1353 VDD.n1254 4.5005
R89817 VDD.n1333 VDD.n1254 4.5005
R89818 VDD.n1354 VDD.n1254 4.5005
R89819 VDD.n1332 VDD.n1254 4.5005
R89820 VDD.n1356 VDD.n1254 4.5005
R89821 VDD.n1331 VDD.n1254 4.5005
R89822 VDD.n1357 VDD.n1254 4.5005
R89823 VDD.n1330 VDD.n1254 4.5005
R89824 VDD.n1359 VDD.n1254 4.5005
R89825 VDD.n1329 VDD.n1254 4.5005
R89826 VDD.n1360 VDD.n1254 4.5005
R89827 VDD.n1328 VDD.n1254 4.5005
R89828 VDD.n1362 VDD.n1254 4.5005
R89829 VDD.n1327 VDD.n1254 4.5005
R89830 VDD.n1363 VDD.n1254 4.5005
R89831 VDD.n1326 VDD.n1254 4.5005
R89832 VDD.n1365 VDD.n1254 4.5005
R89833 VDD.n1325 VDD.n1254 4.5005
R89834 VDD.n1366 VDD.n1254 4.5005
R89835 VDD.n1324 VDD.n1254 4.5005
R89836 VDD.n1368 VDD.n1254 4.5005
R89837 VDD.n1323 VDD.n1254 4.5005
R89838 VDD.n1369 VDD.n1254 4.5005
R89839 VDD.n1322 VDD.n1254 4.5005
R89840 VDD.n1371 VDD.n1254 4.5005
R89841 VDD.n1321 VDD.n1254 4.5005
R89842 VDD.n1372 VDD.n1254 4.5005
R89843 VDD.n1320 VDD.n1254 4.5005
R89844 VDD.n1374 VDD.n1254 4.5005
R89845 VDD.n1319 VDD.n1254 4.5005
R89846 VDD.n1375 VDD.n1254 4.5005
R89847 VDD.n1318 VDD.n1254 4.5005
R89848 VDD.n1376 VDD.n1254 4.5005
R89849 VDD.n1316 VDD.n1254 4.5005
R89850 VDD.n1377 VDD.n1254 4.5005
R89851 VDD.n1315 VDD.n1254 4.5005
R89852 VDD.n1378 VDD.n1254 4.5005
R89853 VDD.n1313 VDD.n1254 4.5005
R89854 VDD.n1379 VDD.n1254 4.5005
R89855 VDD.n1312 VDD.n1254 4.5005
R89856 VDD.n1380 VDD.n1254 4.5005
R89857 VDD.n1310 VDD.n1254 4.5005
R89858 VDD.n1381 VDD.n1254 4.5005
R89859 VDD.n1309 VDD.n1254 4.5005
R89860 VDD.n1382 VDD.n1254 4.5005
R89861 VDD.n1307 VDD.n1254 4.5005
R89862 VDD.n1383 VDD.n1254 4.5005
R89863 VDD.n1306 VDD.n1254 4.5005
R89864 VDD.n1384 VDD.n1254 4.5005
R89865 VDD.n1304 VDD.n1254 4.5005
R89866 VDD.n1385 VDD.n1254 4.5005
R89867 VDD.n1303 VDD.n1254 4.5005
R89868 VDD.n1386 VDD.n1254 4.5005
R89869 VDD.n1301 VDD.n1254 4.5005
R89870 VDD.n1387 VDD.n1254 4.5005
R89871 VDD.n1300 VDD.n1254 4.5005
R89872 VDD.n1388 VDD.n1254 4.5005
R89873 VDD.n1298 VDD.n1254 4.5005
R89874 VDD.n1389 VDD.n1254 4.5005
R89875 VDD.n1297 VDD.n1254 4.5005
R89876 VDD.n1390 VDD.n1254 4.5005
R89877 VDD.n1295 VDD.n1254 4.5005
R89878 VDD.n1391 VDD.n1254 4.5005
R89879 VDD.n1294 VDD.n1254 4.5005
R89880 VDD.n1392 VDD.n1254 4.5005
R89881 VDD.n1292 VDD.n1254 4.5005
R89882 VDD.n1393 VDD.n1254 4.5005
R89883 VDD.n1291 VDD.n1254 4.5005
R89884 VDD.n1394 VDD.n1254 4.5005
R89885 VDD.n1289 VDD.n1254 4.5005
R89886 VDD.n1395 VDD.n1254 4.5005
R89887 VDD.n1288 VDD.n1254 4.5005
R89888 VDD.n1396 VDD.n1254 4.5005
R89889 VDD.n1286 VDD.n1254 4.5005
R89890 VDD.n1397 VDD.n1254 4.5005
R89891 VDD.n1285 VDD.n1254 4.5005
R89892 VDD.n1398 VDD.n1254 4.5005
R89893 VDD.n1283 VDD.n1254 4.5005
R89894 VDD.n1399 VDD.n1254 4.5005
R89895 VDD.n1282 VDD.n1254 4.5005
R89896 VDD.n1400 VDD.n1254 4.5005
R89897 VDD.n1280 VDD.n1254 4.5005
R89898 VDD.n1401 VDD.n1254 4.5005
R89899 VDD.n1279 VDD.n1254 4.5005
R89900 VDD.n1402 VDD.n1254 4.5005
R89901 VDD.n1277 VDD.n1254 4.5005
R89902 VDD.n1403 VDD.n1254 4.5005
R89903 VDD.n1276 VDD.n1254 4.5005
R89904 VDD.n1404 VDD.n1254 4.5005
R89905 VDD.n1274 VDD.n1254 4.5005
R89906 VDD.n1405 VDD.n1254 4.5005
R89907 VDD.n1273 VDD.n1254 4.5005
R89908 VDD.n1406 VDD.n1254 4.5005
R89909 VDD.n1271 VDD.n1254 4.5005
R89910 VDD.n1407 VDD.n1254 4.5005
R89911 VDD.n1270 VDD.n1254 4.5005
R89912 VDD.n1408 VDD.n1254 4.5005
R89913 VDD.n1268 VDD.n1254 4.5005
R89914 VDD.n1409 VDD.n1254 4.5005
R89915 VDD.n1267 VDD.n1254 4.5005
R89916 VDD.n1410 VDD.n1254 4.5005
R89917 VDD.n1265 VDD.n1254 4.5005
R89918 VDD.n1411 VDD.n1254 4.5005
R89919 VDD.n1264 VDD.n1254 4.5005
R89920 VDD.n1412 VDD.n1254 4.5005
R89921 VDD.n1262 VDD.n1254 4.5005
R89922 VDD.n1413 VDD.n1254 4.5005
R89923 VDD.n1261 VDD.n1254 4.5005
R89924 VDD.n1414 VDD.n1254 4.5005
R89925 VDD.n1415 VDD.n1254 4.5005
R89926 VDD.n1674 VDD.n1254 4.5005
R89927 VDD.n1676 VDD.n1135 4.5005
R89928 VDD.n1341 VDD.n1135 4.5005
R89929 VDD.n1342 VDD.n1135 4.5005
R89930 VDD.n1340 VDD.n1135 4.5005
R89931 VDD.n1344 VDD.n1135 4.5005
R89932 VDD.n1339 VDD.n1135 4.5005
R89933 VDD.n1345 VDD.n1135 4.5005
R89934 VDD.n1338 VDD.n1135 4.5005
R89935 VDD.n1347 VDD.n1135 4.5005
R89936 VDD.n1337 VDD.n1135 4.5005
R89937 VDD.n1348 VDD.n1135 4.5005
R89938 VDD.n1336 VDD.n1135 4.5005
R89939 VDD.n1350 VDD.n1135 4.5005
R89940 VDD.n1335 VDD.n1135 4.5005
R89941 VDD.n1351 VDD.n1135 4.5005
R89942 VDD.n1334 VDD.n1135 4.5005
R89943 VDD.n1353 VDD.n1135 4.5005
R89944 VDD.n1333 VDD.n1135 4.5005
R89945 VDD.n1354 VDD.n1135 4.5005
R89946 VDD.n1332 VDD.n1135 4.5005
R89947 VDD.n1356 VDD.n1135 4.5005
R89948 VDD.n1331 VDD.n1135 4.5005
R89949 VDD.n1357 VDD.n1135 4.5005
R89950 VDD.n1330 VDD.n1135 4.5005
R89951 VDD.n1359 VDD.n1135 4.5005
R89952 VDD.n1329 VDD.n1135 4.5005
R89953 VDD.n1360 VDD.n1135 4.5005
R89954 VDD.n1328 VDD.n1135 4.5005
R89955 VDD.n1362 VDD.n1135 4.5005
R89956 VDD.n1327 VDD.n1135 4.5005
R89957 VDD.n1363 VDD.n1135 4.5005
R89958 VDD.n1326 VDD.n1135 4.5005
R89959 VDD.n1365 VDD.n1135 4.5005
R89960 VDD.n1325 VDD.n1135 4.5005
R89961 VDD.n1366 VDD.n1135 4.5005
R89962 VDD.n1324 VDD.n1135 4.5005
R89963 VDD.n1368 VDD.n1135 4.5005
R89964 VDD.n1323 VDD.n1135 4.5005
R89965 VDD.n1369 VDD.n1135 4.5005
R89966 VDD.n1322 VDD.n1135 4.5005
R89967 VDD.n1371 VDD.n1135 4.5005
R89968 VDD.n1321 VDD.n1135 4.5005
R89969 VDD.n1372 VDD.n1135 4.5005
R89970 VDD.n1320 VDD.n1135 4.5005
R89971 VDD.n1374 VDD.n1135 4.5005
R89972 VDD.n1319 VDD.n1135 4.5005
R89973 VDD.n1375 VDD.n1135 4.5005
R89974 VDD.n1318 VDD.n1135 4.5005
R89975 VDD.n1376 VDD.n1135 4.5005
R89976 VDD.n1316 VDD.n1135 4.5005
R89977 VDD.n1377 VDD.n1135 4.5005
R89978 VDD.n1315 VDD.n1135 4.5005
R89979 VDD.n1378 VDD.n1135 4.5005
R89980 VDD.n1313 VDD.n1135 4.5005
R89981 VDD.n1379 VDD.n1135 4.5005
R89982 VDD.n1312 VDD.n1135 4.5005
R89983 VDD.n1380 VDD.n1135 4.5005
R89984 VDD.n1310 VDD.n1135 4.5005
R89985 VDD.n1381 VDD.n1135 4.5005
R89986 VDD.n1309 VDD.n1135 4.5005
R89987 VDD.n1382 VDD.n1135 4.5005
R89988 VDD.n1307 VDD.n1135 4.5005
R89989 VDD.n1383 VDD.n1135 4.5005
R89990 VDD.n1306 VDD.n1135 4.5005
R89991 VDD.n1384 VDD.n1135 4.5005
R89992 VDD.n1304 VDD.n1135 4.5005
R89993 VDD.n1385 VDD.n1135 4.5005
R89994 VDD.n1303 VDD.n1135 4.5005
R89995 VDD.n1386 VDD.n1135 4.5005
R89996 VDD.n1301 VDD.n1135 4.5005
R89997 VDD.n1387 VDD.n1135 4.5005
R89998 VDD.n1300 VDD.n1135 4.5005
R89999 VDD.n1388 VDD.n1135 4.5005
R90000 VDD.n1298 VDD.n1135 4.5005
R90001 VDD.n1389 VDD.n1135 4.5005
R90002 VDD.n1297 VDD.n1135 4.5005
R90003 VDD.n1390 VDD.n1135 4.5005
R90004 VDD.n1295 VDD.n1135 4.5005
R90005 VDD.n1391 VDD.n1135 4.5005
R90006 VDD.n1294 VDD.n1135 4.5005
R90007 VDD.n1392 VDD.n1135 4.5005
R90008 VDD.n1292 VDD.n1135 4.5005
R90009 VDD.n1393 VDD.n1135 4.5005
R90010 VDD.n1291 VDD.n1135 4.5005
R90011 VDD.n1394 VDD.n1135 4.5005
R90012 VDD.n1289 VDD.n1135 4.5005
R90013 VDD.n1395 VDD.n1135 4.5005
R90014 VDD.n1288 VDD.n1135 4.5005
R90015 VDD.n1396 VDD.n1135 4.5005
R90016 VDD.n1286 VDD.n1135 4.5005
R90017 VDD.n1397 VDD.n1135 4.5005
R90018 VDD.n1285 VDD.n1135 4.5005
R90019 VDD.n1398 VDD.n1135 4.5005
R90020 VDD.n1283 VDD.n1135 4.5005
R90021 VDD.n1399 VDD.n1135 4.5005
R90022 VDD.n1282 VDD.n1135 4.5005
R90023 VDD.n1400 VDD.n1135 4.5005
R90024 VDD.n1280 VDD.n1135 4.5005
R90025 VDD.n1401 VDD.n1135 4.5005
R90026 VDD.n1279 VDD.n1135 4.5005
R90027 VDD.n1402 VDD.n1135 4.5005
R90028 VDD.n1277 VDD.n1135 4.5005
R90029 VDD.n1403 VDD.n1135 4.5005
R90030 VDD.n1276 VDD.n1135 4.5005
R90031 VDD.n1404 VDD.n1135 4.5005
R90032 VDD.n1274 VDD.n1135 4.5005
R90033 VDD.n1405 VDD.n1135 4.5005
R90034 VDD.n1273 VDD.n1135 4.5005
R90035 VDD.n1406 VDD.n1135 4.5005
R90036 VDD.n1271 VDD.n1135 4.5005
R90037 VDD.n1407 VDD.n1135 4.5005
R90038 VDD.n1270 VDD.n1135 4.5005
R90039 VDD.n1408 VDD.n1135 4.5005
R90040 VDD.n1268 VDD.n1135 4.5005
R90041 VDD.n1409 VDD.n1135 4.5005
R90042 VDD.n1267 VDD.n1135 4.5005
R90043 VDD.n1410 VDD.n1135 4.5005
R90044 VDD.n1265 VDD.n1135 4.5005
R90045 VDD.n1411 VDD.n1135 4.5005
R90046 VDD.n1264 VDD.n1135 4.5005
R90047 VDD.n1412 VDD.n1135 4.5005
R90048 VDD.n1262 VDD.n1135 4.5005
R90049 VDD.n1413 VDD.n1135 4.5005
R90050 VDD.n1261 VDD.n1135 4.5005
R90051 VDD.n1414 VDD.n1135 4.5005
R90052 VDD.n1415 VDD.n1135 4.5005
R90053 VDD.n1674 VDD.n1135 4.5005
R90054 VDD.n1676 VDD.n1255 4.5005
R90055 VDD.n1341 VDD.n1255 4.5005
R90056 VDD.n1342 VDD.n1255 4.5005
R90057 VDD.n1340 VDD.n1255 4.5005
R90058 VDD.n1344 VDD.n1255 4.5005
R90059 VDD.n1339 VDD.n1255 4.5005
R90060 VDD.n1345 VDD.n1255 4.5005
R90061 VDD.n1338 VDD.n1255 4.5005
R90062 VDD.n1347 VDD.n1255 4.5005
R90063 VDD.n1337 VDD.n1255 4.5005
R90064 VDD.n1348 VDD.n1255 4.5005
R90065 VDD.n1336 VDD.n1255 4.5005
R90066 VDD.n1350 VDD.n1255 4.5005
R90067 VDD.n1335 VDD.n1255 4.5005
R90068 VDD.n1351 VDD.n1255 4.5005
R90069 VDD.n1334 VDD.n1255 4.5005
R90070 VDD.n1353 VDD.n1255 4.5005
R90071 VDD.n1333 VDD.n1255 4.5005
R90072 VDD.n1354 VDD.n1255 4.5005
R90073 VDD.n1332 VDD.n1255 4.5005
R90074 VDD.n1356 VDD.n1255 4.5005
R90075 VDD.n1331 VDD.n1255 4.5005
R90076 VDD.n1357 VDD.n1255 4.5005
R90077 VDD.n1330 VDD.n1255 4.5005
R90078 VDD.n1359 VDD.n1255 4.5005
R90079 VDD.n1329 VDD.n1255 4.5005
R90080 VDD.n1360 VDD.n1255 4.5005
R90081 VDD.n1328 VDD.n1255 4.5005
R90082 VDD.n1362 VDD.n1255 4.5005
R90083 VDD.n1327 VDD.n1255 4.5005
R90084 VDD.n1363 VDD.n1255 4.5005
R90085 VDD.n1326 VDD.n1255 4.5005
R90086 VDD.n1365 VDD.n1255 4.5005
R90087 VDD.n1325 VDD.n1255 4.5005
R90088 VDD.n1366 VDD.n1255 4.5005
R90089 VDD.n1324 VDD.n1255 4.5005
R90090 VDD.n1368 VDD.n1255 4.5005
R90091 VDD.n1323 VDD.n1255 4.5005
R90092 VDD.n1369 VDD.n1255 4.5005
R90093 VDD.n1322 VDD.n1255 4.5005
R90094 VDD.n1371 VDD.n1255 4.5005
R90095 VDD.n1321 VDD.n1255 4.5005
R90096 VDD.n1372 VDD.n1255 4.5005
R90097 VDD.n1320 VDD.n1255 4.5005
R90098 VDD.n1374 VDD.n1255 4.5005
R90099 VDD.n1319 VDD.n1255 4.5005
R90100 VDD.n1375 VDD.n1255 4.5005
R90101 VDD.n1318 VDD.n1255 4.5005
R90102 VDD.n1376 VDD.n1255 4.5005
R90103 VDD.n1316 VDD.n1255 4.5005
R90104 VDD.n1377 VDD.n1255 4.5005
R90105 VDD.n1315 VDD.n1255 4.5005
R90106 VDD.n1378 VDD.n1255 4.5005
R90107 VDD.n1313 VDD.n1255 4.5005
R90108 VDD.n1379 VDD.n1255 4.5005
R90109 VDD.n1312 VDD.n1255 4.5005
R90110 VDD.n1380 VDD.n1255 4.5005
R90111 VDD.n1310 VDD.n1255 4.5005
R90112 VDD.n1381 VDD.n1255 4.5005
R90113 VDD.n1309 VDD.n1255 4.5005
R90114 VDD.n1382 VDD.n1255 4.5005
R90115 VDD.n1307 VDD.n1255 4.5005
R90116 VDD.n1383 VDD.n1255 4.5005
R90117 VDD.n1306 VDD.n1255 4.5005
R90118 VDD.n1384 VDD.n1255 4.5005
R90119 VDD.n1304 VDD.n1255 4.5005
R90120 VDD.n1385 VDD.n1255 4.5005
R90121 VDD.n1303 VDD.n1255 4.5005
R90122 VDD.n1386 VDD.n1255 4.5005
R90123 VDD.n1301 VDD.n1255 4.5005
R90124 VDD.n1387 VDD.n1255 4.5005
R90125 VDD.n1300 VDD.n1255 4.5005
R90126 VDD.n1388 VDD.n1255 4.5005
R90127 VDD.n1298 VDD.n1255 4.5005
R90128 VDD.n1389 VDD.n1255 4.5005
R90129 VDD.n1297 VDD.n1255 4.5005
R90130 VDD.n1390 VDD.n1255 4.5005
R90131 VDD.n1295 VDD.n1255 4.5005
R90132 VDD.n1391 VDD.n1255 4.5005
R90133 VDD.n1294 VDD.n1255 4.5005
R90134 VDD.n1392 VDD.n1255 4.5005
R90135 VDD.n1292 VDD.n1255 4.5005
R90136 VDD.n1393 VDD.n1255 4.5005
R90137 VDD.n1291 VDD.n1255 4.5005
R90138 VDD.n1394 VDD.n1255 4.5005
R90139 VDD.n1289 VDD.n1255 4.5005
R90140 VDD.n1395 VDD.n1255 4.5005
R90141 VDD.n1288 VDD.n1255 4.5005
R90142 VDD.n1396 VDD.n1255 4.5005
R90143 VDD.n1286 VDD.n1255 4.5005
R90144 VDD.n1397 VDD.n1255 4.5005
R90145 VDD.n1285 VDD.n1255 4.5005
R90146 VDD.n1398 VDD.n1255 4.5005
R90147 VDD.n1283 VDD.n1255 4.5005
R90148 VDD.n1399 VDD.n1255 4.5005
R90149 VDD.n1282 VDD.n1255 4.5005
R90150 VDD.n1400 VDD.n1255 4.5005
R90151 VDD.n1280 VDD.n1255 4.5005
R90152 VDD.n1401 VDD.n1255 4.5005
R90153 VDD.n1279 VDD.n1255 4.5005
R90154 VDD.n1402 VDD.n1255 4.5005
R90155 VDD.n1277 VDD.n1255 4.5005
R90156 VDD.n1403 VDD.n1255 4.5005
R90157 VDD.n1276 VDD.n1255 4.5005
R90158 VDD.n1404 VDD.n1255 4.5005
R90159 VDD.n1274 VDD.n1255 4.5005
R90160 VDD.n1405 VDD.n1255 4.5005
R90161 VDD.n1273 VDD.n1255 4.5005
R90162 VDD.n1406 VDD.n1255 4.5005
R90163 VDD.n1271 VDD.n1255 4.5005
R90164 VDD.n1407 VDD.n1255 4.5005
R90165 VDD.n1270 VDD.n1255 4.5005
R90166 VDD.n1408 VDD.n1255 4.5005
R90167 VDD.n1268 VDD.n1255 4.5005
R90168 VDD.n1409 VDD.n1255 4.5005
R90169 VDD.n1267 VDD.n1255 4.5005
R90170 VDD.n1410 VDD.n1255 4.5005
R90171 VDD.n1265 VDD.n1255 4.5005
R90172 VDD.n1411 VDD.n1255 4.5005
R90173 VDD.n1264 VDD.n1255 4.5005
R90174 VDD.n1412 VDD.n1255 4.5005
R90175 VDD.n1262 VDD.n1255 4.5005
R90176 VDD.n1413 VDD.n1255 4.5005
R90177 VDD.n1261 VDD.n1255 4.5005
R90178 VDD.n1414 VDD.n1255 4.5005
R90179 VDD.n1415 VDD.n1255 4.5005
R90180 VDD.n1674 VDD.n1255 4.5005
R90181 VDD.n1676 VDD.n1134 4.5005
R90182 VDD.n1341 VDD.n1134 4.5005
R90183 VDD.n1342 VDD.n1134 4.5005
R90184 VDD.n1340 VDD.n1134 4.5005
R90185 VDD.n1344 VDD.n1134 4.5005
R90186 VDD.n1339 VDD.n1134 4.5005
R90187 VDD.n1345 VDD.n1134 4.5005
R90188 VDD.n1338 VDD.n1134 4.5005
R90189 VDD.n1347 VDD.n1134 4.5005
R90190 VDD.n1337 VDD.n1134 4.5005
R90191 VDD.n1348 VDD.n1134 4.5005
R90192 VDD.n1336 VDD.n1134 4.5005
R90193 VDD.n1350 VDD.n1134 4.5005
R90194 VDD.n1335 VDD.n1134 4.5005
R90195 VDD.n1351 VDD.n1134 4.5005
R90196 VDD.n1334 VDD.n1134 4.5005
R90197 VDD.n1353 VDD.n1134 4.5005
R90198 VDD.n1333 VDD.n1134 4.5005
R90199 VDD.n1354 VDD.n1134 4.5005
R90200 VDD.n1332 VDD.n1134 4.5005
R90201 VDD.n1356 VDD.n1134 4.5005
R90202 VDD.n1331 VDD.n1134 4.5005
R90203 VDD.n1357 VDD.n1134 4.5005
R90204 VDD.n1330 VDD.n1134 4.5005
R90205 VDD.n1359 VDD.n1134 4.5005
R90206 VDD.n1329 VDD.n1134 4.5005
R90207 VDD.n1360 VDD.n1134 4.5005
R90208 VDD.n1328 VDD.n1134 4.5005
R90209 VDD.n1362 VDD.n1134 4.5005
R90210 VDD.n1327 VDD.n1134 4.5005
R90211 VDD.n1363 VDD.n1134 4.5005
R90212 VDD.n1326 VDD.n1134 4.5005
R90213 VDD.n1365 VDD.n1134 4.5005
R90214 VDD.n1325 VDD.n1134 4.5005
R90215 VDD.n1366 VDD.n1134 4.5005
R90216 VDD.n1324 VDD.n1134 4.5005
R90217 VDD.n1368 VDD.n1134 4.5005
R90218 VDD.n1323 VDD.n1134 4.5005
R90219 VDD.n1369 VDD.n1134 4.5005
R90220 VDD.n1322 VDD.n1134 4.5005
R90221 VDD.n1371 VDD.n1134 4.5005
R90222 VDD.n1321 VDD.n1134 4.5005
R90223 VDD.n1372 VDD.n1134 4.5005
R90224 VDD.n1320 VDD.n1134 4.5005
R90225 VDD.n1374 VDD.n1134 4.5005
R90226 VDD.n1319 VDD.n1134 4.5005
R90227 VDD.n1375 VDD.n1134 4.5005
R90228 VDD.n1318 VDD.n1134 4.5005
R90229 VDD.n1376 VDD.n1134 4.5005
R90230 VDD.n1316 VDD.n1134 4.5005
R90231 VDD.n1377 VDD.n1134 4.5005
R90232 VDD.n1315 VDD.n1134 4.5005
R90233 VDD.n1378 VDD.n1134 4.5005
R90234 VDD.n1313 VDD.n1134 4.5005
R90235 VDD.n1379 VDD.n1134 4.5005
R90236 VDD.n1312 VDD.n1134 4.5005
R90237 VDD.n1380 VDD.n1134 4.5005
R90238 VDD.n1310 VDD.n1134 4.5005
R90239 VDD.n1381 VDD.n1134 4.5005
R90240 VDD.n1309 VDD.n1134 4.5005
R90241 VDD.n1382 VDD.n1134 4.5005
R90242 VDD.n1307 VDD.n1134 4.5005
R90243 VDD.n1383 VDD.n1134 4.5005
R90244 VDD.n1306 VDD.n1134 4.5005
R90245 VDD.n1384 VDD.n1134 4.5005
R90246 VDD.n1304 VDD.n1134 4.5005
R90247 VDD.n1385 VDD.n1134 4.5005
R90248 VDD.n1303 VDD.n1134 4.5005
R90249 VDD.n1386 VDD.n1134 4.5005
R90250 VDD.n1301 VDD.n1134 4.5005
R90251 VDD.n1387 VDD.n1134 4.5005
R90252 VDD.n1300 VDD.n1134 4.5005
R90253 VDD.n1388 VDD.n1134 4.5005
R90254 VDD.n1298 VDD.n1134 4.5005
R90255 VDD.n1389 VDD.n1134 4.5005
R90256 VDD.n1297 VDD.n1134 4.5005
R90257 VDD.n1390 VDD.n1134 4.5005
R90258 VDD.n1295 VDD.n1134 4.5005
R90259 VDD.n1391 VDD.n1134 4.5005
R90260 VDD.n1294 VDD.n1134 4.5005
R90261 VDD.n1392 VDD.n1134 4.5005
R90262 VDD.n1292 VDD.n1134 4.5005
R90263 VDD.n1393 VDD.n1134 4.5005
R90264 VDD.n1291 VDD.n1134 4.5005
R90265 VDD.n1394 VDD.n1134 4.5005
R90266 VDD.n1289 VDD.n1134 4.5005
R90267 VDD.n1395 VDD.n1134 4.5005
R90268 VDD.n1288 VDD.n1134 4.5005
R90269 VDD.n1396 VDD.n1134 4.5005
R90270 VDD.n1286 VDD.n1134 4.5005
R90271 VDD.n1397 VDD.n1134 4.5005
R90272 VDD.n1285 VDD.n1134 4.5005
R90273 VDD.n1398 VDD.n1134 4.5005
R90274 VDD.n1283 VDD.n1134 4.5005
R90275 VDD.n1399 VDD.n1134 4.5005
R90276 VDD.n1282 VDD.n1134 4.5005
R90277 VDD.n1400 VDD.n1134 4.5005
R90278 VDD.n1280 VDD.n1134 4.5005
R90279 VDD.n1401 VDD.n1134 4.5005
R90280 VDD.n1279 VDD.n1134 4.5005
R90281 VDD.n1402 VDD.n1134 4.5005
R90282 VDD.n1277 VDD.n1134 4.5005
R90283 VDD.n1403 VDD.n1134 4.5005
R90284 VDD.n1276 VDD.n1134 4.5005
R90285 VDD.n1404 VDD.n1134 4.5005
R90286 VDD.n1274 VDD.n1134 4.5005
R90287 VDD.n1405 VDD.n1134 4.5005
R90288 VDD.n1273 VDD.n1134 4.5005
R90289 VDD.n1406 VDD.n1134 4.5005
R90290 VDD.n1271 VDD.n1134 4.5005
R90291 VDD.n1407 VDD.n1134 4.5005
R90292 VDD.n1270 VDD.n1134 4.5005
R90293 VDD.n1408 VDD.n1134 4.5005
R90294 VDD.n1268 VDD.n1134 4.5005
R90295 VDD.n1409 VDD.n1134 4.5005
R90296 VDD.n1267 VDD.n1134 4.5005
R90297 VDD.n1410 VDD.n1134 4.5005
R90298 VDD.n1265 VDD.n1134 4.5005
R90299 VDD.n1411 VDD.n1134 4.5005
R90300 VDD.n1264 VDD.n1134 4.5005
R90301 VDD.n1412 VDD.n1134 4.5005
R90302 VDD.n1262 VDD.n1134 4.5005
R90303 VDD.n1413 VDD.n1134 4.5005
R90304 VDD.n1261 VDD.n1134 4.5005
R90305 VDD.n1414 VDD.n1134 4.5005
R90306 VDD.n1415 VDD.n1134 4.5005
R90307 VDD.n1674 VDD.n1134 4.5005
R90308 VDD.n1676 VDD.n1256 4.5005
R90309 VDD.n1341 VDD.n1256 4.5005
R90310 VDD.n1342 VDD.n1256 4.5005
R90311 VDD.n1340 VDD.n1256 4.5005
R90312 VDD.n1344 VDD.n1256 4.5005
R90313 VDD.n1339 VDD.n1256 4.5005
R90314 VDD.n1345 VDD.n1256 4.5005
R90315 VDD.n1338 VDD.n1256 4.5005
R90316 VDD.n1347 VDD.n1256 4.5005
R90317 VDD.n1337 VDD.n1256 4.5005
R90318 VDD.n1348 VDD.n1256 4.5005
R90319 VDD.n1336 VDD.n1256 4.5005
R90320 VDD.n1350 VDD.n1256 4.5005
R90321 VDD.n1335 VDD.n1256 4.5005
R90322 VDD.n1351 VDD.n1256 4.5005
R90323 VDD.n1334 VDD.n1256 4.5005
R90324 VDD.n1353 VDD.n1256 4.5005
R90325 VDD.n1333 VDD.n1256 4.5005
R90326 VDD.n1354 VDD.n1256 4.5005
R90327 VDD.n1332 VDD.n1256 4.5005
R90328 VDD.n1356 VDD.n1256 4.5005
R90329 VDD.n1331 VDD.n1256 4.5005
R90330 VDD.n1357 VDD.n1256 4.5005
R90331 VDD.n1330 VDD.n1256 4.5005
R90332 VDD.n1359 VDD.n1256 4.5005
R90333 VDD.n1329 VDD.n1256 4.5005
R90334 VDD.n1360 VDD.n1256 4.5005
R90335 VDD.n1328 VDD.n1256 4.5005
R90336 VDD.n1362 VDD.n1256 4.5005
R90337 VDD.n1327 VDD.n1256 4.5005
R90338 VDD.n1363 VDD.n1256 4.5005
R90339 VDD.n1326 VDD.n1256 4.5005
R90340 VDD.n1365 VDD.n1256 4.5005
R90341 VDD.n1325 VDD.n1256 4.5005
R90342 VDD.n1366 VDD.n1256 4.5005
R90343 VDD.n1324 VDD.n1256 4.5005
R90344 VDD.n1368 VDD.n1256 4.5005
R90345 VDD.n1323 VDD.n1256 4.5005
R90346 VDD.n1369 VDD.n1256 4.5005
R90347 VDD.n1322 VDD.n1256 4.5005
R90348 VDD.n1371 VDD.n1256 4.5005
R90349 VDD.n1321 VDD.n1256 4.5005
R90350 VDD.n1372 VDD.n1256 4.5005
R90351 VDD.n1320 VDD.n1256 4.5005
R90352 VDD.n1374 VDD.n1256 4.5005
R90353 VDD.n1319 VDD.n1256 4.5005
R90354 VDD.n1375 VDD.n1256 4.5005
R90355 VDD.n1318 VDD.n1256 4.5005
R90356 VDD.n1376 VDD.n1256 4.5005
R90357 VDD.n1316 VDD.n1256 4.5005
R90358 VDD.n1377 VDD.n1256 4.5005
R90359 VDD.n1315 VDD.n1256 4.5005
R90360 VDD.n1378 VDD.n1256 4.5005
R90361 VDD.n1313 VDD.n1256 4.5005
R90362 VDD.n1379 VDD.n1256 4.5005
R90363 VDD.n1312 VDD.n1256 4.5005
R90364 VDD.n1380 VDD.n1256 4.5005
R90365 VDD.n1310 VDD.n1256 4.5005
R90366 VDD.n1381 VDD.n1256 4.5005
R90367 VDD.n1309 VDD.n1256 4.5005
R90368 VDD.n1382 VDD.n1256 4.5005
R90369 VDD.n1307 VDD.n1256 4.5005
R90370 VDD.n1383 VDD.n1256 4.5005
R90371 VDD.n1306 VDD.n1256 4.5005
R90372 VDD.n1384 VDD.n1256 4.5005
R90373 VDD.n1304 VDD.n1256 4.5005
R90374 VDD.n1385 VDD.n1256 4.5005
R90375 VDD.n1303 VDD.n1256 4.5005
R90376 VDD.n1386 VDD.n1256 4.5005
R90377 VDD.n1301 VDD.n1256 4.5005
R90378 VDD.n1387 VDD.n1256 4.5005
R90379 VDD.n1300 VDD.n1256 4.5005
R90380 VDD.n1388 VDD.n1256 4.5005
R90381 VDD.n1298 VDD.n1256 4.5005
R90382 VDD.n1389 VDD.n1256 4.5005
R90383 VDD.n1297 VDD.n1256 4.5005
R90384 VDD.n1390 VDD.n1256 4.5005
R90385 VDD.n1295 VDD.n1256 4.5005
R90386 VDD.n1391 VDD.n1256 4.5005
R90387 VDD.n1294 VDD.n1256 4.5005
R90388 VDD.n1392 VDD.n1256 4.5005
R90389 VDD.n1292 VDD.n1256 4.5005
R90390 VDD.n1393 VDD.n1256 4.5005
R90391 VDD.n1291 VDD.n1256 4.5005
R90392 VDD.n1394 VDD.n1256 4.5005
R90393 VDD.n1289 VDD.n1256 4.5005
R90394 VDD.n1395 VDD.n1256 4.5005
R90395 VDD.n1288 VDD.n1256 4.5005
R90396 VDD.n1396 VDD.n1256 4.5005
R90397 VDD.n1286 VDD.n1256 4.5005
R90398 VDD.n1397 VDD.n1256 4.5005
R90399 VDD.n1285 VDD.n1256 4.5005
R90400 VDD.n1398 VDD.n1256 4.5005
R90401 VDD.n1283 VDD.n1256 4.5005
R90402 VDD.n1399 VDD.n1256 4.5005
R90403 VDD.n1282 VDD.n1256 4.5005
R90404 VDD.n1400 VDD.n1256 4.5005
R90405 VDD.n1280 VDD.n1256 4.5005
R90406 VDD.n1401 VDD.n1256 4.5005
R90407 VDD.n1279 VDD.n1256 4.5005
R90408 VDD.n1402 VDD.n1256 4.5005
R90409 VDD.n1277 VDD.n1256 4.5005
R90410 VDD.n1403 VDD.n1256 4.5005
R90411 VDD.n1276 VDD.n1256 4.5005
R90412 VDD.n1404 VDD.n1256 4.5005
R90413 VDD.n1274 VDD.n1256 4.5005
R90414 VDD.n1405 VDD.n1256 4.5005
R90415 VDD.n1273 VDD.n1256 4.5005
R90416 VDD.n1406 VDD.n1256 4.5005
R90417 VDD.n1271 VDD.n1256 4.5005
R90418 VDD.n1407 VDD.n1256 4.5005
R90419 VDD.n1270 VDD.n1256 4.5005
R90420 VDD.n1408 VDD.n1256 4.5005
R90421 VDD.n1268 VDD.n1256 4.5005
R90422 VDD.n1409 VDD.n1256 4.5005
R90423 VDD.n1267 VDD.n1256 4.5005
R90424 VDD.n1410 VDD.n1256 4.5005
R90425 VDD.n1265 VDD.n1256 4.5005
R90426 VDD.n1411 VDD.n1256 4.5005
R90427 VDD.n1264 VDD.n1256 4.5005
R90428 VDD.n1412 VDD.n1256 4.5005
R90429 VDD.n1262 VDD.n1256 4.5005
R90430 VDD.n1413 VDD.n1256 4.5005
R90431 VDD.n1261 VDD.n1256 4.5005
R90432 VDD.n1414 VDD.n1256 4.5005
R90433 VDD.n1415 VDD.n1256 4.5005
R90434 VDD.n1674 VDD.n1256 4.5005
R90435 VDD.n1676 VDD.n1133 4.5005
R90436 VDD.n1341 VDD.n1133 4.5005
R90437 VDD.n1342 VDD.n1133 4.5005
R90438 VDD.n1340 VDD.n1133 4.5005
R90439 VDD.n1344 VDD.n1133 4.5005
R90440 VDD.n1339 VDD.n1133 4.5005
R90441 VDD.n1345 VDD.n1133 4.5005
R90442 VDD.n1338 VDD.n1133 4.5005
R90443 VDD.n1347 VDD.n1133 4.5005
R90444 VDD.n1337 VDD.n1133 4.5005
R90445 VDD.n1348 VDD.n1133 4.5005
R90446 VDD.n1336 VDD.n1133 4.5005
R90447 VDD.n1350 VDD.n1133 4.5005
R90448 VDD.n1335 VDD.n1133 4.5005
R90449 VDD.n1351 VDD.n1133 4.5005
R90450 VDD.n1334 VDD.n1133 4.5005
R90451 VDD.n1353 VDD.n1133 4.5005
R90452 VDD.n1333 VDD.n1133 4.5005
R90453 VDD.n1354 VDD.n1133 4.5005
R90454 VDD.n1332 VDD.n1133 4.5005
R90455 VDD.n1356 VDD.n1133 4.5005
R90456 VDD.n1331 VDD.n1133 4.5005
R90457 VDD.n1357 VDD.n1133 4.5005
R90458 VDD.n1330 VDD.n1133 4.5005
R90459 VDD.n1359 VDD.n1133 4.5005
R90460 VDD.n1329 VDD.n1133 4.5005
R90461 VDD.n1360 VDD.n1133 4.5005
R90462 VDD.n1328 VDD.n1133 4.5005
R90463 VDD.n1362 VDD.n1133 4.5005
R90464 VDD.n1327 VDD.n1133 4.5005
R90465 VDD.n1363 VDD.n1133 4.5005
R90466 VDD.n1326 VDD.n1133 4.5005
R90467 VDD.n1365 VDD.n1133 4.5005
R90468 VDD.n1325 VDD.n1133 4.5005
R90469 VDD.n1366 VDD.n1133 4.5005
R90470 VDD.n1324 VDD.n1133 4.5005
R90471 VDD.n1368 VDD.n1133 4.5005
R90472 VDD.n1323 VDD.n1133 4.5005
R90473 VDD.n1369 VDD.n1133 4.5005
R90474 VDD.n1322 VDD.n1133 4.5005
R90475 VDD.n1371 VDD.n1133 4.5005
R90476 VDD.n1321 VDD.n1133 4.5005
R90477 VDD.n1372 VDD.n1133 4.5005
R90478 VDD.n1320 VDD.n1133 4.5005
R90479 VDD.n1374 VDD.n1133 4.5005
R90480 VDD.n1319 VDD.n1133 4.5005
R90481 VDD.n1375 VDD.n1133 4.5005
R90482 VDD.n1318 VDD.n1133 4.5005
R90483 VDD.n1376 VDD.n1133 4.5005
R90484 VDD.n1316 VDD.n1133 4.5005
R90485 VDD.n1377 VDD.n1133 4.5005
R90486 VDD.n1315 VDD.n1133 4.5005
R90487 VDD.n1378 VDD.n1133 4.5005
R90488 VDD.n1313 VDD.n1133 4.5005
R90489 VDD.n1379 VDD.n1133 4.5005
R90490 VDD.n1312 VDD.n1133 4.5005
R90491 VDD.n1380 VDD.n1133 4.5005
R90492 VDD.n1310 VDD.n1133 4.5005
R90493 VDD.n1381 VDD.n1133 4.5005
R90494 VDD.n1309 VDD.n1133 4.5005
R90495 VDD.n1382 VDD.n1133 4.5005
R90496 VDD.n1307 VDD.n1133 4.5005
R90497 VDD.n1383 VDD.n1133 4.5005
R90498 VDD.n1306 VDD.n1133 4.5005
R90499 VDD.n1384 VDD.n1133 4.5005
R90500 VDD.n1304 VDD.n1133 4.5005
R90501 VDD.n1385 VDD.n1133 4.5005
R90502 VDD.n1303 VDD.n1133 4.5005
R90503 VDD.n1386 VDD.n1133 4.5005
R90504 VDD.n1301 VDD.n1133 4.5005
R90505 VDD.n1387 VDD.n1133 4.5005
R90506 VDD.n1300 VDD.n1133 4.5005
R90507 VDD.n1388 VDD.n1133 4.5005
R90508 VDD.n1298 VDD.n1133 4.5005
R90509 VDD.n1389 VDD.n1133 4.5005
R90510 VDD.n1297 VDD.n1133 4.5005
R90511 VDD.n1390 VDD.n1133 4.5005
R90512 VDD.n1295 VDD.n1133 4.5005
R90513 VDD.n1391 VDD.n1133 4.5005
R90514 VDD.n1294 VDD.n1133 4.5005
R90515 VDD.n1392 VDD.n1133 4.5005
R90516 VDD.n1292 VDD.n1133 4.5005
R90517 VDD.n1393 VDD.n1133 4.5005
R90518 VDD.n1291 VDD.n1133 4.5005
R90519 VDD.n1394 VDD.n1133 4.5005
R90520 VDD.n1289 VDD.n1133 4.5005
R90521 VDD.n1395 VDD.n1133 4.5005
R90522 VDD.n1288 VDD.n1133 4.5005
R90523 VDD.n1396 VDD.n1133 4.5005
R90524 VDD.n1286 VDD.n1133 4.5005
R90525 VDD.n1397 VDD.n1133 4.5005
R90526 VDD.n1285 VDD.n1133 4.5005
R90527 VDD.n1398 VDD.n1133 4.5005
R90528 VDD.n1283 VDD.n1133 4.5005
R90529 VDD.n1399 VDD.n1133 4.5005
R90530 VDD.n1282 VDD.n1133 4.5005
R90531 VDD.n1400 VDD.n1133 4.5005
R90532 VDD.n1280 VDD.n1133 4.5005
R90533 VDD.n1401 VDD.n1133 4.5005
R90534 VDD.n1279 VDD.n1133 4.5005
R90535 VDD.n1402 VDD.n1133 4.5005
R90536 VDD.n1277 VDD.n1133 4.5005
R90537 VDD.n1403 VDD.n1133 4.5005
R90538 VDD.n1276 VDD.n1133 4.5005
R90539 VDD.n1404 VDD.n1133 4.5005
R90540 VDD.n1274 VDD.n1133 4.5005
R90541 VDD.n1405 VDD.n1133 4.5005
R90542 VDD.n1273 VDD.n1133 4.5005
R90543 VDD.n1406 VDD.n1133 4.5005
R90544 VDD.n1271 VDD.n1133 4.5005
R90545 VDD.n1407 VDD.n1133 4.5005
R90546 VDD.n1270 VDD.n1133 4.5005
R90547 VDD.n1408 VDD.n1133 4.5005
R90548 VDD.n1268 VDD.n1133 4.5005
R90549 VDD.n1409 VDD.n1133 4.5005
R90550 VDD.n1267 VDD.n1133 4.5005
R90551 VDD.n1410 VDD.n1133 4.5005
R90552 VDD.n1265 VDD.n1133 4.5005
R90553 VDD.n1411 VDD.n1133 4.5005
R90554 VDD.n1264 VDD.n1133 4.5005
R90555 VDD.n1412 VDD.n1133 4.5005
R90556 VDD.n1262 VDD.n1133 4.5005
R90557 VDD.n1413 VDD.n1133 4.5005
R90558 VDD.n1261 VDD.n1133 4.5005
R90559 VDD.n1414 VDD.n1133 4.5005
R90560 VDD.n1415 VDD.n1133 4.5005
R90561 VDD.n1674 VDD.n1133 4.5005
R90562 VDD.n1676 VDD.n1257 4.5005
R90563 VDD.n1341 VDD.n1257 4.5005
R90564 VDD.n1342 VDD.n1257 4.5005
R90565 VDD.n1340 VDD.n1257 4.5005
R90566 VDD.n1344 VDD.n1257 4.5005
R90567 VDD.n1339 VDD.n1257 4.5005
R90568 VDD.n1345 VDD.n1257 4.5005
R90569 VDD.n1338 VDD.n1257 4.5005
R90570 VDD.n1347 VDD.n1257 4.5005
R90571 VDD.n1337 VDD.n1257 4.5005
R90572 VDD.n1348 VDD.n1257 4.5005
R90573 VDD.n1336 VDD.n1257 4.5005
R90574 VDD.n1350 VDD.n1257 4.5005
R90575 VDD.n1335 VDD.n1257 4.5005
R90576 VDD.n1351 VDD.n1257 4.5005
R90577 VDD.n1334 VDD.n1257 4.5005
R90578 VDD.n1353 VDD.n1257 4.5005
R90579 VDD.n1333 VDD.n1257 4.5005
R90580 VDD.n1354 VDD.n1257 4.5005
R90581 VDD.n1332 VDD.n1257 4.5005
R90582 VDD.n1356 VDD.n1257 4.5005
R90583 VDD.n1331 VDD.n1257 4.5005
R90584 VDD.n1357 VDD.n1257 4.5005
R90585 VDD.n1330 VDD.n1257 4.5005
R90586 VDD.n1359 VDD.n1257 4.5005
R90587 VDD.n1329 VDD.n1257 4.5005
R90588 VDD.n1360 VDD.n1257 4.5005
R90589 VDD.n1328 VDD.n1257 4.5005
R90590 VDD.n1362 VDD.n1257 4.5005
R90591 VDD.n1327 VDD.n1257 4.5005
R90592 VDD.n1363 VDD.n1257 4.5005
R90593 VDD.n1326 VDD.n1257 4.5005
R90594 VDD.n1365 VDD.n1257 4.5005
R90595 VDD.n1325 VDD.n1257 4.5005
R90596 VDD.n1366 VDD.n1257 4.5005
R90597 VDD.n1324 VDD.n1257 4.5005
R90598 VDD.n1368 VDD.n1257 4.5005
R90599 VDD.n1323 VDD.n1257 4.5005
R90600 VDD.n1369 VDD.n1257 4.5005
R90601 VDD.n1322 VDD.n1257 4.5005
R90602 VDD.n1371 VDD.n1257 4.5005
R90603 VDD.n1321 VDD.n1257 4.5005
R90604 VDD.n1372 VDD.n1257 4.5005
R90605 VDD.n1320 VDD.n1257 4.5005
R90606 VDD.n1374 VDD.n1257 4.5005
R90607 VDD.n1319 VDD.n1257 4.5005
R90608 VDD.n1375 VDD.n1257 4.5005
R90609 VDD.n1318 VDD.n1257 4.5005
R90610 VDD.n1376 VDD.n1257 4.5005
R90611 VDD.n1316 VDD.n1257 4.5005
R90612 VDD.n1377 VDD.n1257 4.5005
R90613 VDD.n1315 VDD.n1257 4.5005
R90614 VDD.n1378 VDD.n1257 4.5005
R90615 VDD.n1313 VDD.n1257 4.5005
R90616 VDD.n1379 VDD.n1257 4.5005
R90617 VDD.n1312 VDD.n1257 4.5005
R90618 VDD.n1380 VDD.n1257 4.5005
R90619 VDD.n1310 VDD.n1257 4.5005
R90620 VDD.n1381 VDD.n1257 4.5005
R90621 VDD.n1309 VDD.n1257 4.5005
R90622 VDD.n1382 VDD.n1257 4.5005
R90623 VDD.n1307 VDD.n1257 4.5005
R90624 VDD.n1383 VDD.n1257 4.5005
R90625 VDD.n1306 VDD.n1257 4.5005
R90626 VDD.n1384 VDD.n1257 4.5005
R90627 VDD.n1304 VDD.n1257 4.5005
R90628 VDD.n1385 VDD.n1257 4.5005
R90629 VDD.n1303 VDD.n1257 4.5005
R90630 VDD.n1386 VDD.n1257 4.5005
R90631 VDD.n1301 VDD.n1257 4.5005
R90632 VDD.n1387 VDD.n1257 4.5005
R90633 VDD.n1300 VDD.n1257 4.5005
R90634 VDD.n1388 VDD.n1257 4.5005
R90635 VDD.n1298 VDD.n1257 4.5005
R90636 VDD.n1389 VDD.n1257 4.5005
R90637 VDD.n1297 VDD.n1257 4.5005
R90638 VDD.n1390 VDD.n1257 4.5005
R90639 VDD.n1295 VDD.n1257 4.5005
R90640 VDD.n1391 VDD.n1257 4.5005
R90641 VDD.n1294 VDD.n1257 4.5005
R90642 VDD.n1392 VDD.n1257 4.5005
R90643 VDD.n1292 VDD.n1257 4.5005
R90644 VDD.n1393 VDD.n1257 4.5005
R90645 VDD.n1291 VDD.n1257 4.5005
R90646 VDD.n1394 VDD.n1257 4.5005
R90647 VDD.n1289 VDD.n1257 4.5005
R90648 VDD.n1395 VDD.n1257 4.5005
R90649 VDD.n1288 VDD.n1257 4.5005
R90650 VDD.n1396 VDD.n1257 4.5005
R90651 VDD.n1286 VDD.n1257 4.5005
R90652 VDD.n1397 VDD.n1257 4.5005
R90653 VDD.n1285 VDD.n1257 4.5005
R90654 VDD.n1398 VDD.n1257 4.5005
R90655 VDD.n1283 VDD.n1257 4.5005
R90656 VDD.n1399 VDD.n1257 4.5005
R90657 VDD.n1282 VDD.n1257 4.5005
R90658 VDD.n1400 VDD.n1257 4.5005
R90659 VDD.n1280 VDD.n1257 4.5005
R90660 VDD.n1401 VDD.n1257 4.5005
R90661 VDD.n1279 VDD.n1257 4.5005
R90662 VDD.n1402 VDD.n1257 4.5005
R90663 VDD.n1277 VDD.n1257 4.5005
R90664 VDD.n1403 VDD.n1257 4.5005
R90665 VDD.n1276 VDD.n1257 4.5005
R90666 VDD.n1404 VDD.n1257 4.5005
R90667 VDD.n1274 VDD.n1257 4.5005
R90668 VDD.n1405 VDD.n1257 4.5005
R90669 VDD.n1273 VDD.n1257 4.5005
R90670 VDD.n1406 VDD.n1257 4.5005
R90671 VDD.n1271 VDD.n1257 4.5005
R90672 VDD.n1407 VDD.n1257 4.5005
R90673 VDD.n1270 VDD.n1257 4.5005
R90674 VDD.n1408 VDD.n1257 4.5005
R90675 VDD.n1268 VDD.n1257 4.5005
R90676 VDD.n1409 VDD.n1257 4.5005
R90677 VDD.n1267 VDD.n1257 4.5005
R90678 VDD.n1410 VDD.n1257 4.5005
R90679 VDD.n1265 VDD.n1257 4.5005
R90680 VDD.n1411 VDD.n1257 4.5005
R90681 VDD.n1264 VDD.n1257 4.5005
R90682 VDD.n1412 VDD.n1257 4.5005
R90683 VDD.n1262 VDD.n1257 4.5005
R90684 VDD.n1413 VDD.n1257 4.5005
R90685 VDD.n1261 VDD.n1257 4.5005
R90686 VDD.n1414 VDD.n1257 4.5005
R90687 VDD.n1415 VDD.n1257 4.5005
R90688 VDD.n1674 VDD.n1257 4.5005
R90689 VDD.n1676 VDD.n1132 4.5005
R90690 VDD.n1341 VDD.n1132 4.5005
R90691 VDD.n1342 VDD.n1132 4.5005
R90692 VDD.n1340 VDD.n1132 4.5005
R90693 VDD.n1344 VDD.n1132 4.5005
R90694 VDD.n1339 VDD.n1132 4.5005
R90695 VDD.n1345 VDD.n1132 4.5005
R90696 VDD.n1338 VDD.n1132 4.5005
R90697 VDD.n1347 VDD.n1132 4.5005
R90698 VDD.n1337 VDD.n1132 4.5005
R90699 VDD.n1348 VDD.n1132 4.5005
R90700 VDD.n1336 VDD.n1132 4.5005
R90701 VDD.n1350 VDD.n1132 4.5005
R90702 VDD.n1335 VDD.n1132 4.5005
R90703 VDD.n1351 VDD.n1132 4.5005
R90704 VDD.n1334 VDD.n1132 4.5005
R90705 VDD.n1353 VDD.n1132 4.5005
R90706 VDD.n1333 VDD.n1132 4.5005
R90707 VDD.n1354 VDD.n1132 4.5005
R90708 VDD.n1332 VDD.n1132 4.5005
R90709 VDD.n1356 VDD.n1132 4.5005
R90710 VDD.n1331 VDD.n1132 4.5005
R90711 VDD.n1357 VDD.n1132 4.5005
R90712 VDD.n1330 VDD.n1132 4.5005
R90713 VDD.n1359 VDD.n1132 4.5005
R90714 VDD.n1329 VDD.n1132 4.5005
R90715 VDD.n1360 VDD.n1132 4.5005
R90716 VDD.n1328 VDD.n1132 4.5005
R90717 VDD.n1362 VDD.n1132 4.5005
R90718 VDD.n1327 VDD.n1132 4.5005
R90719 VDD.n1363 VDD.n1132 4.5005
R90720 VDD.n1326 VDD.n1132 4.5005
R90721 VDD.n1365 VDD.n1132 4.5005
R90722 VDD.n1325 VDD.n1132 4.5005
R90723 VDD.n1366 VDD.n1132 4.5005
R90724 VDD.n1324 VDD.n1132 4.5005
R90725 VDD.n1368 VDD.n1132 4.5005
R90726 VDD.n1323 VDD.n1132 4.5005
R90727 VDD.n1369 VDD.n1132 4.5005
R90728 VDD.n1322 VDD.n1132 4.5005
R90729 VDD.n1371 VDD.n1132 4.5005
R90730 VDD.n1321 VDD.n1132 4.5005
R90731 VDD.n1372 VDD.n1132 4.5005
R90732 VDD.n1320 VDD.n1132 4.5005
R90733 VDD.n1374 VDD.n1132 4.5005
R90734 VDD.n1319 VDD.n1132 4.5005
R90735 VDD.n1375 VDD.n1132 4.5005
R90736 VDD.n1318 VDD.n1132 4.5005
R90737 VDD.n1376 VDD.n1132 4.5005
R90738 VDD.n1316 VDD.n1132 4.5005
R90739 VDD.n1377 VDD.n1132 4.5005
R90740 VDD.n1315 VDD.n1132 4.5005
R90741 VDD.n1378 VDD.n1132 4.5005
R90742 VDD.n1313 VDD.n1132 4.5005
R90743 VDD.n1379 VDD.n1132 4.5005
R90744 VDD.n1312 VDD.n1132 4.5005
R90745 VDD.n1380 VDD.n1132 4.5005
R90746 VDD.n1310 VDD.n1132 4.5005
R90747 VDD.n1381 VDD.n1132 4.5005
R90748 VDD.n1309 VDD.n1132 4.5005
R90749 VDD.n1382 VDD.n1132 4.5005
R90750 VDD.n1307 VDD.n1132 4.5005
R90751 VDD.n1383 VDD.n1132 4.5005
R90752 VDD.n1306 VDD.n1132 4.5005
R90753 VDD.n1384 VDD.n1132 4.5005
R90754 VDD.n1304 VDD.n1132 4.5005
R90755 VDD.n1385 VDD.n1132 4.5005
R90756 VDD.n1303 VDD.n1132 4.5005
R90757 VDD.n1386 VDD.n1132 4.5005
R90758 VDD.n1301 VDD.n1132 4.5005
R90759 VDD.n1387 VDD.n1132 4.5005
R90760 VDD.n1300 VDD.n1132 4.5005
R90761 VDD.n1388 VDD.n1132 4.5005
R90762 VDD.n1298 VDD.n1132 4.5005
R90763 VDD.n1389 VDD.n1132 4.5005
R90764 VDD.n1297 VDD.n1132 4.5005
R90765 VDD.n1390 VDD.n1132 4.5005
R90766 VDD.n1295 VDD.n1132 4.5005
R90767 VDD.n1391 VDD.n1132 4.5005
R90768 VDD.n1294 VDD.n1132 4.5005
R90769 VDD.n1392 VDD.n1132 4.5005
R90770 VDD.n1292 VDD.n1132 4.5005
R90771 VDD.n1393 VDD.n1132 4.5005
R90772 VDD.n1291 VDD.n1132 4.5005
R90773 VDD.n1394 VDD.n1132 4.5005
R90774 VDD.n1289 VDD.n1132 4.5005
R90775 VDD.n1395 VDD.n1132 4.5005
R90776 VDD.n1288 VDD.n1132 4.5005
R90777 VDD.n1396 VDD.n1132 4.5005
R90778 VDD.n1286 VDD.n1132 4.5005
R90779 VDD.n1397 VDD.n1132 4.5005
R90780 VDD.n1285 VDD.n1132 4.5005
R90781 VDD.n1398 VDD.n1132 4.5005
R90782 VDD.n1283 VDD.n1132 4.5005
R90783 VDD.n1399 VDD.n1132 4.5005
R90784 VDD.n1282 VDD.n1132 4.5005
R90785 VDD.n1400 VDD.n1132 4.5005
R90786 VDD.n1280 VDD.n1132 4.5005
R90787 VDD.n1401 VDD.n1132 4.5005
R90788 VDD.n1279 VDD.n1132 4.5005
R90789 VDD.n1402 VDD.n1132 4.5005
R90790 VDD.n1277 VDD.n1132 4.5005
R90791 VDD.n1403 VDD.n1132 4.5005
R90792 VDD.n1276 VDD.n1132 4.5005
R90793 VDD.n1404 VDD.n1132 4.5005
R90794 VDD.n1274 VDD.n1132 4.5005
R90795 VDD.n1405 VDD.n1132 4.5005
R90796 VDD.n1273 VDD.n1132 4.5005
R90797 VDD.n1406 VDD.n1132 4.5005
R90798 VDD.n1271 VDD.n1132 4.5005
R90799 VDD.n1407 VDD.n1132 4.5005
R90800 VDD.n1270 VDD.n1132 4.5005
R90801 VDD.n1408 VDD.n1132 4.5005
R90802 VDD.n1268 VDD.n1132 4.5005
R90803 VDD.n1409 VDD.n1132 4.5005
R90804 VDD.n1267 VDD.n1132 4.5005
R90805 VDD.n1410 VDD.n1132 4.5005
R90806 VDD.n1265 VDD.n1132 4.5005
R90807 VDD.n1411 VDD.n1132 4.5005
R90808 VDD.n1264 VDD.n1132 4.5005
R90809 VDD.n1412 VDD.n1132 4.5005
R90810 VDD.n1262 VDD.n1132 4.5005
R90811 VDD.n1413 VDD.n1132 4.5005
R90812 VDD.n1261 VDD.n1132 4.5005
R90813 VDD.n1414 VDD.n1132 4.5005
R90814 VDD.n1415 VDD.n1132 4.5005
R90815 VDD.n1674 VDD.n1132 4.5005
R90816 VDD.n1676 VDD.n1675 4.5005
R90817 VDD.n1675 VDD.n1341 4.5005
R90818 VDD.n1675 VDD.n1342 4.5005
R90819 VDD.n1675 VDD.n1340 4.5005
R90820 VDD.n1675 VDD.n1344 4.5005
R90821 VDD.n1675 VDD.n1339 4.5005
R90822 VDD.n1675 VDD.n1345 4.5005
R90823 VDD.n1675 VDD.n1338 4.5005
R90824 VDD.n1675 VDD.n1347 4.5005
R90825 VDD.n1675 VDD.n1337 4.5005
R90826 VDD.n1675 VDD.n1348 4.5005
R90827 VDD.n1675 VDD.n1336 4.5005
R90828 VDD.n1675 VDD.n1350 4.5005
R90829 VDD.n1675 VDD.n1335 4.5005
R90830 VDD.n1675 VDD.n1351 4.5005
R90831 VDD.n1675 VDD.n1334 4.5005
R90832 VDD.n1675 VDD.n1353 4.5005
R90833 VDD.n1675 VDD.n1333 4.5005
R90834 VDD.n1675 VDD.n1354 4.5005
R90835 VDD.n1675 VDD.n1332 4.5005
R90836 VDD.n1675 VDD.n1356 4.5005
R90837 VDD.n1675 VDD.n1331 4.5005
R90838 VDD.n1675 VDD.n1357 4.5005
R90839 VDD.n1675 VDD.n1330 4.5005
R90840 VDD.n1675 VDD.n1359 4.5005
R90841 VDD.n1675 VDD.n1329 4.5005
R90842 VDD.n1675 VDD.n1360 4.5005
R90843 VDD.n1675 VDD.n1328 4.5005
R90844 VDD.n1675 VDD.n1362 4.5005
R90845 VDD.n1675 VDD.n1327 4.5005
R90846 VDD.n1675 VDD.n1363 4.5005
R90847 VDD.n1675 VDD.n1326 4.5005
R90848 VDD.n1675 VDD.n1365 4.5005
R90849 VDD.n1675 VDD.n1325 4.5005
R90850 VDD.n1675 VDD.n1366 4.5005
R90851 VDD.n1675 VDD.n1324 4.5005
R90852 VDD.n1675 VDD.n1368 4.5005
R90853 VDD.n1675 VDD.n1323 4.5005
R90854 VDD.n1675 VDD.n1369 4.5005
R90855 VDD.n1675 VDD.n1322 4.5005
R90856 VDD.n1675 VDD.n1371 4.5005
R90857 VDD.n1675 VDD.n1321 4.5005
R90858 VDD.n1675 VDD.n1372 4.5005
R90859 VDD.n1675 VDD.n1320 4.5005
R90860 VDD.n1675 VDD.n1374 4.5005
R90861 VDD.n1675 VDD.n1319 4.5005
R90862 VDD.n1675 VDD.n1375 4.5005
R90863 VDD.n1675 VDD.n1318 4.5005
R90864 VDD.n1675 VDD.n1376 4.5005
R90865 VDD.n1675 VDD.n1316 4.5005
R90866 VDD.n1675 VDD.n1377 4.5005
R90867 VDD.n1675 VDD.n1315 4.5005
R90868 VDD.n1675 VDD.n1378 4.5005
R90869 VDD.n1675 VDD.n1313 4.5005
R90870 VDD.n1675 VDD.n1379 4.5005
R90871 VDD.n1675 VDD.n1312 4.5005
R90872 VDD.n1675 VDD.n1380 4.5005
R90873 VDD.n1675 VDD.n1310 4.5005
R90874 VDD.n1675 VDD.n1381 4.5005
R90875 VDD.n1675 VDD.n1309 4.5005
R90876 VDD.n1675 VDD.n1382 4.5005
R90877 VDD.n1675 VDD.n1307 4.5005
R90878 VDD.n1675 VDD.n1383 4.5005
R90879 VDD.n1675 VDD.n1306 4.5005
R90880 VDD.n1675 VDD.n1384 4.5005
R90881 VDD.n1675 VDD.n1304 4.5005
R90882 VDD.n1675 VDD.n1385 4.5005
R90883 VDD.n1675 VDD.n1303 4.5005
R90884 VDD.n1675 VDD.n1386 4.5005
R90885 VDD.n1675 VDD.n1301 4.5005
R90886 VDD.n1675 VDD.n1387 4.5005
R90887 VDD.n1675 VDD.n1300 4.5005
R90888 VDD.n1675 VDD.n1388 4.5005
R90889 VDD.n1675 VDD.n1298 4.5005
R90890 VDD.n1675 VDD.n1389 4.5005
R90891 VDD.n1675 VDD.n1297 4.5005
R90892 VDD.n1675 VDD.n1390 4.5005
R90893 VDD.n1675 VDD.n1295 4.5005
R90894 VDD.n1675 VDD.n1391 4.5005
R90895 VDD.n1675 VDD.n1294 4.5005
R90896 VDD.n1675 VDD.n1392 4.5005
R90897 VDD.n1675 VDD.n1292 4.5005
R90898 VDD.n1675 VDD.n1393 4.5005
R90899 VDD.n1675 VDD.n1291 4.5005
R90900 VDD.n1675 VDD.n1394 4.5005
R90901 VDD.n1675 VDD.n1289 4.5005
R90902 VDD.n1675 VDD.n1395 4.5005
R90903 VDD.n1675 VDD.n1288 4.5005
R90904 VDD.n1675 VDD.n1396 4.5005
R90905 VDD.n1675 VDD.n1286 4.5005
R90906 VDD.n1675 VDD.n1397 4.5005
R90907 VDD.n1675 VDD.n1285 4.5005
R90908 VDD.n1675 VDD.n1398 4.5005
R90909 VDD.n1675 VDD.n1283 4.5005
R90910 VDD.n1675 VDD.n1399 4.5005
R90911 VDD.n1675 VDD.n1282 4.5005
R90912 VDD.n1675 VDD.n1400 4.5005
R90913 VDD.n1675 VDD.n1280 4.5005
R90914 VDD.n1675 VDD.n1401 4.5005
R90915 VDD.n1675 VDD.n1279 4.5005
R90916 VDD.n1675 VDD.n1402 4.5005
R90917 VDD.n1675 VDD.n1277 4.5005
R90918 VDD.n1675 VDD.n1403 4.5005
R90919 VDD.n1675 VDD.n1276 4.5005
R90920 VDD.n1675 VDD.n1404 4.5005
R90921 VDD.n1675 VDD.n1274 4.5005
R90922 VDD.n1675 VDD.n1405 4.5005
R90923 VDD.n1675 VDD.n1273 4.5005
R90924 VDD.n1675 VDD.n1406 4.5005
R90925 VDD.n1675 VDD.n1271 4.5005
R90926 VDD.n1675 VDD.n1407 4.5005
R90927 VDD.n1675 VDD.n1270 4.5005
R90928 VDD.n1675 VDD.n1408 4.5005
R90929 VDD.n1675 VDD.n1268 4.5005
R90930 VDD.n1675 VDD.n1409 4.5005
R90931 VDD.n1675 VDD.n1267 4.5005
R90932 VDD.n1675 VDD.n1410 4.5005
R90933 VDD.n1675 VDD.n1265 4.5005
R90934 VDD.n1675 VDD.n1411 4.5005
R90935 VDD.n1675 VDD.n1264 4.5005
R90936 VDD.n1675 VDD.n1412 4.5005
R90937 VDD.n1675 VDD.n1262 4.5005
R90938 VDD.n1675 VDD.n1413 4.5005
R90939 VDD.n1675 VDD.n1261 4.5005
R90940 VDD.n1675 VDD.n1414 4.5005
R90941 VDD.n1675 VDD.n1415 4.5005
R90942 VDD.n1675 VDD.n1674 4.5005
R90943 VDD.n1676 VDD.n1131 4.5005
R90944 VDD.n1341 VDD.n1131 4.5005
R90945 VDD.n1342 VDD.n1131 4.5005
R90946 VDD.n1340 VDD.n1131 4.5005
R90947 VDD.n1344 VDD.n1131 4.5005
R90948 VDD.n1339 VDD.n1131 4.5005
R90949 VDD.n1345 VDD.n1131 4.5005
R90950 VDD.n1338 VDD.n1131 4.5005
R90951 VDD.n1347 VDD.n1131 4.5005
R90952 VDD.n1337 VDD.n1131 4.5005
R90953 VDD.n1348 VDD.n1131 4.5005
R90954 VDD.n1336 VDD.n1131 4.5005
R90955 VDD.n1350 VDD.n1131 4.5005
R90956 VDD.n1335 VDD.n1131 4.5005
R90957 VDD.n1351 VDD.n1131 4.5005
R90958 VDD.n1334 VDD.n1131 4.5005
R90959 VDD.n1353 VDD.n1131 4.5005
R90960 VDD.n1333 VDD.n1131 4.5005
R90961 VDD.n1354 VDD.n1131 4.5005
R90962 VDD.n1332 VDD.n1131 4.5005
R90963 VDD.n1356 VDD.n1131 4.5005
R90964 VDD.n1331 VDD.n1131 4.5005
R90965 VDD.n1357 VDD.n1131 4.5005
R90966 VDD.n1330 VDD.n1131 4.5005
R90967 VDD.n1359 VDD.n1131 4.5005
R90968 VDD.n1329 VDD.n1131 4.5005
R90969 VDD.n1360 VDD.n1131 4.5005
R90970 VDD.n1328 VDD.n1131 4.5005
R90971 VDD.n1362 VDD.n1131 4.5005
R90972 VDD.n1327 VDD.n1131 4.5005
R90973 VDD.n1363 VDD.n1131 4.5005
R90974 VDD.n1326 VDD.n1131 4.5005
R90975 VDD.n1365 VDD.n1131 4.5005
R90976 VDD.n1325 VDD.n1131 4.5005
R90977 VDD.n1366 VDD.n1131 4.5005
R90978 VDD.n1324 VDD.n1131 4.5005
R90979 VDD.n1368 VDD.n1131 4.5005
R90980 VDD.n1323 VDD.n1131 4.5005
R90981 VDD.n1369 VDD.n1131 4.5005
R90982 VDD.n1322 VDD.n1131 4.5005
R90983 VDD.n1371 VDD.n1131 4.5005
R90984 VDD.n1321 VDD.n1131 4.5005
R90985 VDD.n1372 VDD.n1131 4.5005
R90986 VDD.n1320 VDD.n1131 4.5005
R90987 VDD.n1374 VDD.n1131 4.5005
R90988 VDD.n1319 VDD.n1131 4.5005
R90989 VDD.n1375 VDD.n1131 4.5005
R90990 VDD.n1318 VDD.n1131 4.5005
R90991 VDD.n1376 VDD.n1131 4.5005
R90992 VDD.n1316 VDD.n1131 4.5005
R90993 VDD.n1377 VDD.n1131 4.5005
R90994 VDD.n1315 VDD.n1131 4.5005
R90995 VDD.n1378 VDD.n1131 4.5005
R90996 VDD.n1313 VDD.n1131 4.5005
R90997 VDD.n1379 VDD.n1131 4.5005
R90998 VDD.n1312 VDD.n1131 4.5005
R90999 VDD.n1380 VDD.n1131 4.5005
R91000 VDD.n1310 VDD.n1131 4.5005
R91001 VDD.n1381 VDD.n1131 4.5005
R91002 VDD.n1309 VDD.n1131 4.5005
R91003 VDD.n1382 VDD.n1131 4.5005
R91004 VDD.n1307 VDD.n1131 4.5005
R91005 VDD.n1383 VDD.n1131 4.5005
R91006 VDD.n1306 VDD.n1131 4.5005
R91007 VDD.n1384 VDD.n1131 4.5005
R91008 VDD.n1304 VDD.n1131 4.5005
R91009 VDD.n1385 VDD.n1131 4.5005
R91010 VDD.n1303 VDD.n1131 4.5005
R91011 VDD.n1386 VDD.n1131 4.5005
R91012 VDD.n1301 VDD.n1131 4.5005
R91013 VDD.n1387 VDD.n1131 4.5005
R91014 VDD.n1300 VDD.n1131 4.5005
R91015 VDD.n1388 VDD.n1131 4.5005
R91016 VDD.n1298 VDD.n1131 4.5005
R91017 VDD.n1389 VDD.n1131 4.5005
R91018 VDD.n1297 VDD.n1131 4.5005
R91019 VDD.n1390 VDD.n1131 4.5005
R91020 VDD.n1295 VDD.n1131 4.5005
R91021 VDD.n1391 VDD.n1131 4.5005
R91022 VDD.n1294 VDD.n1131 4.5005
R91023 VDD.n1392 VDD.n1131 4.5005
R91024 VDD.n1292 VDD.n1131 4.5005
R91025 VDD.n1393 VDD.n1131 4.5005
R91026 VDD.n1291 VDD.n1131 4.5005
R91027 VDD.n1394 VDD.n1131 4.5005
R91028 VDD.n1289 VDD.n1131 4.5005
R91029 VDD.n1395 VDD.n1131 4.5005
R91030 VDD.n1288 VDD.n1131 4.5005
R91031 VDD.n1396 VDD.n1131 4.5005
R91032 VDD.n1286 VDD.n1131 4.5005
R91033 VDD.n1397 VDD.n1131 4.5005
R91034 VDD.n1285 VDD.n1131 4.5005
R91035 VDD.n1398 VDD.n1131 4.5005
R91036 VDD.n1283 VDD.n1131 4.5005
R91037 VDD.n1399 VDD.n1131 4.5005
R91038 VDD.n1282 VDD.n1131 4.5005
R91039 VDD.n1400 VDD.n1131 4.5005
R91040 VDD.n1280 VDD.n1131 4.5005
R91041 VDD.n1401 VDD.n1131 4.5005
R91042 VDD.n1279 VDD.n1131 4.5005
R91043 VDD.n1402 VDD.n1131 4.5005
R91044 VDD.n1277 VDD.n1131 4.5005
R91045 VDD.n1403 VDD.n1131 4.5005
R91046 VDD.n1276 VDD.n1131 4.5005
R91047 VDD.n1404 VDD.n1131 4.5005
R91048 VDD.n1274 VDD.n1131 4.5005
R91049 VDD.n1405 VDD.n1131 4.5005
R91050 VDD.n1273 VDD.n1131 4.5005
R91051 VDD.n1406 VDD.n1131 4.5005
R91052 VDD.n1271 VDD.n1131 4.5005
R91053 VDD.n1407 VDD.n1131 4.5005
R91054 VDD.n1270 VDD.n1131 4.5005
R91055 VDD.n1408 VDD.n1131 4.5005
R91056 VDD.n1268 VDD.n1131 4.5005
R91057 VDD.n1409 VDD.n1131 4.5005
R91058 VDD.n1267 VDD.n1131 4.5005
R91059 VDD.n1410 VDD.n1131 4.5005
R91060 VDD.n1265 VDD.n1131 4.5005
R91061 VDD.n1411 VDD.n1131 4.5005
R91062 VDD.n1264 VDD.n1131 4.5005
R91063 VDD.n1412 VDD.n1131 4.5005
R91064 VDD.n1262 VDD.n1131 4.5005
R91065 VDD.n1413 VDD.n1131 4.5005
R91066 VDD.n1261 VDD.n1131 4.5005
R91067 VDD.n1414 VDD.n1131 4.5005
R91068 VDD.n1544 VDD.n1131 4.5005
R91069 VDD.n1415 VDD.n1131 4.5005
R91070 VDD.n1674 VDD.n1131 4.5005
R91071 VDD.n1676 VDD.n1195 2.25083
R91072 VDD.n1480 VDD.n1479 2.25083
R91073 VDD.n1480 VDD.n1478 2.25083
R91074 VDD.n1480 VDD.n1477 2.25083
R91075 VDD.n1480 VDD.n1476 2.25083
R91076 VDD.n1480 VDD.n1475 2.25083
R91077 VDD.n1480 VDD.n1474 2.25083
R91078 VDD.n1480 VDD.n1473 2.25083
R91079 VDD.n1480 VDD.n1472 2.25083
R91080 VDD.n1480 VDD.n1471 2.25083
R91081 VDD.n1480 VDD.n1470 2.25083
R91082 VDD.n1480 VDD.n1469 2.25083
R91083 VDD.n1480 VDD.n1468 2.25083
R91084 VDD.n1480 VDD.n1467 2.25083
R91085 VDD.n1480 VDD.n1466 2.25083
R91086 VDD.n1480 VDD.n1465 2.25083
R91087 VDD.n1480 VDD.n1464 2.25083
R91088 VDD.n1480 VDD.n1463 2.25083
R91089 VDD.n1480 VDD.n1462 2.25083
R91090 VDD.n1480 VDD.n1461 2.25083
R91091 VDD.n1480 VDD.n1460 2.25083
R91092 VDD.n1480 VDD.n1459 2.25083
R91093 VDD.n1480 VDD.n1458 2.25083
R91094 VDD.n1480 VDD.n1457 2.25083
R91095 VDD.n1480 VDD.n1456 2.25083
R91096 VDD.n1480 VDD.n1455 2.25083
R91097 VDD.n1480 VDD.n1454 2.25083
R91098 VDD.n1480 VDD.n1453 2.25083
R91099 VDD.n1480 VDD.n1452 2.25083
R91100 VDD.n1480 VDD.n1451 2.25083
R91101 VDD.n1480 VDD.n1450 2.25083
R91102 VDD.n1480 VDD.n1449 2.25083
R91103 VDD.n1480 VDD.n1448 2.25083
R91104 VDD.n1480 VDD.n1447 2.25083
R91105 VDD.n1480 VDD.n1446 2.25083
R91106 VDD.n1480 VDD.n1445 2.25083
R91107 VDD.n1480 VDD.n1444 2.25083
R91108 VDD.n1480 VDD.n1443 2.25083
R91109 VDD.n1480 VDD.n1442 2.25083
R91110 VDD.n1480 VDD.n1441 2.25083
R91111 VDD.n1480 VDD.n1440 2.25083
R91112 VDD.n1480 VDD.n1439 2.25083
R91113 VDD.n1480 VDD.n1438 2.25083
R91114 VDD.n1480 VDD.n1437 2.25083
R91115 VDD.n1480 VDD.n1436 2.25083
R91116 VDD.n1480 VDD.n1435 2.25083
R91117 VDD.n1480 VDD.n1434 2.25083
R91118 VDD.n1480 VDD.n1433 2.25083
R91119 VDD.n1480 VDD.n1432 2.25083
R91120 VDD.n1480 VDD.n1431 2.25083
R91121 VDD.n1480 VDD.n1430 2.25083
R91122 VDD.n1480 VDD.n1429 2.25083
R91123 VDD.n1480 VDD.n1428 2.25083
R91124 VDD.n1480 VDD.n1427 2.25083
R91125 VDD.n1480 VDD.n1426 2.25083
R91126 VDD.n1480 VDD.n1425 2.25083
R91127 VDD.n1480 VDD.n1424 2.25083
R91128 VDD.n1480 VDD.n1423 2.25083
R91129 VDD.n1480 VDD.n1422 2.25083
R91130 VDD.n1480 VDD.n1421 2.25083
R91131 VDD.n1480 VDD.n1420 2.25083
R91132 VDD.n1480 VDD.n1419 2.25083
R91133 VDD.n1480 VDD.n1418 2.25083
R91134 VDD.n1481 VDD.n1480 2.25083
R91135 VDD.n1480 VDD.n1417 2.25083
R91136 VDD.n1607 VDD.n1606 2.25083
R91137 VDD.n1607 VDD.n1605 2.25083
R91138 VDD.n1607 VDD.n1604 2.25083
R91139 VDD.n1607 VDD.n1603 2.25083
R91140 VDD.n1607 VDD.n1602 2.25083
R91141 VDD.n1607 VDD.n1601 2.25083
R91142 VDD.n1607 VDD.n1600 2.25083
R91143 VDD.n1607 VDD.n1599 2.25083
R91144 VDD.n1607 VDD.n1598 2.25083
R91145 VDD.n1607 VDD.n1597 2.25083
R91146 VDD.n1607 VDD.n1596 2.25083
R91147 VDD.n1607 VDD.n1595 2.25083
R91148 VDD.n1607 VDD.n1594 2.25083
R91149 VDD.n1607 VDD.n1593 2.25083
R91150 VDD.n1607 VDD.n1592 2.25083
R91151 VDD.n1607 VDD.n1591 2.25083
R91152 VDD.n1607 VDD.n1590 2.25083
R91153 VDD.n1607 VDD.n1589 2.25083
R91154 VDD.n1607 VDD.n1588 2.25083
R91155 VDD.n1607 VDD.n1587 2.25083
R91156 VDD.n1607 VDD.n1586 2.25083
R91157 VDD.n1607 VDD.n1585 2.25083
R91158 VDD.n1607 VDD.n1584 2.25083
R91159 VDD.n1607 VDD.n1583 2.25083
R91160 VDD.n1607 VDD.n1582 2.25083
R91161 VDD.n1607 VDD.n1581 2.25083
R91162 VDD.n1607 VDD.n1580 2.25083
R91163 VDD.n1607 VDD.n1579 2.25083
R91164 VDD.n1607 VDD.n1578 2.25083
R91165 VDD.n1607 VDD.n1577 2.25083
R91166 VDD.n1607 VDD.n1576 2.25083
R91167 VDD.n1607 VDD.n1575 2.25083
R91168 VDD.n1607 VDD.n1574 2.25083
R91169 VDD.n1607 VDD.n1573 2.25083
R91170 VDD.n1607 VDD.n1572 2.25083
R91171 VDD.n1607 VDD.n1571 2.25083
R91172 VDD.n1607 VDD.n1570 2.25083
R91173 VDD.n1607 VDD.n1569 2.25083
R91174 VDD.n1607 VDD.n1568 2.25083
R91175 VDD.n1607 VDD.n1567 2.25083
R91176 VDD.n1607 VDD.n1566 2.25083
R91177 VDD.n1607 VDD.n1565 2.25083
R91178 VDD.n1607 VDD.n1564 2.25083
R91179 VDD.n1607 VDD.n1563 2.25083
R91180 VDD.n1607 VDD.n1562 2.25083
R91181 VDD.n1607 VDD.n1561 2.25083
R91182 VDD.n1607 VDD.n1560 2.25083
R91183 VDD.n1607 VDD.n1559 2.25083
R91184 VDD.n1607 VDD.n1558 2.25083
R91185 VDD.n1607 VDD.n1557 2.25083
R91186 VDD.n1607 VDD.n1556 2.25083
R91187 VDD.n1607 VDD.n1555 2.25083
R91188 VDD.n1607 VDD.n1554 2.25083
R91189 VDD.n1607 VDD.n1553 2.25083
R91190 VDD.n1607 VDD.n1552 2.25083
R91191 VDD.n1607 VDD.n1551 2.25083
R91192 VDD.n1607 VDD.n1550 2.25083
R91193 VDD.n1607 VDD.n1549 2.25083
R91194 VDD.n1607 VDD.n1548 2.25083
R91195 VDD.n1607 VDD.n1547 2.25083
R91196 VDD.n1607 VDD.n1546 2.25083
R91197 VDD.n1607 VDD.n1545 2.25083
R91198 VDD.n1416 VDD.n1194 2.25083
R91199 VDD.n1671 VDD.n1670 2.25083
R91200 VDD.n1544 VDD.n1482 2.25083
R91201 VDD.n1671 VDD.n1669 2.25083
R91202 VDD.n1544 VDD.n1483 2.25083
R91203 VDD.n1671 VDD.n1668 2.25083
R91204 VDD.n1544 VDD.n1484 2.25083
R91205 VDD.n1671 VDD.n1667 2.25083
R91206 VDD.n1544 VDD.n1485 2.25083
R91207 VDD.n1671 VDD.n1666 2.25083
R91208 VDD.n1544 VDD.n1486 2.25083
R91209 VDD.n1671 VDD.n1665 2.25083
R91210 VDD.n1544 VDD.n1487 2.25083
R91211 VDD.n1671 VDD.n1664 2.25083
R91212 VDD.n1544 VDD.n1488 2.25083
R91213 VDD.n1671 VDD.n1663 2.25083
R91214 VDD.n1544 VDD.n1489 2.25083
R91215 VDD.n1671 VDD.n1662 2.25083
R91216 VDD.n1544 VDD.n1490 2.25083
R91217 VDD.n1671 VDD.n1661 2.25083
R91218 VDD.n1544 VDD.n1491 2.25083
R91219 VDD.n1671 VDD.n1660 2.25083
R91220 VDD.n1544 VDD.n1492 2.25083
R91221 VDD.n1671 VDD.n1659 2.25083
R91222 VDD.n1544 VDD.n1493 2.25083
R91223 VDD.n1671 VDD.n1658 2.25083
R91224 VDD.n1544 VDD.n1494 2.25083
R91225 VDD.n1671 VDD.n1657 2.25083
R91226 VDD.n1544 VDD.n1495 2.25083
R91227 VDD.n1671 VDD.n1656 2.25083
R91228 VDD.n1544 VDD.n1496 2.25083
R91229 VDD.n1671 VDD.n1655 2.25083
R91230 VDD.n1544 VDD.n1497 2.25083
R91231 VDD.n1671 VDD.n1654 2.25083
R91232 VDD.n1544 VDD.n1498 2.25083
R91233 VDD.n1671 VDD.n1653 2.25083
R91234 VDD.n1544 VDD.n1499 2.25083
R91235 VDD.n1671 VDD.n1652 2.25083
R91236 VDD.n1544 VDD.n1500 2.25083
R91237 VDD.n1671 VDD.n1651 2.25083
R91238 VDD.n1544 VDD.n1501 2.25083
R91239 VDD.n1671 VDD.n1650 2.25083
R91240 VDD.n1544 VDD.n1502 2.25083
R91241 VDD.n1671 VDD.n1649 2.25083
R91242 VDD.n1544 VDD.n1503 2.25083
R91243 VDD.n1671 VDD.n1648 2.25083
R91244 VDD.n1544 VDD.n1504 2.25083
R91245 VDD.n1671 VDD.n1647 2.25083
R91246 VDD.n1544 VDD.n1505 2.25083
R91247 VDD.n1671 VDD.n1646 2.25083
R91248 VDD.n1544 VDD.n1506 2.25083
R91249 VDD.n1671 VDD.n1645 2.25083
R91250 VDD.n1544 VDD.n1507 2.25083
R91251 VDD.n1671 VDD.n1644 2.25083
R91252 VDD.n1544 VDD.n1508 2.25083
R91253 VDD.n1671 VDD.n1643 2.25083
R91254 VDD.n1544 VDD.n1509 2.25083
R91255 VDD.n1671 VDD.n1642 2.25083
R91256 VDD.n1544 VDD.n1510 2.25083
R91257 VDD.n1671 VDD.n1641 2.25083
R91258 VDD.n1544 VDD.n1511 2.25083
R91259 VDD.n1671 VDD.n1640 2.25083
R91260 VDD.n1544 VDD.n1512 2.25083
R91261 VDD.n1671 VDD.n1639 2.25083
R91262 VDD.n1544 VDD.n1513 2.25083
R91263 VDD.n1671 VDD.n1638 2.25083
R91264 VDD.n1544 VDD.n1514 2.25083
R91265 VDD.n1671 VDD.n1637 2.25083
R91266 VDD.n1544 VDD.n1515 2.25083
R91267 VDD.n1671 VDD.n1636 2.25083
R91268 VDD.n1544 VDD.n1516 2.25083
R91269 VDD.n1671 VDD.n1635 2.25083
R91270 VDD.n1544 VDD.n1517 2.25083
R91271 VDD.n1671 VDD.n1634 2.25083
R91272 VDD.n1544 VDD.n1518 2.25083
R91273 VDD.n1671 VDD.n1633 2.25083
R91274 VDD.n1544 VDD.n1519 2.25083
R91275 VDD.n1671 VDD.n1632 2.25083
R91276 VDD.n1544 VDD.n1520 2.25083
R91277 VDD.n1671 VDD.n1631 2.25083
R91278 VDD.n1544 VDD.n1521 2.25083
R91279 VDD.n1671 VDD.n1630 2.25083
R91280 VDD.n1544 VDD.n1522 2.25083
R91281 VDD.n1671 VDD.n1629 2.25083
R91282 VDD.n1544 VDD.n1523 2.25083
R91283 VDD.n1671 VDD.n1628 2.25083
R91284 VDD.n1544 VDD.n1524 2.25083
R91285 VDD.n1671 VDD.n1627 2.25083
R91286 VDD.n1544 VDD.n1525 2.25083
R91287 VDD.n1671 VDD.n1626 2.25083
R91288 VDD.n1544 VDD.n1526 2.25083
R91289 VDD.n1671 VDD.n1625 2.25083
R91290 VDD.n1544 VDD.n1527 2.25083
R91291 VDD.n1671 VDD.n1624 2.25083
R91292 VDD.n1544 VDD.n1528 2.25083
R91293 VDD.n1671 VDD.n1623 2.25083
R91294 VDD.n1544 VDD.n1529 2.25083
R91295 VDD.n1671 VDD.n1622 2.25083
R91296 VDD.n1544 VDD.n1530 2.25083
R91297 VDD.n1671 VDD.n1621 2.25083
R91298 VDD.n1544 VDD.n1531 2.25083
R91299 VDD.n1671 VDD.n1620 2.25083
R91300 VDD.n1544 VDD.n1532 2.25083
R91301 VDD.n1671 VDD.n1619 2.25083
R91302 VDD.n1544 VDD.n1533 2.25083
R91303 VDD.n1671 VDD.n1618 2.25083
R91304 VDD.n1544 VDD.n1534 2.25083
R91305 VDD.n1671 VDD.n1617 2.25083
R91306 VDD.n1544 VDD.n1535 2.25083
R91307 VDD.n1671 VDD.n1616 2.25083
R91308 VDD.n1544 VDD.n1536 2.25083
R91309 VDD.n1671 VDD.n1615 2.25083
R91310 VDD.n1544 VDD.n1537 2.25083
R91311 VDD.n1671 VDD.n1614 2.25083
R91312 VDD.n1544 VDD.n1538 2.25083
R91313 VDD.n1671 VDD.n1613 2.25083
R91314 VDD.n1544 VDD.n1539 2.25083
R91315 VDD.n1671 VDD.n1612 2.25083
R91316 VDD.n1544 VDD.n1540 2.25083
R91317 VDD.n1671 VDD.n1611 2.25083
R91318 VDD.n1544 VDD.n1541 2.25083
R91319 VDD.n1671 VDD.n1610 2.25083
R91320 VDD.n1544 VDD.n1542 2.25083
R91321 VDD.n1671 VDD.n1609 2.25083
R91322 VDD.n1544 VDD.n1543 2.25083
R91323 VDD.n1671 VDD.n1608 2.25083
R91324 VDD.n1544 VDD.n1258 2.25083
R91325 VDD.n1671 VDD.n1259 2.25083
R91326 VDD.n487 VDD.n486 1.51655
R91327 VDD.n481 VDD.n480 1.51655
R91328 VDD.n477 VDD.n476 1.51655
R91329 VDD.n471 VDD.n470 1.51655
R91330 VDD.n465 VDD.n464 1.51655
R91331 VDD.n459 VDD.n458 1.51655
R91332 VDD.n453 VDD.n452 1.51655
R91333 VDD.n449 VDD.n448 1.51655
R91334 VDD.n443 VDD.n442 1.51655
R91335 VDD.n439 VDD.n438 1.51655
R91336 VDD.n691 VDD.n690 1.51655
R91337 VDD.n949 VDD.n406 1.51655
R91338 VDD.n428 VDD.n427 1.51655
R91339 VDD.n425 VDD.n424 1.50629
R91340 VDD.n767 VDD.n766 0.9005
R91341 VDD.n694 VDD.n693 0.9005
R91342 VDD.n719 VDD.n694 0.9005
R91343 VDD.n718 VDD.n717 0.9005
R91344 VDD.n953 VDD.n952 0.9005
R91345 VDD.n952 VDD.n951 0.9005
R91346 VDD.n708 VDD.n403 0.9005
R91347 VDD.n950 VDD.n949 0.9005
R91348 VDD.n951 VDD.n950 0.9005
R91349 VDD.n692 VDD.n691 0.9005
R91350 VDD.n719 VDD.n692 0.9005
R91351 VDD.n721 VDD.n720 0.9005
R91352 VDD.n731 VDD.n730 0.9005
R91353 VDD.n734 VDD.n733 0.9005
R91354 VDD.n764 VDD.n763 0.9005
R91355 VDD.n405 VDD.n404 0.9005
R91356 VDD.n734 VDD.n383 0.684974
R91357 VDD.n486 VDD.t43 0.6505
R91358 VDD.n486 VDD.t27 0.6505
R91359 VDD.n480 VDD.t11 0.6505
R91360 VDD.n480 VDD.t1 0.6505
R91361 VDD.n476 VDD.t41 0.6505
R91362 VDD.n476 VDD.t5 0.6505
R91363 VDD.n470 VDD.t51 0.6505
R91364 VDD.n470 VDD.t33 0.6505
R91365 VDD.n464 VDD.t23 0.6505
R91366 VDD.n464 VDD.t7 0.6505
R91367 VDD.n458 VDD.t25 0.6505
R91368 VDD.n458 VDD.t9 0.6505
R91369 VDD.n452 VDD.t13 0.6505
R91370 VDD.n452 VDD.t37 0.6505
R91371 VDD.n448 VDD.t19 0.6505
R91372 VDD.n448 VDD.t49 0.6505
R91373 VDD.n442 VDD.t21 0.6505
R91374 VDD.n442 VDD.t35 0.6505
R91375 VDD.n438 VDD.t55 0.6505
R91376 VDD.n438 VDD.t47 0.6505
R91377 VDD.n424 VDD.t39 0.6505
R91378 VDD.n424 VDD.t15 0.6505
R91379 VDD.n690 VDD.t31 0.6505
R91380 VDD.n690 VDD.t17 0.6505
R91381 VDD.n406 VDD.t29 0.6505
R91382 VDD.n406 VDD.t53 0.6505
R91383 VDD.n427 VDD.t3 0.6505
R91384 VDD.n427 VDD.t45 0.6505
R91385 VDD.n763 VDD.n762 0.611553
R91386 VDD.n674 VDD.n385 0.573227
R91387 VDD.n732 VDD.n674 0.573227
R91388 VDD.n673 VDD.n426 0.573227
R91389 VDD.n732 VDD.n673 0.573227
R91390 VDD.n699 VDD.n696 0.3965
R91391 VDD.n716 VDD.n715 0.3965
R91392 VDD.n698 VDD.n697 0.3965
R91393 VDD.n695 VDD.n412 0.3965
R91394 VDD.n770 VDD.n663 0.365
R91395 VDD.n769 VDD.n768 0.365
R91396 VDD.n667 VDD.n665 0.365
R91397 VDD.n666 VDD.n493 0.365
R91398 VDD.n1069 VDD.n277 0.355706
R91399 VDD.n1073 VDD.n277 0.355706
R91400 VDD.n980 VDD.n979 0.345348
R91401 VDD.n798 VDD.n639 0.345348
R91402 VDD.n672 VDD.n431 0.34025
R91403 VDD.n761 VDD.n640 0.32225
R91404 VDD.n760 VDD.n641 0.32225
R91405 VDD.n759 VDD.n642 0.32225
R91406 VDD.n758 VDD.n643 0.32225
R91407 VDD.n757 VDD.n644 0.32225
R91408 VDD.n756 VDD.n645 0.32225
R91409 VDD.n755 VDD.n646 0.32225
R91410 VDD.n754 VDD.n647 0.32225
R91411 VDD.n753 VDD.n648 0.32225
R91412 VDD.n751 VDD.n649 0.32225
R91413 VDD.n750 VDD.n650 0.32225
R91414 VDD.n749 VDD.n651 0.32225
R91415 VDD.n748 VDD.n652 0.32225
R91416 VDD.n747 VDD.n653 0.32225
R91417 VDD.n746 VDD.n654 0.32225
R91418 VDD.n745 VDD.n655 0.32225
R91419 VDD.n744 VDD.n656 0.32225
R91420 VDD.n743 VDD.n657 0.32225
R91421 VDD.n742 VDD.n658 0.32225
R91422 VDD.n964 VDD.n396 0.32225
R91423 VDD.n965 VDD.n395 0.32225
R91424 VDD.n978 VDD.n383 0.32225
R91425 VDD.n977 VDD.n384 0.32225
R91426 VDD.n976 VDD.n385 0.32225
R91427 VDD.n975 VDD.n386 0.32225
R91428 VDD.n974 VDD.n387 0.32225
R91429 VDD.n966 VDD.n394 0.32225
R91430 VDD.n957 VDD.n402 0.32225
R91431 VDD.n956 VDD.n953 0.32225
R91432 VDD.n955 VDD.n954 0.32225
R91433 VDD.n736 VDD.n735 0.31775
R91434 VDD.n679 VDD.n677 0.31775
R91435 VDD.n675 VDD.n421 0.31775
R91436 VDD.n678 VDD.n676 0.31775
R91437 VDD.n729 VDD.n728 0.31775
R91438 VDD.n874 VDD.n565 0.292176
R91439 VDD.n707 VDD.n704 0.2885
R91440 VDD.n712 VDD.n711 0.2885
R91441 VDD.n710 VDD.n705 0.2885
R91442 VDD.n706 VDD.n409 0.2885
R91443 VDD.n878 VDD.n565 0.282618
R91444 VDD.n954 VDD.n266 0.279974
R91445 VDD.n967 VDD.n393 0.2795
R91446 VDD.n762 VDD.n639 0.2795
R91447 VDD.n677 VDD.n387 0.277605
R91448 VDD.n566 VDD.n563 0.2705
R91449 VDD.n772 VDD.n555 0.2705
R91450 VDD.n772 VDD.n661 0.2705
R91451 VDD.n771 VDD.n554 0.2705
R91452 VDD.n771 VDD.n770 0.2705
R91453 VDD.n662 VDD.n553 0.2705
R91454 VDD.n769 VDD.n662 0.2705
R91455 VDD.n664 VDD.n552 0.2705
R91456 VDD.n665 VDD.n664 0.2705
R91457 VDD.n497 VDD.n495 0.2705
R91458 VDD.n495 VDD.n493 0.2705
R91459 VDD.n389 VDD.n388 0.2705
R91460 VDD.n390 VDD.n389 0.2705
R91461 VDD.n391 VDD.n390 0.2705
R91462 VDD.n392 VDD.n391 0.2705
R91463 VDD.n681 VDD.n679 0.2705
R91464 VDD.n683 VDD.n681 0.2705
R91465 VDD.n685 VDD.n683 0.2705
R91466 VDD.n686 VDD.n685 0.2705
R91467 VDD.n701 VDD.n699 0.2705
R91468 VDD.n703 VDD.n701 0.2705
R91469 VDD.n704 VDD.n703 0.2705
R91470 VDD.n715 VDD.n714 0.2705
R91471 VDD.n714 VDD.n713 0.2705
R91472 VDD.n713 VDD.n712 0.2705
R91473 VDD.n700 VDD.n698 0.2705
R91474 VDD.n702 VDD.n700 0.2705
R91475 VDD.n705 VDD.n702 0.2705
R91476 VDD.n398 VDD.n397 0.2705
R91477 VDD.n399 VDD.n398 0.2705
R91478 VDD.n400 VDD.n399 0.2705
R91479 VDD.n401 VDD.n400 0.2705
R91480 VDD.n412 VDD.n411 0.2705
R91481 VDD.n411 VDD.n410 0.2705
R91482 VDD.n410 VDD.n409 0.2705
R91483 VDD.n421 VDD.n420 0.2705
R91484 VDD.n420 VDD.n419 0.2705
R91485 VDD.n419 VDD.n418 0.2705
R91486 VDD.n418 VDD.n417 0.2705
R91487 VDD.n680 VDD.n678 0.2705
R91488 VDD.n682 VDD.n680 0.2705
R91489 VDD.n684 VDD.n682 0.2705
R91490 VDD.n687 VDD.n684 0.2705
R91491 VDD.n728 VDD.n727 0.2705
R91492 VDD.n727 VDD.n726 0.2705
R91493 VDD.n726 VDD.n725 0.2705
R91494 VDD.n725 VDD.n724 0.2705
R91495 VDD.n435 VDD.n434 0.2705
R91496 VDD.n434 VDD.n433 0.2705
R91497 VDD.n433 VDD.n432 0.2705
R91498 VDD.n432 VDD.n431 0.2705
R91499 VDD.n773 VDD.n556 0.2705
R91500 VDD.n773 VDD.n660 0.2705
R91501 VDD.n660 VDD.n659 0.2705
R91502 VDD.n659 VDD.n658 0.2705
R91503 VDD.n658 VDD.n657 0.2705
R91504 VDD.n657 VDD.n656 0.2705
R91505 VDD.n656 VDD.n655 0.2705
R91506 VDD.n655 VDD.n654 0.2705
R91507 VDD.n654 VDD.n653 0.2705
R91508 VDD.n653 VDD.n652 0.2705
R91509 VDD.n652 VDD.n651 0.2705
R91510 VDD.n651 VDD.n650 0.2705
R91511 VDD.n650 VDD.n649 0.2705
R91512 VDD.n649 VDD.n648 0.2705
R91513 VDD.n648 VDD.n647 0.2705
R91514 VDD.n647 VDD.n646 0.2705
R91515 VDD.n646 VDD.n645 0.2705
R91516 VDD.n645 VDD.n644 0.2705
R91517 VDD.n644 VDD.n643 0.2705
R91518 VDD.n643 VDD.n642 0.2705
R91519 VDD.n642 VDD.n641 0.2705
R91520 VDD.n641 VDD.n640 0.2705
R91521 VDD.n640 VDD.n639 0.2705
R91522 VDD.n774 VDD.n557 0.2705
R91523 VDD.n775 VDD.n774 0.2705
R91524 VDD.n776 VDD.n775 0.2705
R91525 VDD.n777 VDD.n776 0.2705
R91526 VDD.n778 VDD.n777 0.2705
R91527 VDD.n779 VDD.n778 0.2705
R91528 VDD.n780 VDD.n779 0.2705
R91529 VDD.n781 VDD.n780 0.2705
R91530 VDD.n782 VDD.n781 0.2705
R91531 VDD.n783 VDD.n782 0.2705
R91532 VDD.n784 VDD.n783 0.2705
R91533 VDD.n785 VDD.n784 0.2705
R91534 VDD.n786 VDD.n785 0.2705
R91535 VDD.n787 VDD.n786 0.2705
R91536 VDD.n788 VDD.n787 0.2705
R91537 VDD.n789 VDD.n788 0.2705
R91538 VDD.n790 VDD.n789 0.2705
R91539 VDD.n791 VDD.n790 0.2705
R91540 VDD.n792 VDD.n791 0.2705
R91541 VDD.n793 VDD.n792 0.2705
R91542 VDD.n794 VDD.n793 0.2705
R91543 VDD.n795 VDD.n794 0.2705
R91544 VDD.n796 VDD.n795 0.2705
R91545 VDD.n797 VDD.n796 0.2705
R91546 VDD.n615 VDD.n558 0.2705
R91547 VDD.n616 VDD.n615 0.2705
R91548 VDD.n617 VDD.n616 0.2705
R91549 VDD.n618 VDD.n617 0.2705
R91550 VDD.n619 VDD.n618 0.2705
R91551 VDD.n620 VDD.n619 0.2705
R91552 VDD.n621 VDD.n620 0.2705
R91553 VDD.n622 VDD.n621 0.2705
R91554 VDD.n623 VDD.n622 0.2705
R91555 VDD.n624 VDD.n623 0.2705
R91556 VDD.n625 VDD.n624 0.2705
R91557 VDD.n626 VDD.n625 0.2705
R91558 VDD.n627 VDD.n626 0.2705
R91559 VDD.n628 VDD.n627 0.2705
R91560 VDD.n629 VDD.n628 0.2705
R91561 VDD.n630 VDD.n629 0.2705
R91562 VDD.n631 VDD.n630 0.2705
R91563 VDD.n632 VDD.n631 0.2705
R91564 VDD.n633 VDD.n632 0.2705
R91565 VDD.n634 VDD.n633 0.2705
R91566 VDD.n635 VDD.n634 0.2705
R91567 VDD.n636 VDD.n635 0.2705
R91568 VDD.n637 VDD.n636 0.2705
R91569 VDD.n638 VDD.n637 0.2705
R91570 VDD.n824 VDD.n559 0.2705
R91571 VDD.n824 VDD.n823 0.2705
R91572 VDD.n823 VDD.n822 0.2705
R91573 VDD.n822 VDD.n821 0.2705
R91574 VDD.n821 VDD.n820 0.2705
R91575 VDD.n820 VDD.n819 0.2705
R91576 VDD.n819 VDD.n818 0.2705
R91577 VDD.n818 VDD.n817 0.2705
R91578 VDD.n817 VDD.n816 0.2705
R91579 VDD.n816 VDD.n815 0.2705
R91580 VDD.n815 VDD.n814 0.2705
R91581 VDD.n814 VDD.n813 0.2705
R91582 VDD.n813 VDD.n812 0.2705
R91583 VDD.n812 VDD.n811 0.2705
R91584 VDD.n811 VDD.n810 0.2705
R91585 VDD.n810 VDD.n809 0.2705
R91586 VDD.n809 VDD.n808 0.2705
R91587 VDD.n808 VDD.n807 0.2705
R91588 VDD.n807 VDD.n806 0.2705
R91589 VDD.n806 VDD.n805 0.2705
R91590 VDD.n805 VDD.n804 0.2705
R91591 VDD.n804 VDD.n803 0.2705
R91592 VDD.n803 VDD.n802 0.2705
R91593 VDD.n802 VDD.n801 0.2705
R91594 VDD.n825 VDD.n560 0.2705
R91595 VDD.n825 VDD.n613 0.2705
R91596 VDD.n613 VDD.n612 0.2705
R91597 VDD.n612 VDD.n611 0.2705
R91598 VDD.n611 VDD.n610 0.2705
R91599 VDD.n610 VDD.n609 0.2705
R91600 VDD.n609 VDD.n608 0.2705
R91601 VDD.n608 VDD.n607 0.2705
R91602 VDD.n607 VDD.n606 0.2705
R91603 VDD.n606 VDD.n605 0.2705
R91604 VDD.n605 VDD.n604 0.2705
R91605 VDD.n604 VDD.n603 0.2705
R91606 VDD.n603 VDD.n602 0.2705
R91607 VDD.n602 VDD.n601 0.2705
R91608 VDD.n601 VDD.n600 0.2705
R91609 VDD.n600 VDD.n599 0.2705
R91610 VDD.n599 VDD.n598 0.2705
R91611 VDD.n598 VDD.n597 0.2705
R91612 VDD.n597 VDD.n596 0.2705
R91613 VDD.n596 VDD.n595 0.2705
R91614 VDD.n595 VDD.n594 0.2705
R91615 VDD.n594 VDD.n593 0.2705
R91616 VDD.n593 VDD.n592 0.2705
R91617 VDD.n592 VDD.n591 0.2705
R91618 VDD.n826 VDD.n561 0.2705
R91619 VDD.n827 VDD.n826 0.2705
R91620 VDD.n828 VDD.n827 0.2705
R91621 VDD.n829 VDD.n828 0.2705
R91622 VDD.n830 VDD.n829 0.2705
R91623 VDD.n831 VDD.n830 0.2705
R91624 VDD.n832 VDD.n831 0.2705
R91625 VDD.n833 VDD.n832 0.2705
R91626 VDD.n834 VDD.n833 0.2705
R91627 VDD.n835 VDD.n834 0.2705
R91628 VDD.n836 VDD.n835 0.2705
R91629 VDD.n837 VDD.n836 0.2705
R91630 VDD.n838 VDD.n837 0.2705
R91631 VDD.n839 VDD.n838 0.2705
R91632 VDD.n840 VDD.n839 0.2705
R91633 VDD.n841 VDD.n840 0.2705
R91634 VDD.n842 VDD.n841 0.2705
R91635 VDD.n843 VDD.n842 0.2705
R91636 VDD.n844 VDD.n843 0.2705
R91637 VDD.n845 VDD.n844 0.2705
R91638 VDD.n846 VDD.n845 0.2705
R91639 VDD.n847 VDD.n846 0.2705
R91640 VDD.n848 VDD.n847 0.2705
R91641 VDD.n849 VDD.n848 0.2705
R91642 VDD.n614 VDD.n562 0.2705
R91643 VDD.n614 VDD.n567 0.2705
R91644 VDD.n568 VDD.n567 0.2705
R91645 VDD.n569 VDD.n568 0.2705
R91646 VDD.n570 VDD.n569 0.2705
R91647 VDD.n571 VDD.n570 0.2705
R91648 VDD.n572 VDD.n571 0.2705
R91649 VDD.n573 VDD.n572 0.2705
R91650 VDD.n574 VDD.n573 0.2705
R91651 VDD.n575 VDD.n574 0.2705
R91652 VDD.n576 VDD.n575 0.2705
R91653 VDD.n577 VDD.n576 0.2705
R91654 VDD.n578 VDD.n577 0.2705
R91655 VDD.n579 VDD.n578 0.2705
R91656 VDD.n580 VDD.n579 0.2705
R91657 VDD.n581 VDD.n580 0.2705
R91658 VDD.n582 VDD.n581 0.2705
R91659 VDD.n583 VDD.n582 0.2705
R91660 VDD.n584 VDD.n583 0.2705
R91661 VDD.n585 VDD.n584 0.2705
R91662 VDD.n586 VDD.n585 0.2705
R91663 VDD.n587 VDD.n586 0.2705
R91664 VDD.n588 VDD.n587 0.2705
R91665 VDD.n589 VDD.n588 0.2705
R91666 VDD.n875 VDD.n564 0.2705
R91667 VDD.n875 VDD.n874 0.2705
R91668 VDD.n877 VDD.n876 0.2705
R91669 VDD.n549 VDD.n548 0.2705
R91670 VDD.n548 VDD.n547 0.2705
R91671 VDD.n547 VDD.n546 0.2705
R91672 VDD.n546 VDD.n545 0.2705
R91673 VDD.n545 VDD.n544 0.2705
R91674 VDD.n544 VDD.n543 0.2705
R91675 VDD.n543 VDD.n542 0.2705
R91676 VDD.n542 VDD.n541 0.2705
R91677 VDD.n541 VDD.n540 0.2705
R91678 VDD.n540 VDD.n539 0.2705
R91679 VDD.n539 VDD.n538 0.2705
R91680 VDD.n538 VDD.n537 0.2705
R91681 VDD.n537 VDD.n536 0.2705
R91682 VDD.n536 VDD.n535 0.2705
R91683 VDD.n535 VDD.n534 0.2705
R91684 VDD.n534 VDD.n533 0.2705
R91685 VDD.n533 VDD.n532 0.2705
R91686 VDD.n532 VDD.n169 0.2705
R91687 VDD.n1126 VDD.n169 0.2705
R91688 VDD.n1126 VDD.n1125 0.2705
R91689 VDD.n1125 VDD.n1124 0.2705
R91690 VDD.n1124 VDD.n1123 0.2705
R91691 VDD.n1123 VDD.n1122 0.2705
R91692 VDD.n1122 VDD.n1121 0.2705
R91693 VDD.n1121 VDD.n1120 0.2705
R91694 VDD.n1120 VDD.n1119 0.2705
R91695 VDD.n1119 VDD.n1118 0.2705
R91696 VDD.n1118 VDD.n1117 0.2705
R91697 VDD.n1117 VDD.n1116 0.2705
R91698 VDD.n1116 VDD.n1115 0.2705
R91699 VDD.n1115 VDD.n1114 0.2705
R91700 VDD.n1114 VDD.n1113 0.2705
R91701 VDD.n1113 VDD.n1112 0.2705
R91702 VDD.n1112 VDD.n1111 0.2705
R91703 VDD.n1111 VDD.n1110 0.2705
R91704 VDD.n1110 VDD.n1109 0.2705
R91705 VDD.n1109 VDD.n1108 0.2705
R91706 VDD.n1108 VDD.n1107 0.2705
R91707 VDD.n1107 VDD.n1106 0.2705
R91708 VDD.n1106 VDD.n1105 0.2705
R91709 VDD.n1105 VDD.n1104 0.2705
R91710 VDD.n1104 VDD.n1103 0.2705
R91711 VDD.n1103 VDD.n1102 0.2705
R91712 VDD.n1102 VDD.n1101 0.2705
R91713 VDD.n1101 VDD.n1100 0.2705
R91714 VDD.n1100 VDD.n1099 0.2705
R91715 VDD.n1099 VDD.n1098 0.2705
R91716 VDD.n1098 VDD.n1097 0.2705
R91717 VDD.n1097 VDD.n1096 0.2705
R91718 VDD.n1096 VDD.n1095 0.2705
R91719 VDD.n1095 VDD.n1094 0.2705
R91720 VDD.n1094 VDD.n1093 0.2705
R91721 VDD.n1093 VDD.n1092 0.2705
R91722 VDD.n1092 VDD.n239 0.2705
R91723 VDD.n496 VDD.n494 0.2705
R91724 VDD.n494 VDD.n492 0.2705
R91725 VDD.n492 VDD.n491 0.2705
R91726 VDD.n491 VDD.n489 0.2705
R91727 VDD.n489 VDD.n485 0.2705
R91728 VDD.n485 VDD.n483 0.2705
R91729 VDD.n483 VDD.n479 0.2705
R91730 VDD.n479 VDD.n475 0.2705
R91731 VDD.n475 VDD.n473 0.2705
R91732 VDD.n473 VDD.n469 0.2705
R91733 VDD.n469 VDD.n467 0.2705
R91734 VDD.n467 VDD.n463 0.2705
R91735 VDD.n463 VDD.n461 0.2705
R91736 VDD.n461 VDD.n457 0.2705
R91737 VDD.n457 VDD.n455 0.2705
R91738 VDD.n455 VDD.n451 0.2705
R91739 VDD.n451 VDD.n447 0.2705
R91740 VDD.n447 VDD.n445 0.2705
R91741 VDD.n445 VDD.n171 0.2705
R91742 VDD.n173 VDD.n171 0.2705
R91743 VDD.n175 VDD.n173 0.2705
R91744 VDD.n177 VDD.n175 0.2705
R91745 VDD.n179 VDD.n177 0.2705
R91746 VDD.n181 VDD.n179 0.2705
R91747 VDD.n183 VDD.n181 0.2705
R91748 VDD.n185 VDD.n183 0.2705
R91749 VDD.n187 VDD.n185 0.2705
R91750 VDD.n189 VDD.n187 0.2705
R91751 VDD.n191 VDD.n189 0.2705
R91752 VDD.n193 VDD.n191 0.2705
R91753 VDD.n195 VDD.n193 0.2705
R91754 VDD.n197 VDD.n195 0.2705
R91755 VDD.n199 VDD.n197 0.2705
R91756 VDD.n201 VDD.n199 0.2705
R91757 VDD.n203 VDD.n201 0.2705
R91758 VDD.n205 VDD.n203 0.2705
R91759 VDD.n207 VDD.n205 0.2705
R91760 VDD.n209 VDD.n207 0.2705
R91761 VDD.n211 VDD.n209 0.2705
R91762 VDD.n213 VDD.n211 0.2705
R91763 VDD.n215 VDD.n213 0.2705
R91764 VDD.n217 VDD.n215 0.2705
R91765 VDD.n219 VDD.n217 0.2705
R91766 VDD.n221 VDD.n219 0.2705
R91767 VDD.n223 VDD.n221 0.2705
R91768 VDD.n225 VDD.n223 0.2705
R91769 VDD.n227 VDD.n225 0.2705
R91770 VDD.n229 VDD.n227 0.2705
R91771 VDD.n231 VDD.n229 0.2705
R91772 VDD.n233 VDD.n231 0.2705
R91773 VDD.n235 VDD.n233 0.2705
R91774 VDD.n237 VDD.n235 0.2705
R91775 VDD.n1091 VDD.n237 0.2705
R91776 VDD.n1091 VDD.n1090 0.2705
R91777 VDD.n895 VDD.n894 0.2705
R91778 VDD.n896 VDD.n895 0.2705
R91779 VDD.n897 VDD.n896 0.2705
R91780 VDD.n898 VDD.n897 0.2705
R91781 VDD.n899 VDD.n898 0.2705
R91782 VDD.n900 VDD.n899 0.2705
R91783 VDD.n901 VDD.n900 0.2705
R91784 VDD.n902 VDD.n901 0.2705
R91785 VDD.n903 VDD.n902 0.2705
R91786 VDD.n904 VDD.n903 0.2705
R91787 VDD.n905 VDD.n904 0.2705
R91788 VDD.n906 VDD.n905 0.2705
R91789 VDD.n907 VDD.n906 0.2705
R91790 VDD.n908 VDD.n907 0.2705
R91791 VDD.n909 VDD.n908 0.2705
R91792 VDD.n910 VDD.n909 0.2705
R91793 VDD.n911 VDD.n910 0.2705
R91794 VDD.n912 VDD.n911 0.2705
R91795 VDD.n913 VDD.n912 0.2705
R91796 VDD.n914 VDD.n913 0.2705
R91797 VDD.n915 VDD.n914 0.2705
R91798 VDD.n916 VDD.n915 0.2705
R91799 VDD.n917 VDD.n916 0.2705
R91800 VDD.n918 VDD.n917 0.2705
R91801 VDD.n919 VDD.n918 0.2705
R91802 VDD.n920 VDD.n919 0.2705
R91803 VDD.n921 VDD.n920 0.2705
R91804 VDD.n922 VDD.n921 0.2705
R91805 VDD.n923 VDD.n922 0.2705
R91806 VDD.n924 VDD.n923 0.2705
R91807 VDD.n925 VDD.n924 0.2705
R91808 VDD.n926 VDD.n925 0.2705
R91809 VDD.n927 VDD.n926 0.2705
R91810 VDD.n928 VDD.n927 0.2705
R91811 VDD.n929 VDD.n928 0.2705
R91812 VDD.n930 VDD.n929 0.2705
R91813 VDD.n931 VDD.n930 0.2705
R91814 VDD.n932 VDD.n931 0.2705
R91815 VDD.n933 VDD.n932 0.2705
R91816 VDD.n934 VDD.n933 0.2705
R91817 VDD.n935 VDD.n934 0.2705
R91818 VDD.n936 VDD.n935 0.2705
R91819 VDD.n937 VDD.n936 0.2705
R91820 VDD.n938 VDD.n937 0.2705
R91821 VDD.n939 VDD.n938 0.2705
R91822 VDD.n940 VDD.n939 0.2705
R91823 VDD.n941 VDD.n940 0.2705
R91824 VDD.n942 VDD.n941 0.2705
R91825 VDD.n943 VDD.n942 0.2705
R91826 VDD.n944 VDD.n943 0.2705
R91827 VDD.n945 VDD.n944 0.2705
R91828 VDD.n946 VDD.n945 0.2705
R91829 VDD.n946 VDD.n240 0.2705
R91830 VDD.n1089 VDD.n240 0.2705
R91831 VDD.n1087 VDD.n263 0.2705
R91832 VDD.n1086 VDD.n264 0.2705
R91833 VDD.n1085 VDD.n265 0.2705
R91834 VDD.n1084 VDD.n266 0.2705
R91835 VDD.n979 VDD.n978 0.2705
R91836 VDD.n978 VDD.n977 0.2705
R91837 VDD.n977 VDD.n976 0.2705
R91838 VDD.n976 VDD.n975 0.2705
R91839 VDD.n975 VDD.n974 0.2705
R91840 VDD.n974 VDD.n973 0.2705
R91841 VDD.n973 VDD.n972 0.2705
R91842 VDD.n972 VDD.n971 0.2705
R91843 VDD.n971 VDD.n970 0.2705
R91844 VDD.n970 VDD.n969 0.2705
R91845 VDD.n969 VDD.n968 0.2705
R91846 VDD.n968 VDD.n967 0.2705
R91847 VDD.n967 VDD.n966 0.2705
R91848 VDD.n966 VDD.n965 0.2705
R91849 VDD.n965 VDD.n964 0.2705
R91850 VDD.n964 VDD.n963 0.2705
R91851 VDD.n963 VDD.n962 0.2705
R91852 VDD.n962 VDD.n961 0.2705
R91853 VDD.n961 VDD.n960 0.2705
R91854 VDD.n960 VDD.n959 0.2705
R91855 VDD.n959 VDD.n958 0.2705
R91856 VDD.n958 VDD.n957 0.2705
R91857 VDD.n957 VDD.n956 0.2705
R91858 VDD.n956 VDD.n955 0.2705
R91859 VDD.n955 VDD.n267 0.2705
R91860 VDD.n382 VDD.n381 0.2705
R91861 VDD.n381 VDD.n380 0.2705
R91862 VDD.n380 VDD.n379 0.2705
R91863 VDD.n379 VDD.n378 0.2705
R91864 VDD.n378 VDD.n377 0.2705
R91865 VDD.n377 VDD.n376 0.2705
R91866 VDD.n376 VDD.n375 0.2705
R91867 VDD.n375 VDD.n374 0.2705
R91868 VDD.n374 VDD.n373 0.2705
R91869 VDD.n373 VDD.n372 0.2705
R91870 VDD.n372 VDD.n371 0.2705
R91871 VDD.n371 VDD.n370 0.2705
R91872 VDD.n370 VDD.n369 0.2705
R91873 VDD.n369 VDD.n368 0.2705
R91874 VDD.n368 VDD.n367 0.2705
R91875 VDD.n367 VDD.n366 0.2705
R91876 VDD.n366 VDD.n365 0.2705
R91877 VDD.n365 VDD.n364 0.2705
R91878 VDD.n364 VDD.n363 0.2705
R91879 VDD.n363 VDD.n362 0.2705
R91880 VDD.n362 VDD.n361 0.2705
R91881 VDD.n361 VDD.n360 0.2705
R91882 VDD.n360 VDD.n359 0.2705
R91883 VDD.n359 VDD.n358 0.2705
R91884 VDD.n358 VDD.n357 0.2705
R91885 VDD.n357 VDD.n268 0.2705
R91886 VDD.n983 VDD.n982 0.2705
R91887 VDD.n984 VDD.n983 0.2705
R91888 VDD.n985 VDD.n984 0.2705
R91889 VDD.n986 VDD.n985 0.2705
R91890 VDD.n987 VDD.n986 0.2705
R91891 VDD.n988 VDD.n987 0.2705
R91892 VDD.n989 VDD.n988 0.2705
R91893 VDD.n990 VDD.n989 0.2705
R91894 VDD.n991 VDD.n990 0.2705
R91895 VDD.n992 VDD.n991 0.2705
R91896 VDD.n993 VDD.n992 0.2705
R91897 VDD.n994 VDD.n993 0.2705
R91898 VDD.n995 VDD.n994 0.2705
R91899 VDD.n996 VDD.n995 0.2705
R91900 VDD.n997 VDD.n996 0.2705
R91901 VDD.n998 VDD.n997 0.2705
R91902 VDD.n999 VDD.n998 0.2705
R91903 VDD.n1000 VDD.n999 0.2705
R91904 VDD.n1001 VDD.n1000 0.2705
R91905 VDD.n1002 VDD.n1001 0.2705
R91906 VDD.n1003 VDD.n1002 0.2705
R91907 VDD.n1004 VDD.n1003 0.2705
R91908 VDD.n1005 VDD.n1004 0.2705
R91909 VDD.n1006 VDD.n1005 0.2705
R91910 VDD.n1007 VDD.n1006 0.2705
R91911 VDD.n1007 VDD.n269 0.2705
R91912 VDD.n333 VDD.n332 0.2705
R91913 VDD.n334 VDD.n333 0.2705
R91914 VDD.n335 VDD.n334 0.2705
R91915 VDD.n336 VDD.n335 0.2705
R91916 VDD.n337 VDD.n336 0.2705
R91917 VDD.n338 VDD.n337 0.2705
R91918 VDD.n339 VDD.n338 0.2705
R91919 VDD.n340 VDD.n339 0.2705
R91920 VDD.n341 VDD.n340 0.2705
R91921 VDD.n342 VDD.n341 0.2705
R91922 VDD.n343 VDD.n342 0.2705
R91923 VDD.n344 VDD.n343 0.2705
R91924 VDD.n345 VDD.n344 0.2705
R91925 VDD.n346 VDD.n345 0.2705
R91926 VDD.n347 VDD.n346 0.2705
R91927 VDD.n348 VDD.n347 0.2705
R91928 VDD.n349 VDD.n348 0.2705
R91929 VDD.n350 VDD.n349 0.2705
R91930 VDD.n351 VDD.n350 0.2705
R91931 VDD.n352 VDD.n351 0.2705
R91932 VDD.n353 VDD.n352 0.2705
R91933 VDD.n354 VDD.n353 0.2705
R91934 VDD.n355 VDD.n354 0.2705
R91935 VDD.n356 VDD.n355 0.2705
R91936 VDD.n1008 VDD.n356 0.2705
R91937 VDD.n1008 VDD.n270 0.2705
R91938 VDD.n1034 VDD.n1033 0.2705
R91939 VDD.n1033 VDD.n1032 0.2705
R91940 VDD.n1032 VDD.n1031 0.2705
R91941 VDD.n1031 VDD.n1030 0.2705
R91942 VDD.n1030 VDD.n1029 0.2705
R91943 VDD.n1029 VDD.n1028 0.2705
R91944 VDD.n1028 VDD.n1027 0.2705
R91945 VDD.n1027 VDD.n1026 0.2705
R91946 VDD.n1026 VDD.n1025 0.2705
R91947 VDD.n1025 VDD.n1024 0.2705
R91948 VDD.n1024 VDD.n1023 0.2705
R91949 VDD.n1023 VDD.n1022 0.2705
R91950 VDD.n1022 VDD.n1021 0.2705
R91951 VDD.n1021 VDD.n1020 0.2705
R91952 VDD.n1020 VDD.n1019 0.2705
R91953 VDD.n1019 VDD.n1018 0.2705
R91954 VDD.n1018 VDD.n1017 0.2705
R91955 VDD.n1017 VDD.n1016 0.2705
R91956 VDD.n1016 VDD.n1015 0.2705
R91957 VDD.n1015 VDD.n1014 0.2705
R91958 VDD.n1014 VDD.n1013 0.2705
R91959 VDD.n1013 VDD.n1012 0.2705
R91960 VDD.n1012 VDD.n1011 0.2705
R91961 VDD.n1011 VDD.n1010 0.2705
R91962 VDD.n1010 VDD.n1009 0.2705
R91963 VDD.n1009 VDD.n271 0.2705
R91964 VDD.n330 VDD.n328 0.2705
R91965 VDD.n328 VDD.n326 0.2705
R91966 VDD.n326 VDD.n324 0.2705
R91967 VDD.n324 VDD.n322 0.2705
R91968 VDD.n322 VDD.n320 0.2705
R91969 VDD.n320 VDD.n318 0.2705
R91970 VDD.n318 VDD.n316 0.2705
R91971 VDD.n316 VDD.n314 0.2705
R91972 VDD.n314 VDD.n312 0.2705
R91973 VDD.n312 VDD.n310 0.2705
R91974 VDD.n310 VDD.n308 0.2705
R91975 VDD.n308 VDD.n306 0.2705
R91976 VDD.n306 VDD.n304 0.2705
R91977 VDD.n304 VDD.n302 0.2705
R91978 VDD.n302 VDD.n300 0.2705
R91979 VDD.n300 VDD.n298 0.2705
R91980 VDD.n298 VDD.n296 0.2705
R91981 VDD.n296 VDD.n294 0.2705
R91982 VDD.n294 VDD.n292 0.2705
R91983 VDD.n292 VDD.n290 0.2705
R91984 VDD.n290 VDD.n288 0.2705
R91985 VDD.n288 VDD.n286 0.2705
R91986 VDD.n286 VDD.n284 0.2705
R91987 VDD.n284 VDD.n283 0.2705
R91988 VDD.n283 VDD.n282 0.2705
R91989 VDD.n282 VDD.n272 0.2705
R91990 VDD.n1039 VDD.n1038 0.2705
R91991 VDD.n1040 VDD.n1039 0.2705
R91992 VDD.n1041 VDD.n1040 0.2705
R91993 VDD.n1042 VDD.n1041 0.2705
R91994 VDD.n1043 VDD.n1042 0.2705
R91995 VDD.n1044 VDD.n1043 0.2705
R91996 VDD.n1045 VDD.n1044 0.2705
R91997 VDD.n1046 VDD.n1045 0.2705
R91998 VDD.n1047 VDD.n1046 0.2705
R91999 VDD.n1048 VDD.n1047 0.2705
R92000 VDD.n1049 VDD.n1048 0.2705
R92001 VDD.n1050 VDD.n1049 0.2705
R92002 VDD.n1051 VDD.n1050 0.2705
R92003 VDD.n1052 VDD.n1051 0.2705
R92004 VDD.n1053 VDD.n1052 0.2705
R92005 VDD.n1054 VDD.n1053 0.2705
R92006 VDD.n1055 VDD.n1054 0.2705
R92007 VDD.n1056 VDD.n1055 0.2705
R92008 VDD.n1057 VDD.n1056 0.2705
R92009 VDD.n1058 VDD.n1057 0.2705
R92010 VDD.n1059 VDD.n1058 0.2705
R92011 VDD.n1060 VDD.n1059 0.2705
R92012 VDD.n1061 VDD.n1060 0.2705
R92013 VDD.n1062 VDD.n1061 0.2705
R92014 VDD.n1063 VDD.n1062 0.2705
R92015 VDD.n1063 VDD.n273 0.2705
R92016 VDD.n1064 VDD.n281 0.2705
R92017 VDD.n1064 VDD.n274 0.2705
R92018 VDD.n1066 VDD.n1065 0.2705
R92019 VDD.n1065 VDD.n275 0.2705
R92020 VDD.n279 VDD.n278 0.2705
R92021 VDD.n278 VDD.n276 0.2705
R92022 VDD.n1071 VDD.n1070 0.2705
R92023 VDD.n1072 VDD.n1071 0.2705
R92024 VDD.n1084 VDD.n1083 0.2705
R92025 VDD.n500 VDD.n499 0.2705
R92026 VDD.n501 VDD.n500 0.2705
R92027 VDD.n502 VDD.n501 0.2705
R92028 VDD.n503 VDD.n502 0.2705
R92029 VDD.n504 VDD.n503 0.2705
R92030 VDD.n505 VDD.n504 0.2705
R92031 VDD.n506 VDD.n505 0.2705
R92032 VDD.n507 VDD.n506 0.2705
R92033 VDD.n508 VDD.n507 0.2705
R92034 VDD.n509 VDD.n508 0.2705
R92035 VDD.n510 VDD.n509 0.2705
R92036 VDD.n511 VDD.n510 0.2705
R92037 VDD.n512 VDD.n511 0.2705
R92038 VDD.n513 VDD.n512 0.2705
R92039 VDD.n514 VDD.n513 0.2705
R92040 VDD.n531 VDD.n514 0.2705
R92041 VDD.n531 VDD.n170 0.2705
R92042 VDD.n1128 VDD.n170 0.2705
R92043 VDD.n1128 VDD.n1127 0.2705
R92044 VDD.n174 VDD.n172 0.2705
R92045 VDD.n178 VDD.n176 0.2705
R92046 VDD.n182 VDD.n180 0.2705
R92047 VDD.n186 VDD.n184 0.2705
R92048 VDD.n190 VDD.n188 0.2705
R92049 VDD.n194 VDD.n192 0.2705
R92050 VDD.n198 VDD.n196 0.2705
R92051 VDD.n202 VDD.n200 0.2705
R92052 VDD.n204 VDD.n202 0.2705
R92053 VDD.n206 VDD.n204 0.2705
R92054 VDD.n208 VDD.n206 0.2705
R92055 VDD.n210 VDD.n208 0.2705
R92056 VDD.n212 VDD.n210 0.2705
R92057 VDD.n214 VDD.n212 0.2705
R92058 VDD.n216 VDD.n214 0.2705
R92059 VDD.n218 VDD.n216 0.2705
R92060 VDD.n220 VDD.n218 0.2705
R92061 VDD.n222 VDD.n220 0.2705
R92062 VDD.n224 VDD.n222 0.2705
R92063 VDD.n226 VDD.n224 0.2705
R92064 VDD.n228 VDD.n226 0.2705
R92065 VDD.n230 VDD.n228 0.2705
R92066 VDD.n232 VDD.n230 0.2705
R92067 VDD.n234 VDD.n232 0.2705
R92068 VDD.n236 VDD.n234 0.2705
R92069 VDD.n238 VDD.n236 0.2705
R92070 VDD.n259 VDD.n238 0.2705
R92071 VDD.n285 VDD.n281 0.248
R92072 VDD.n873 VDD.n566 0.248
R92073 VDD.n1069 VDD.n1068 0.241882
R92074 VDD.n1074 VDD.n1073 0.241882
R92075 VDD.n762 VDD.n761 0.237342
R92076 VDD.n490 VDD.n488 0.237342
R92077 VDD.n484 VDD.n482 0.237342
R92078 VDD.n474 VDD.n472 0.237342
R92079 VDD.n456 VDD.n454 0.237342
R92080 VDD.n446 VDD.n444 0.237342
R92081 VDD.n437 VDD.n436 0.237342
R92082 VDD.n423 VDD.n422 0.237342
R92083 VDD.n394 VDD.n393 0.237342
R92084 VDD.n948 VDD.n947 0.237342
R92085 VDD.n416 VDD.n415 0.237342
R92086 VDD.n430 VDD.n429 0.237342
R92087 VDD.n981 VDD.n980 0.228935
R92088 VDD.n799 VDD.n798 0.228935
R92089 VDD.n742 VDD.n663 0.227868
R92090 VDD.n481 VDD.n478 0.227868
R92091 VDD.n453 VDD.n450 0.227868
R92092 VDD.n1037 VDD.n1036 0.226
R92093 VDD.n550 VDD.n498 0.226
R92094 VDD.n851 VDD.n850 0.226
R92095 VDD.n879 VDD.n878 0.226
R92096 VDD.n261 VDD.n260 0.226
R92097 VDD.n880 VDD.n563 0.2255
R92098 VDD.n888 VDD.n555 0.2255
R92099 VDD.n889 VDD.n554 0.2255
R92100 VDD.n890 VDD.n553 0.2255
R92101 VDD.n891 VDD.n552 0.2255
R92102 VDD.n892 VDD.n497 0.2255
R92103 VDD.n887 VDD.n556 0.2255
R92104 VDD.n886 VDD.n557 0.2255
R92105 VDD.n885 VDD.n558 0.2255
R92106 VDD.n799 VDD.n638 0.2255
R92107 VDD.n884 VDD.n559 0.2255
R92108 VDD.n801 VDD.n800 0.2255
R92109 VDD.n883 VDD.n560 0.2255
R92110 VDD.n591 VDD.n590 0.2255
R92111 VDD.n882 VDD.n561 0.2255
R92112 VDD.n850 VDD.n849 0.2255
R92113 VDD.n881 VDD.n562 0.2255
R92114 VDD.n879 VDD.n564 0.2255
R92115 VDD.n550 VDD.n549 0.2255
R92116 VDD.n261 VDD.n239 0.2255
R92117 VDD.n551 VDD.n496 0.2255
R92118 VDD.n1090 VDD.n262 0.2255
R92119 VDD.n894 VDD.n893 0.2255
R92120 VDD.n1089 VDD.n1088 0.2255
R92121 VDD.n1083 VDD.n267 0.2255
R92122 VDD.n1082 VDD.n268 0.2255
R92123 VDD.n982 VDD.n981 0.2255
R92124 VDD.n1081 VDD.n269 0.2255
R92125 VDD.n332 VDD.n331 0.2255
R92126 VDD.n1080 VDD.n270 0.2255
R92127 VDD.n1035 VDD.n1034 0.2255
R92128 VDD.n1079 VDD.n271 0.2255
R92129 VDD.n1036 VDD.n330 0.2255
R92130 VDD.n1078 VDD.n272 0.2255
R92131 VDD.n1077 VDD.n273 0.2255
R92132 VDD.n1076 VDD.n274 0.2255
R92133 VDD.n1067 VDD.n1066 0.2255
R92134 VDD.n1075 VDD.n275 0.2255
R92135 VDD.n1068 VDD.n279 0.2255
R92136 VDD.n1074 VDD.n276 0.2255
R92137 VDD.n949 VDD.n407 0.223132
R92138 VDD.n426 VDD.n425 0.221947
R92139 VDD.n709 VDD.n402 0.218395
R92140 VDD.n408 VDD.n407 0.218395
R92141 VDD.n1037 VDD.n329 0.208
R92142 VDD.n515 VDD.n498 0.208
R92143 VDD.n852 VDD.n851 0.208
R92144 VDD.n260 VDD.n258 0.208
R92145 VDD.n722 VDD.n686 0.2075
R92146 VDD.n688 VDD.n417 0.2075
R92147 VDD.n689 VDD.n687 0.2075
R92148 VDD.n724 VDD.n723 0.2075
R92149 VDD.n428 VDD.n426 0.197079
R92150 VDD.n697 VDD.n396 0.194711
R92151 VDD.n947 VDD.n263 0.194711
R92152 VDD.n675 VDD.n422 0.192342
R92153 VDD.n668 VDD.n460 0.189974
R92154 VDD.n761 VDD.n760 0.189974
R92155 VDD.n760 VDD.n759 0.189974
R92156 VDD.n759 VDD.n758 0.189974
R92157 VDD.n758 VDD.n757 0.189974
R92158 VDD.n757 VDD.n756 0.189974
R92159 VDD.n756 VDD.n755 0.189974
R92160 VDD.n755 VDD.n754 0.189974
R92161 VDD.n754 VDD.n753 0.189974
R92162 VDD.n751 VDD.n750 0.189974
R92163 VDD.n750 VDD.n749 0.189974
R92164 VDD.n749 VDD.n748 0.189974
R92165 VDD.n748 VDD.n747 0.189974
R92166 VDD.n747 VDD.n746 0.189974
R92167 VDD.n746 VDD.n745 0.189974
R92168 VDD.n745 VDD.n744 0.189974
R92169 VDD.n744 VDD.n743 0.189974
R92170 VDD.n743 VDD.n742 0.189974
R92171 VDD.n768 VDD.n663 0.189974
R92172 VDD.n667 VDD.n666 0.189974
R92173 VDD.n478 VDD.n477 0.189974
R92174 VDD.n468 VDD.n466 0.189974
R92175 VDD.n450 VDD.n449 0.189974
R92176 VDD.n441 VDD.n440 0.189974
R92177 VDD.n741 VDD.n671 0.189974
R92178 VDD.n676 VDD.n675 0.189974
R92179 VDD.n716 VDD.n697 0.189974
R92180 VDD.n396 VDD.n395 0.189974
R92181 VDD.n384 VDD.n383 0.189974
R92182 VDD.n385 VDD.n384 0.189974
R92183 VDD.n386 VDD.n385 0.189974
R92184 VDD.n387 VDD.n386 0.189974
R92185 VDD.n729 VDD.n677 0.189974
R92186 VDD.n696 VDD.n695 0.189974
R92187 VDD.n711 VDD.n710 0.189974
R92188 VDD.n953 VDD.n402 0.189974
R92189 VDD.n707 VDD.n706 0.189974
R92190 VDD.n414 VDD.n413 0.189974
R92191 VDD.n689 VDD.n688 0.189974
R92192 VDD.n723 VDD.n722 0.189974
R92193 VDD.n735 VDD.n672 0.189974
R92194 VDD.n264 VDD.n263 0.189974
R92195 VDD.n266 VDD.n265 0.189974
R92196 VDD.n954 VDD.n953 0.189974
R92197 VDD.n671 VDD.n435 0.185
R92198 VDD.n1070 VDD.n279 0.1805
R92199 VDD.n1066 VDD.n279 0.1805
R92200 VDD.n1066 VDD.n281 0.1805
R92201 VDD.n1062 VDD.n281 0.1805
R92202 VDD.n1038 VDD.n330 0.1805
R92203 VDD.n1039 VDD.n328 0.1805
R92204 VDD.n1040 VDD.n326 0.1805
R92205 VDD.n1041 VDD.n324 0.1805
R92206 VDD.n1042 VDD.n322 0.1805
R92207 VDD.n1043 VDD.n320 0.1805
R92208 VDD.n1044 VDD.n318 0.1805
R92209 VDD.n1045 VDD.n316 0.1805
R92210 VDD.n1046 VDD.n314 0.1805
R92211 VDD.n1047 VDD.n312 0.1805
R92212 VDD.n1048 VDD.n310 0.1805
R92213 VDD.n1049 VDD.n308 0.1805
R92214 VDD.n1050 VDD.n306 0.1805
R92215 VDD.n1051 VDD.n304 0.1805
R92216 VDD.n1052 VDD.n302 0.1805
R92217 VDD.n1053 VDD.n300 0.1805
R92218 VDD.n1054 VDD.n298 0.1805
R92219 VDD.n1055 VDD.n296 0.1805
R92220 VDD.n1056 VDD.n294 0.1805
R92221 VDD.n1057 VDD.n292 0.1805
R92222 VDD.n1058 VDD.n290 0.1805
R92223 VDD.n1059 VDD.n288 0.1805
R92224 VDD.n1060 VDD.n286 0.1805
R92225 VDD.n1061 VDD.n284 0.1805
R92226 VDD.n1062 VDD.n283 0.1805
R92227 VDD.n1034 VDD.n330 0.1805
R92228 VDD.n1033 VDD.n328 0.1805
R92229 VDD.n1032 VDD.n326 0.1805
R92230 VDD.n1031 VDD.n324 0.1805
R92231 VDD.n1030 VDD.n322 0.1805
R92232 VDD.n1029 VDD.n320 0.1805
R92233 VDD.n1028 VDD.n318 0.1805
R92234 VDD.n1027 VDD.n316 0.1805
R92235 VDD.n1026 VDD.n314 0.1805
R92236 VDD.n1025 VDD.n312 0.1805
R92237 VDD.n1024 VDD.n310 0.1805
R92238 VDD.n1023 VDD.n308 0.1805
R92239 VDD.n1022 VDD.n306 0.1805
R92240 VDD.n1021 VDD.n304 0.1805
R92241 VDD.n1020 VDD.n302 0.1805
R92242 VDD.n1019 VDD.n300 0.1805
R92243 VDD.n1018 VDD.n298 0.1805
R92244 VDD.n1017 VDD.n296 0.1805
R92245 VDD.n1016 VDD.n294 0.1805
R92246 VDD.n1015 VDD.n292 0.1805
R92247 VDD.n1014 VDD.n290 0.1805
R92248 VDD.n1013 VDD.n288 0.1805
R92249 VDD.n1012 VDD.n286 0.1805
R92250 VDD.n1011 VDD.n284 0.1805
R92251 VDD.n1010 VDD.n283 0.1805
R92252 VDD.n1034 VDD.n332 0.1805
R92253 VDD.n1033 VDD.n333 0.1805
R92254 VDD.n1032 VDD.n334 0.1805
R92255 VDD.n1031 VDD.n335 0.1805
R92256 VDD.n1030 VDD.n336 0.1805
R92257 VDD.n1029 VDD.n337 0.1805
R92258 VDD.n1028 VDD.n338 0.1805
R92259 VDD.n1027 VDD.n339 0.1805
R92260 VDD.n1026 VDD.n340 0.1805
R92261 VDD.n1025 VDD.n341 0.1805
R92262 VDD.n1024 VDD.n342 0.1805
R92263 VDD.n1023 VDD.n343 0.1805
R92264 VDD.n1022 VDD.n344 0.1805
R92265 VDD.n1021 VDD.n345 0.1805
R92266 VDD.n1020 VDD.n346 0.1805
R92267 VDD.n1019 VDD.n347 0.1805
R92268 VDD.n1018 VDD.n348 0.1805
R92269 VDD.n1017 VDD.n349 0.1805
R92270 VDD.n1016 VDD.n350 0.1805
R92271 VDD.n1015 VDD.n351 0.1805
R92272 VDD.n1014 VDD.n352 0.1805
R92273 VDD.n1013 VDD.n353 0.1805
R92274 VDD.n1012 VDD.n354 0.1805
R92275 VDD.n1011 VDD.n355 0.1805
R92276 VDD.n1010 VDD.n356 0.1805
R92277 VDD.n982 VDD.n332 0.1805
R92278 VDD.n983 VDD.n333 0.1805
R92279 VDD.n984 VDD.n334 0.1805
R92280 VDD.n985 VDD.n335 0.1805
R92281 VDD.n986 VDD.n336 0.1805
R92282 VDD.n987 VDD.n337 0.1805
R92283 VDD.n988 VDD.n338 0.1805
R92284 VDD.n989 VDD.n339 0.1805
R92285 VDD.n990 VDD.n340 0.1805
R92286 VDD.n991 VDD.n341 0.1805
R92287 VDD.n992 VDD.n342 0.1805
R92288 VDD.n993 VDD.n343 0.1805
R92289 VDD.n994 VDD.n344 0.1805
R92290 VDD.n995 VDD.n345 0.1805
R92291 VDD.n996 VDD.n346 0.1805
R92292 VDD.n997 VDD.n347 0.1805
R92293 VDD.n998 VDD.n348 0.1805
R92294 VDD.n999 VDD.n349 0.1805
R92295 VDD.n1000 VDD.n350 0.1805
R92296 VDD.n1001 VDD.n351 0.1805
R92297 VDD.n1002 VDD.n352 0.1805
R92298 VDD.n1003 VDD.n353 0.1805
R92299 VDD.n1004 VDD.n354 0.1805
R92300 VDD.n1005 VDD.n355 0.1805
R92301 VDD.n1006 VDD.n356 0.1805
R92302 VDD.n982 VDD.n382 0.1805
R92303 VDD.n983 VDD.n381 0.1805
R92304 VDD.n984 VDD.n380 0.1805
R92305 VDD.n985 VDD.n379 0.1805
R92306 VDD.n986 VDD.n378 0.1805
R92307 VDD.n987 VDD.n377 0.1805
R92308 VDD.n988 VDD.n376 0.1805
R92309 VDD.n989 VDD.n375 0.1805
R92310 VDD.n990 VDD.n374 0.1805
R92311 VDD.n991 VDD.n373 0.1805
R92312 VDD.n992 VDD.n372 0.1805
R92313 VDD.n993 VDD.n371 0.1805
R92314 VDD.n994 VDD.n370 0.1805
R92315 VDD.n995 VDD.n369 0.1805
R92316 VDD.n996 VDD.n368 0.1805
R92317 VDD.n997 VDD.n367 0.1805
R92318 VDD.n998 VDD.n366 0.1805
R92319 VDD.n999 VDD.n365 0.1805
R92320 VDD.n1000 VDD.n364 0.1805
R92321 VDD.n1001 VDD.n363 0.1805
R92322 VDD.n1002 VDD.n362 0.1805
R92323 VDD.n1003 VDD.n361 0.1805
R92324 VDD.n1004 VDD.n360 0.1805
R92325 VDD.n1005 VDD.n359 0.1805
R92326 VDD.n1006 VDD.n358 0.1805
R92327 VDD.n1039 VDD.n329 0.1805
R92328 VDD.n1040 VDD.n327 0.1805
R92329 VDD.n1041 VDD.n325 0.1805
R92330 VDD.n1042 VDD.n323 0.1805
R92331 VDD.n1043 VDD.n321 0.1805
R92332 VDD.n1044 VDD.n319 0.1805
R92333 VDD.n1045 VDD.n317 0.1805
R92334 VDD.n1046 VDD.n315 0.1805
R92335 VDD.n1047 VDD.n313 0.1805
R92336 VDD.n1048 VDD.n311 0.1805
R92337 VDD.n1049 VDD.n309 0.1805
R92338 VDD.n1050 VDD.n307 0.1805
R92339 VDD.n1051 VDD.n305 0.1805
R92340 VDD.n1052 VDD.n303 0.1805
R92341 VDD.n1053 VDD.n301 0.1805
R92342 VDD.n1054 VDD.n299 0.1805
R92343 VDD.n1055 VDD.n297 0.1805
R92344 VDD.n1056 VDD.n295 0.1805
R92345 VDD.n1057 VDD.n293 0.1805
R92346 VDD.n1058 VDD.n291 0.1805
R92347 VDD.n1059 VDD.n289 0.1805
R92348 VDD.n1060 VDD.n287 0.1805
R92349 VDD.n1061 VDD.n285 0.1805
R92350 VDD.n978 VDD.n380 0.1805
R92351 VDD.n977 VDD.n379 0.1805
R92352 VDD.n976 VDD.n378 0.1805
R92353 VDD.n975 VDD.n377 0.1805
R92354 VDD.n974 VDD.n376 0.1805
R92355 VDD.n973 VDD.n375 0.1805
R92356 VDD.n972 VDD.n374 0.1805
R92357 VDD.n971 VDD.n373 0.1805
R92358 VDD.n970 VDD.n372 0.1805
R92359 VDD.n969 VDD.n371 0.1805
R92360 VDD.n968 VDD.n370 0.1805
R92361 VDD.n967 VDD.n369 0.1805
R92362 VDD.n966 VDD.n368 0.1805
R92363 VDD.n965 VDD.n367 0.1805
R92364 VDD.n964 VDD.n366 0.1805
R92365 VDD.n963 VDD.n365 0.1805
R92366 VDD.n962 VDD.n364 0.1805
R92367 VDD.n961 VDD.n363 0.1805
R92368 VDD.n960 VDD.n362 0.1805
R92369 VDD.n959 VDD.n361 0.1805
R92370 VDD.n958 VDD.n360 0.1805
R92371 VDD.n957 VDD.n359 0.1805
R92372 VDD.n956 VDD.n358 0.1805
R92373 VDD.n1090 VDD.n239 0.1805
R92374 VDD.n894 VDD.n496 0.1805
R92375 VDD.n895 VDD.n494 0.1805
R92376 VDD.n896 VDD.n492 0.1805
R92377 VDD.n897 VDD.n491 0.1805
R92378 VDD.n898 VDD.n489 0.1805
R92379 VDD.n899 VDD.n485 0.1805
R92380 VDD.n900 VDD.n483 0.1805
R92381 VDD.n901 VDD.n479 0.1805
R92382 VDD.n902 VDD.n475 0.1805
R92383 VDD.n903 VDD.n473 0.1805
R92384 VDD.n904 VDD.n469 0.1805
R92385 VDD.n905 VDD.n467 0.1805
R92386 VDD.n906 VDD.n463 0.1805
R92387 VDD.n907 VDD.n461 0.1805
R92388 VDD.n908 VDD.n457 0.1805
R92389 VDD.n909 VDD.n455 0.1805
R92390 VDD.n910 VDD.n451 0.1805
R92391 VDD.n911 VDD.n447 0.1805
R92392 VDD.n912 VDD.n445 0.1805
R92393 VDD.n913 VDD.n171 0.1805
R92394 VDD.n914 VDD.n173 0.1805
R92395 VDD.n915 VDD.n175 0.1805
R92396 VDD.n916 VDD.n177 0.1805
R92397 VDD.n917 VDD.n179 0.1805
R92398 VDD.n918 VDD.n181 0.1805
R92399 VDD.n919 VDD.n183 0.1805
R92400 VDD.n920 VDD.n185 0.1805
R92401 VDD.n921 VDD.n187 0.1805
R92402 VDD.n922 VDD.n189 0.1805
R92403 VDD.n923 VDD.n191 0.1805
R92404 VDD.n924 VDD.n193 0.1805
R92405 VDD.n925 VDD.n195 0.1805
R92406 VDD.n926 VDD.n197 0.1805
R92407 VDD.n927 VDD.n199 0.1805
R92408 VDD.n928 VDD.n201 0.1805
R92409 VDD.n929 VDD.n203 0.1805
R92410 VDD.n930 VDD.n205 0.1805
R92411 VDD.n931 VDD.n207 0.1805
R92412 VDD.n932 VDD.n209 0.1805
R92413 VDD.n933 VDD.n211 0.1805
R92414 VDD.n934 VDD.n213 0.1805
R92415 VDD.n935 VDD.n215 0.1805
R92416 VDD.n936 VDD.n217 0.1805
R92417 VDD.n937 VDD.n219 0.1805
R92418 VDD.n938 VDD.n221 0.1805
R92419 VDD.n939 VDD.n223 0.1805
R92420 VDD.n940 VDD.n225 0.1805
R92421 VDD.n941 VDD.n227 0.1805
R92422 VDD.n942 VDD.n229 0.1805
R92423 VDD.n943 VDD.n231 0.1805
R92424 VDD.n944 VDD.n233 0.1805
R92425 VDD.n945 VDD.n235 0.1805
R92426 VDD.n946 VDD.n237 0.1805
R92427 VDD.n1092 VDD.n238 0.1805
R92428 VDD.n170 VDD.n159 0.1805
R92429 VDD.n531 VDD.n530 0.1805
R92430 VDD.n529 VDD.n514 0.1805
R92431 VDD.n528 VDD.n513 0.1805
R92432 VDD.n527 VDD.n512 0.1805
R92433 VDD.n526 VDD.n511 0.1805
R92434 VDD.n525 VDD.n510 0.1805
R92435 VDD.n524 VDD.n509 0.1805
R92436 VDD.n523 VDD.n508 0.1805
R92437 VDD.n522 VDD.n507 0.1805
R92438 VDD.n521 VDD.n506 0.1805
R92439 VDD.n520 VDD.n505 0.1805
R92440 VDD.n519 VDD.n504 0.1805
R92441 VDD.n518 VDD.n503 0.1805
R92442 VDD.n517 VDD.n502 0.1805
R92443 VDD.n516 VDD.n501 0.1805
R92444 VDD.n515 VDD.n500 0.1805
R92445 VDD.n877 VDD.n564 0.1805
R92446 VDD.n875 VDD.n566 0.1805
R92447 VDD.n563 VDD.n562 0.1805
R92448 VDD.n564 VDD.n563 0.1805
R92449 VDD.n614 VDD.n566 0.1805
R92450 VDD.n873 VDD.n567 0.1805
R92451 VDD.n872 VDD.n568 0.1805
R92452 VDD.n871 VDD.n569 0.1805
R92453 VDD.n870 VDD.n570 0.1805
R92454 VDD.n869 VDD.n571 0.1805
R92455 VDD.n868 VDD.n572 0.1805
R92456 VDD.n867 VDD.n573 0.1805
R92457 VDD.n866 VDD.n574 0.1805
R92458 VDD.n865 VDD.n575 0.1805
R92459 VDD.n864 VDD.n576 0.1805
R92460 VDD.n863 VDD.n577 0.1805
R92461 VDD.n862 VDD.n578 0.1805
R92462 VDD.n861 VDD.n579 0.1805
R92463 VDD.n860 VDD.n580 0.1805
R92464 VDD.n859 VDD.n581 0.1805
R92465 VDD.n858 VDD.n582 0.1805
R92466 VDD.n857 VDD.n583 0.1805
R92467 VDD.n856 VDD.n584 0.1805
R92468 VDD.n855 VDD.n585 0.1805
R92469 VDD.n854 VDD.n586 0.1805
R92470 VDD.n853 VDD.n587 0.1805
R92471 VDD.n562 VDD.n561 0.1805
R92472 VDD.n826 VDD.n614 0.1805
R92473 VDD.n827 VDD.n567 0.1805
R92474 VDD.n828 VDD.n568 0.1805
R92475 VDD.n829 VDD.n569 0.1805
R92476 VDD.n830 VDD.n570 0.1805
R92477 VDD.n831 VDD.n571 0.1805
R92478 VDD.n832 VDD.n572 0.1805
R92479 VDD.n833 VDD.n573 0.1805
R92480 VDD.n834 VDD.n574 0.1805
R92481 VDD.n835 VDD.n575 0.1805
R92482 VDD.n836 VDD.n576 0.1805
R92483 VDD.n837 VDD.n577 0.1805
R92484 VDD.n838 VDD.n578 0.1805
R92485 VDD.n839 VDD.n579 0.1805
R92486 VDD.n840 VDD.n580 0.1805
R92487 VDD.n841 VDD.n581 0.1805
R92488 VDD.n842 VDD.n582 0.1805
R92489 VDD.n843 VDD.n583 0.1805
R92490 VDD.n844 VDD.n584 0.1805
R92491 VDD.n845 VDD.n585 0.1805
R92492 VDD.n846 VDD.n586 0.1805
R92493 VDD.n847 VDD.n587 0.1805
R92494 VDD.n561 VDD.n560 0.1805
R92495 VDD.n826 VDD.n825 0.1805
R92496 VDD.n827 VDD.n613 0.1805
R92497 VDD.n828 VDD.n612 0.1805
R92498 VDD.n829 VDD.n611 0.1805
R92499 VDD.n830 VDD.n610 0.1805
R92500 VDD.n831 VDD.n609 0.1805
R92501 VDD.n832 VDD.n608 0.1805
R92502 VDD.n833 VDD.n607 0.1805
R92503 VDD.n834 VDD.n606 0.1805
R92504 VDD.n835 VDD.n605 0.1805
R92505 VDD.n836 VDD.n604 0.1805
R92506 VDD.n837 VDD.n603 0.1805
R92507 VDD.n838 VDD.n602 0.1805
R92508 VDD.n839 VDD.n601 0.1805
R92509 VDD.n840 VDD.n600 0.1805
R92510 VDD.n841 VDD.n599 0.1805
R92511 VDD.n842 VDD.n598 0.1805
R92512 VDD.n843 VDD.n597 0.1805
R92513 VDD.n844 VDD.n596 0.1805
R92514 VDD.n845 VDD.n595 0.1805
R92515 VDD.n846 VDD.n594 0.1805
R92516 VDD.n847 VDD.n593 0.1805
R92517 VDD.n560 VDD.n559 0.1805
R92518 VDD.n825 VDD.n824 0.1805
R92519 VDD.n823 VDD.n613 0.1805
R92520 VDD.n822 VDD.n612 0.1805
R92521 VDD.n821 VDD.n611 0.1805
R92522 VDD.n820 VDD.n610 0.1805
R92523 VDD.n819 VDD.n609 0.1805
R92524 VDD.n818 VDD.n608 0.1805
R92525 VDD.n817 VDD.n607 0.1805
R92526 VDD.n816 VDD.n606 0.1805
R92527 VDD.n815 VDD.n605 0.1805
R92528 VDD.n814 VDD.n604 0.1805
R92529 VDD.n813 VDD.n603 0.1805
R92530 VDD.n812 VDD.n602 0.1805
R92531 VDD.n811 VDD.n601 0.1805
R92532 VDD.n810 VDD.n600 0.1805
R92533 VDD.n809 VDD.n599 0.1805
R92534 VDD.n808 VDD.n598 0.1805
R92535 VDD.n807 VDD.n597 0.1805
R92536 VDD.n806 VDD.n596 0.1805
R92537 VDD.n805 VDD.n595 0.1805
R92538 VDD.n804 VDD.n594 0.1805
R92539 VDD.n803 VDD.n593 0.1805
R92540 VDD.n559 VDD.n558 0.1805
R92541 VDD.n824 VDD.n615 0.1805
R92542 VDD.n823 VDD.n616 0.1805
R92543 VDD.n822 VDD.n617 0.1805
R92544 VDD.n821 VDD.n618 0.1805
R92545 VDD.n820 VDD.n619 0.1805
R92546 VDD.n819 VDD.n620 0.1805
R92547 VDD.n818 VDD.n621 0.1805
R92548 VDD.n817 VDD.n622 0.1805
R92549 VDD.n816 VDD.n623 0.1805
R92550 VDD.n815 VDD.n624 0.1805
R92551 VDD.n814 VDD.n625 0.1805
R92552 VDD.n813 VDD.n626 0.1805
R92553 VDD.n812 VDD.n627 0.1805
R92554 VDD.n811 VDD.n628 0.1805
R92555 VDD.n810 VDD.n629 0.1805
R92556 VDD.n809 VDD.n630 0.1805
R92557 VDD.n808 VDD.n631 0.1805
R92558 VDD.n807 VDD.n632 0.1805
R92559 VDD.n806 VDD.n633 0.1805
R92560 VDD.n805 VDD.n634 0.1805
R92561 VDD.n804 VDD.n635 0.1805
R92562 VDD.n803 VDD.n636 0.1805
R92563 VDD.n558 VDD.n557 0.1805
R92564 VDD.n774 VDD.n615 0.1805
R92565 VDD.n775 VDD.n616 0.1805
R92566 VDD.n776 VDD.n617 0.1805
R92567 VDD.n777 VDD.n618 0.1805
R92568 VDD.n778 VDD.n619 0.1805
R92569 VDD.n779 VDD.n620 0.1805
R92570 VDD.n780 VDD.n621 0.1805
R92571 VDD.n781 VDD.n622 0.1805
R92572 VDD.n782 VDD.n623 0.1805
R92573 VDD.n783 VDD.n624 0.1805
R92574 VDD.n784 VDD.n625 0.1805
R92575 VDD.n785 VDD.n626 0.1805
R92576 VDD.n786 VDD.n627 0.1805
R92577 VDD.n787 VDD.n628 0.1805
R92578 VDD.n788 VDD.n629 0.1805
R92579 VDD.n789 VDD.n630 0.1805
R92580 VDD.n790 VDD.n631 0.1805
R92581 VDD.n791 VDD.n632 0.1805
R92582 VDD.n792 VDD.n633 0.1805
R92583 VDD.n793 VDD.n634 0.1805
R92584 VDD.n794 VDD.n635 0.1805
R92585 VDD.n795 VDD.n636 0.1805
R92586 VDD.n557 VDD.n556 0.1805
R92587 VDD.n774 VDD.n773 0.1805
R92588 VDD.n775 VDD.n660 0.1805
R92589 VDD.n777 VDD.n658 0.1805
R92590 VDD.n778 VDD.n657 0.1805
R92591 VDD.n779 VDD.n656 0.1805
R92592 VDD.n780 VDD.n655 0.1805
R92593 VDD.n781 VDD.n654 0.1805
R92594 VDD.n782 VDD.n653 0.1805
R92595 VDD.n783 VDD.n652 0.1805
R92596 VDD.n784 VDD.n651 0.1805
R92597 VDD.n785 VDD.n650 0.1805
R92598 VDD.n786 VDD.n649 0.1805
R92599 VDD.n787 VDD.n648 0.1805
R92600 VDD.n788 VDD.n647 0.1805
R92601 VDD.n789 VDD.n646 0.1805
R92602 VDD.n790 VDD.n645 0.1805
R92603 VDD.n791 VDD.n644 0.1805
R92604 VDD.n792 VDD.n643 0.1805
R92605 VDD.n793 VDD.n642 0.1805
R92606 VDD.n794 VDD.n641 0.1805
R92607 VDD.n795 VDD.n640 0.1805
R92608 VDD.n922 VDD.n431 0.1805
R92609 VDD.n894 VDD.n497 0.1805
R92610 VDD.n895 VDD.n495 0.1805
R92611 VDD.n552 VDD.n497 0.1805
R92612 VDD.n664 VDD.n495 0.1805
R92613 VDD.n553 VDD.n552 0.1805
R92614 VDD.n664 VDD.n662 0.1805
R92615 VDD.n554 VDD.n553 0.1805
R92616 VDD.n773 VDD.n772 0.1805
R92617 VDD.n555 VDD.n554 0.1805
R92618 VDD.n556 VDD.n555 0.1805
R92619 VDD.n770 VDD.n661 0.1805
R92620 VDD.n661 VDD.n660 0.1805
R92621 VDD.n771 VDD.n662 0.1805
R92622 VDD.n772 VDD.n771 0.1805
R92623 VDD.n769 VDD.n665 0.1805
R92624 VDD.n770 VDD.n769 0.1805
R92625 VDD.n896 VDD.n493 0.1805
R92626 VDD.n665 VDD.n493 0.1805
R92627 VDD.n918 VDD.n435 0.1805
R92628 VDD.n740 VDD.n435 0.1805
R92629 VDD.n919 VDD.n434 0.1805
R92630 VDD.n739 VDD.n434 0.1805
R92631 VDD.n920 VDD.n433 0.1805
R92632 VDD.n738 VDD.n433 0.1805
R92633 VDD.n921 VDD.n432 0.1805
R92634 VDD.n737 VDD.n432 0.1805
R92635 VDD.n728 VDD.n678 0.1805
R92636 VDD.n727 VDD.n680 0.1805
R92637 VDD.n726 VDD.n682 0.1805
R92638 VDD.n725 VDD.n684 0.1805
R92639 VDD.n934 VDD.n417 0.1805
R92640 VDD.n930 VDD.n421 0.1805
R92641 VDD.n678 VDD.n421 0.1805
R92642 VDD.n931 VDD.n420 0.1805
R92643 VDD.n680 VDD.n420 0.1805
R92644 VDD.n932 VDD.n419 0.1805
R92645 VDD.n682 VDD.n419 0.1805
R92646 VDD.n933 VDD.n418 0.1805
R92647 VDD.n684 VDD.n418 0.1805
R92648 VDD.n940 VDD.n412 0.1805
R92649 VDD.n941 VDD.n411 0.1805
R92650 VDD.n942 VDD.n410 0.1805
R92651 VDD.n943 VDD.n409 0.1805
R92652 VDD.n958 VDD.n401 0.1805
R92653 VDD.n962 VDD.n397 0.1805
R92654 VDD.n961 VDD.n398 0.1805
R92655 VDD.n960 VDD.n399 0.1805
R92656 VDD.n698 VDD.n397 0.1805
R92657 VDD.n700 VDD.n398 0.1805
R92658 VDD.n702 VDD.n399 0.1805
R92659 VDD.n715 VDD.n698 0.1805
R92660 VDD.n714 VDD.n700 0.1805
R92661 VDD.n713 VDD.n702 0.1805
R92662 VDD.n704 VDD.n409 0.1805
R92663 VDD.n728 VDD.n679 0.1805
R92664 VDD.n727 VDD.n681 0.1805
R92665 VDD.n726 VDD.n683 0.1805
R92666 VDD.n725 VDD.n685 0.1805
R92667 VDD.n968 VDD.n392 0.1805
R92668 VDD.n679 VDD.n388 0.1805
R92669 VDD.n972 VDD.n388 0.1805
R92670 VDD.n681 VDD.n389 0.1805
R92671 VDD.n971 VDD.n389 0.1805
R92672 VDD.n683 VDD.n390 0.1805
R92673 VDD.n970 VDD.n390 0.1805
R92674 VDD.n685 VDD.n391 0.1805
R92675 VDD.n969 VDD.n391 0.1805
R92676 VDD.n724 VDD.n686 0.1805
R92677 VDD.n686 VDD.n392 0.1805
R92678 VDD.n699 VDD.n412 0.1805
R92679 VDD.n715 VDD.n699 0.1805
R92680 VDD.n701 VDD.n411 0.1805
R92681 VDD.n714 VDD.n701 0.1805
R92682 VDD.n703 VDD.n410 0.1805
R92683 VDD.n713 VDD.n703 0.1805
R92684 VDD.n712 VDD.n704 0.1805
R92685 VDD.n712 VDD.n705 0.1805
R92686 VDD.n705 VDD.n400 0.1805
R92687 VDD.n959 VDD.n400 0.1805
R92688 VDD.n687 VDD.n417 0.1805
R92689 VDD.n724 VDD.n687 0.1805
R92690 VDD.n736 VDD.n431 0.1805
R92691 VDD.n796 VDD.n639 0.1805
R92692 VDD.n776 VDD.n659 0.1805
R92693 VDD.n797 VDD.n638 0.1805
R92694 VDD.n796 VDD.n637 0.1805
R92695 VDD.n802 VDD.n637 0.1805
R92696 VDD.n801 VDD.n638 0.1805
R92697 VDD.n801 VDD.n591 0.1805
R92698 VDD.n802 VDD.n592 0.1805
R92699 VDD.n848 VDD.n592 0.1805
R92700 VDD.n849 VDD.n591 0.1805
R92701 VDD.n849 VDD.n589 0.1805
R92702 VDD.n848 VDD.n588 0.1805
R92703 VDD.n852 VDD.n588 0.1805
R92704 VDD.n876 VDD.n875 0.1805
R92705 VDD.n549 VDD.n499 0.1805
R92706 VDD.n549 VDD.n496 0.1805
R92707 VDD.n548 VDD.n500 0.1805
R92708 VDD.n548 VDD.n494 0.1805
R92709 VDD.n547 VDD.n501 0.1805
R92710 VDD.n547 VDD.n492 0.1805
R92711 VDD.n546 VDD.n502 0.1805
R92712 VDD.n546 VDD.n491 0.1805
R92713 VDD.n545 VDD.n503 0.1805
R92714 VDD.n545 VDD.n489 0.1805
R92715 VDD.n544 VDD.n504 0.1805
R92716 VDD.n544 VDD.n485 0.1805
R92717 VDD.n543 VDD.n505 0.1805
R92718 VDD.n543 VDD.n483 0.1805
R92719 VDD.n542 VDD.n506 0.1805
R92720 VDD.n542 VDD.n479 0.1805
R92721 VDD.n541 VDD.n507 0.1805
R92722 VDD.n541 VDD.n475 0.1805
R92723 VDD.n540 VDD.n508 0.1805
R92724 VDD.n540 VDD.n473 0.1805
R92725 VDD.n539 VDD.n509 0.1805
R92726 VDD.n539 VDD.n469 0.1805
R92727 VDD.n538 VDD.n510 0.1805
R92728 VDD.n538 VDD.n467 0.1805
R92729 VDD.n537 VDD.n511 0.1805
R92730 VDD.n537 VDD.n463 0.1805
R92731 VDD.n536 VDD.n512 0.1805
R92732 VDD.n536 VDD.n461 0.1805
R92733 VDD.n535 VDD.n513 0.1805
R92734 VDD.n535 VDD.n457 0.1805
R92735 VDD.n534 VDD.n514 0.1805
R92736 VDD.n534 VDD.n455 0.1805
R92737 VDD.n533 VDD.n531 0.1805
R92738 VDD.n533 VDD.n451 0.1805
R92739 VDD.n532 VDD.n170 0.1805
R92740 VDD.n532 VDD.n447 0.1805
R92741 VDD.n1128 VDD.n169 0.1805
R92742 VDD.n445 VDD.n169 0.1805
R92743 VDD.n1127 VDD.n1126 0.1805
R92744 VDD.n1126 VDD.n171 0.1805
R92745 VDD.n1125 VDD.n172 0.1805
R92746 VDD.n1125 VDD.n173 0.1805
R92747 VDD.n1124 VDD.n174 0.1805
R92748 VDD.n1124 VDD.n175 0.1805
R92749 VDD.n1123 VDD.n176 0.1805
R92750 VDD.n1123 VDD.n177 0.1805
R92751 VDD.n1122 VDD.n178 0.1805
R92752 VDD.n1122 VDD.n179 0.1805
R92753 VDD.n1121 VDD.n180 0.1805
R92754 VDD.n1121 VDD.n181 0.1805
R92755 VDD.n1120 VDD.n182 0.1805
R92756 VDD.n1120 VDD.n183 0.1805
R92757 VDD.n1119 VDD.n184 0.1805
R92758 VDD.n1119 VDD.n185 0.1805
R92759 VDD.n1118 VDD.n186 0.1805
R92760 VDD.n1118 VDD.n187 0.1805
R92761 VDD.n1117 VDD.n188 0.1805
R92762 VDD.n1117 VDD.n189 0.1805
R92763 VDD.n1116 VDD.n190 0.1805
R92764 VDD.n1116 VDD.n191 0.1805
R92765 VDD.n1115 VDD.n192 0.1805
R92766 VDD.n1115 VDD.n193 0.1805
R92767 VDD.n1114 VDD.n194 0.1805
R92768 VDD.n1114 VDD.n195 0.1805
R92769 VDD.n1113 VDD.n196 0.1805
R92770 VDD.n1113 VDD.n197 0.1805
R92771 VDD.n1112 VDD.n198 0.1805
R92772 VDD.n1112 VDD.n199 0.1805
R92773 VDD.n1111 VDD.n200 0.1805
R92774 VDD.n1111 VDD.n201 0.1805
R92775 VDD.n1110 VDD.n202 0.1805
R92776 VDD.n1110 VDD.n203 0.1805
R92777 VDD.n1109 VDD.n204 0.1805
R92778 VDD.n1109 VDD.n205 0.1805
R92779 VDD.n1108 VDD.n206 0.1805
R92780 VDD.n1108 VDD.n207 0.1805
R92781 VDD.n1107 VDD.n208 0.1805
R92782 VDD.n1107 VDD.n209 0.1805
R92783 VDD.n1106 VDD.n210 0.1805
R92784 VDD.n1106 VDD.n211 0.1805
R92785 VDD.n1105 VDD.n212 0.1805
R92786 VDD.n1105 VDD.n213 0.1805
R92787 VDD.n1104 VDD.n214 0.1805
R92788 VDD.n1104 VDD.n215 0.1805
R92789 VDD.n1103 VDD.n216 0.1805
R92790 VDD.n1103 VDD.n217 0.1805
R92791 VDD.n1102 VDD.n218 0.1805
R92792 VDD.n1102 VDD.n219 0.1805
R92793 VDD.n1101 VDD.n220 0.1805
R92794 VDD.n1101 VDD.n221 0.1805
R92795 VDD.n1100 VDD.n222 0.1805
R92796 VDD.n1100 VDD.n223 0.1805
R92797 VDD.n1099 VDD.n224 0.1805
R92798 VDD.n1099 VDD.n225 0.1805
R92799 VDD.n1098 VDD.n226 0.1805
R92800 VDD.n1098 VDD.n227 0.1805
R92801 VDD.n1097 VDD.n228 0.1805
R92802 VDD.n1097 VDD.n229 0.1805
R92803 VDD.n1096 VDD.n230 0.1805
R92804 VDD.n1096 VDD.n231 0.1805
R92805 VDD.n1095 VDD.n232 0.1805
R92806 VDD.n1095 VDD.n233 0.1805
R92807 VDD.n1094 VDD.n234 0.1805
R92808 VDD.n1094 VDD.n235 0.1805
R92809 VDD.n1093 VDD.n236 0.1805
R92810 VDD.n1093 VDD.n237 0.1805
R92811 VDD.n1092 VDD.n1091 0.1805
R92812 VDD.n1091 VDD.n240 0.1805
R92813 VDD.n1090 VDD.n1089 0.1805
R92814 VDD.n955 VDD.n357 0.1805
R92815 VDD.n979 VDD.n381 0.1805
R92816 VDD.n268 VDD.n267 0.1805
R92817 VDD.n269 VDD.n268 0.1805
R92818 VDD.n1007 VDD.n357 0.1805
R92819 VDD.n1008 VDD.n1007 0.1805
R92820 VDD.n270 VDD.n269 0.1805
R92821 VDD.n271 VDD.n270 0.1805
R92822 VDD.n1009 VDD.n1008 0.1805
R92823 VDD.n1009 VDD.n282 0.1805
R92824 VDD.n272 VDD.n271 0.1805
R92825 VDD.n273 VDD.n272 0.1805
R92826 VDD.n1063 VDD.n282 0.1805
R92827 VDD.n1064 VDD.n1063 0.1805
R92828 VDD.n274 VDD.n273 0.1805
R92829 VDD.n275 VDD.n274 0.1805
R92830 VDD.n1065 VDD.n1064 0.1805
R92831 VDD.n1065 VDD.n278 0.1805
R92832 VDD.n276 VDD.n275 0.1805
R92833 VDD.n1072 VDD.n276 0.1805
R92834 VDD.n1071 VDD.n278 0.1805
R92835 VDD.n1071 VDD.n277 0.1805
R92836 VDD.n258 VDD.n238 0.1805
R92837 VDD.n257 VDD.n236 0.1805
R92838 VDD.n256 VDD.n234 0.1805
R92839 VDD.n255 VDD.n232 0.1805
R92840 VDD.n254 VDD.n230 0.1805
R92841 VDD.n253 VDD.n228 0.1805
R92842 VDD.n252 VDD.n226 0.1805
R92843 VDD.n251 VDD.n224 0.1805
R92844 VDD.n250 VDD.n222 0.1805
R92845 VDD.n249 VDD.n220 0.1805
R92846 VDD.n248 VDD.n218 0.1805
R92847 VDD.n247 VDD.n216 0.1805
R92848 VDD.n246 VDD.n214 0.1805
R92849 VDD.n245 VDD.n212 0.1805
R92850 VDD.n244 VDD.n210 0.1805
R92851 VDD.n243 VDD.n208 0.1805
R92852 VDD.n242 VDD.n206 0.1805
R92853 VDD.n241 VDD.n204 0.1805
R92854 VDD.n202 VDD.n160 0.1805
R92855 VDD.n259 VDD.n239 0.1805
R92856 VDD.n1129 VDD.n1128 0.1805
R92857 VDD.n1131 VDD.n1130 0.175505
R92858 VDD.n487 VDD.n484 0.171026
R92859 VDD.n459 VDD.n456 0.171026
R92860 VDD.n672 VDD.n430 0.168658
R92861 VDD.n741 VDD.n740 0.1625
R92862 VDD.n722 VDD.n393 0.156816
R92863 VDD.n753 VDD.n752 0.142605
R92864 VDD.n666 VDD.n490 0.142605
R92865 VDD.n767 VDD.n667 0.137868
R92866 VDD.n708 VDD.n707 0.137868
R92867 VDD.n735 VDD.n734 0.137868
R92868 VDD.n693 VDD.n394 0.137868
R92869 VDD.n717 VDD.n696 0.137868
R92870 VDD.n691 VDD.n415 0.137868
R92871 VDD.n721 VDD.n689 0.137868
R92872 VDD.n730 VDD.n676 0.137868
R92873 VDD.n763 VDD.n741 0.137868
R92874 VDD.n404 VDD.n264 0.137868
R92875 VDD.n1068 VDD.n1067 0.1355
R92876 VDD.n329 VDD.n327 0.1355
R92877 VDD.n327 VDD.n325 0.1355
R92878 VDD.n325 VDD.n323 0.1355
R92879 VDD.n323 VDD.n321 0.1355
R92880 VDD.n321 VDD.n319 0.1355
R92881 VDD.n319 VDD.n317 0.1355
R92882 VDD.n317 VDD.n315 0.1355
R92883 VDD.n315 VDD.n313 0.1355
R92884 VDD.n313 VDD.n311 0.1355
R92885 VDD.n311 VDD.n309 0.1355
R92886 VDD.n309 VDD.n307 0.1355
R92887 VDD.n307 VDD.n305 0.1355
R92888 VDD.n305 VDD.n303 0.1355
R92889 VDD.n303 VDD.n301 0.1355
R92890 VDD.n301 VDD.n299 0.1355
R92891 VDD.n299 VDD.n297 0.1355
R92892 VDD.n297 VDD.n295 0.1355
R92893 VDD.n295 VDD.n293 0.1355
R92894 VDD.n293 VDD.n291 0.1355
R92895 VDD.n291 VDD.n289 0.1355
R92896 VDD.n289 VDD.n287 0.1355
R92897 VDD.n981 VDD.n331 0.1355
R92898 VDD.n1035 VDD.n331 0.1355
R92899 VDD.n1036 VDD.n1035 0.1355
R92900 VDD.n516 VDD.n515 0.1355
R92901 VDD.n517 VDD.n516 0.1355
R92902 VDD.n518 VDD.n517 0.1355
R92903 VDD.n519 VDD.n518 0.1355
R92904 VDD.n520 VDD.n519 0.1355
R92905 VDD.n521 VDD.n520 0.1355
R92906 VDD.n522 VDD.n521 0.1355
R92907 VDD.n523 VDD.n522 0.1355
R92908 VDD.n524 VDD.n523 0.1355
R92909 VDD.n525 VDD.n524 0.1355
R92910 VDD.n526 VDD.n525 0.1355
R92911 VDD.n527 VDD.n526 0.1355
R92912 VDD.n528 VDD.n527 0.1355
R92913 VDD.n529 VDD.n528 0.1355
R92914 VDD.n530 VDD.n529 0.1355
R92915 VDD.n530 VDD.n159 0.1355
R92916 VDD.n800 VDD.n799 0.1355
R92917 VDD.n800 VDD.n590 0.1355
R92918 VDD.n850 VDD.n590 0.1355
R92919 VDD.n740 VDD.n739 0.1355
R92920 VDD.n739 VDD.n738 0.1355
R92921 VDD.n738 VDD.n737 0.1355
R92922 VDD.n737 VDD.n736 0.1355
R92923 VDD.n873 VDD.n872 0.1355
R92924 VDD.n872 VDD.n871 0.1355
R92925 VDD.n871 VDD.n870 0.1355
R92926 VDD.n870 VDD.n869 0.1355
R92927 VDD.n869 VDD.n868 0.1355
R92928 VDD.n868 VDD.n867 0.1355
R92929 VDD.n867 VDD.n866 0.1355
R92930 VDD.n866 VDD.n865 0.1355
R92931 VDD.n865 VDD.n864 0.1355
R92932 VDD.n864 VDD.n863 0.1355
R92933 VDD.n863 VDD.n862 0.1355
R92934 VDD.n862 VDD.n861 0.1355
R92935 VDD.n861 VDD.n860 0.1355
R92936 VDD.n860 VDD.n859 0.1355
R92937 VDD.n859 VDD.n858 0.1355
R92938 VDD.n858 VDD.n857 0.1355
R92939 VDD.n857 VDD.n856 0.1355
R92940 VDD.n856 VDD.n855 0.1355
R92941 VDD.n855 VDD.n854 0.1355
R92942 VDD.n854 VDD.n853 0.1355
R92943 VDD.n853 VDD.n852 0.1355
R92944 VDD.n551 VDD.n550 0.1355
R92945 VDD.n893 VDD.n551 0.1355
R92946 VDD.n893 VDD.n892 0.1355
R92947 VDD.n892 VDD.n891 0.1355
R92948 VDD.n891 VDD.n890 0.1355
R92949 VDD.n890 VDD.n889 0.1355
R92950 VDD.n889 VDD.n888 0.1355
R92951 VDD.n888 VDD.n887 0.1355
R92952 VDD.n887 VDD.n886 0.1355
R92953 VDD.n886 VDD.n885 0.1355
R92954 VDD.n885 VDD.n884 0.1355
R92955 VDD.n884 VDD.n883 0.1355
R92956 VDD.n883 VDD.n882 0.1355
R92957 VDD.n882 VDD.n881 0.1355
R92958 VDD.n881 VDD.n880 0.1355
R92959 VDD.n880 VDD.n879 0.1355
R92960 VDD.n262 VDD.n261 0.1355
R92961 VDD.n1088 VDD.n262 0.1355
R92962 VDD.n1088 VDD.n1087 0.1355
R92963 VDD.n1087 VDD.n1086 0.1355
R92964 VDD.n1086 VDD.n1085 0.1355
R92965 VDD.n1085 VDD.n1084 0.1355
R92966 VDD.n1083 VDD.n1082 0.1355
R92967 VDD.n1082 VDD.n1081 0.1355
R92968 VDD.n1081 VDD.n1080 0.1355
R92969 VDD.n1080 VDD.n1079 0.1355
R92970 VDD.n1079 VDD.n1078 0.1355
R92971 VDD.n1078 VDD.n1077 0.1355
R92972 VDD.n1077 VDD.n1076 0.1355
R92973 VDD.n1076 VDD.n1075 0.1355
R92974 VDD.n1075 VDD.n1074 0.1355
R92975 VDD.n241 VDD.n160 0.1355
R92976 VDD.n242 VDD.n241 0.1355
R92977 VDD.n243 VDD.n242 0.1355
R92978 VDD.n244 VDD.n243 0.1355
R92979 VDD.n245 VDD.n244 0.1355
R92980 VDD.n246 VDD.n245 0.1355
R92981 VDD.n247 VDD.n246 0.1355
R92982 VDD.n248 VDD.n247 0.1355
R92983 VDD.n249 VDD.n248 0.1355
R92984 VDD.n250 VDD.n249 0.1355
R92985 VDD.n251 VDD.n250 0.1355
R92986 VDD.n252 VDD.n251 0.1355
R92987 VDD.n253 VDD.n252 0.1355
R92988 VDD.n254 VDD.n253 0.1355
R92989 VDD.n255 VDD.n254 0.1355
R92990 VDD.n256 VDD.n255 0.1355
R92991 VDD.n257 VDD.n256 0.1355
R92992 VDD.n258 VDD.n257 0.1355
R92993 VDD.n898 VDD.n490 0.13325
R92994 VDD.n900 VDD.n484 0.13325
R92995 VDD.n902 VDD.n478 0.13325
R92996 VDD.n904 VDD.n472 0.13325
R92997 VDD.n905 VDD.n468 0.13325
R92998 VDD.n906 VDD.n466 0.13325
R92999 VDD.n907 VDD.n462 0.13325
R93000 VDD.n909 VDD.n456 0.13325
R93001 VDD.n911 VDD.n450 0.13325
R93002 VDD.n913 VDD.n444 0.13325
R93003 VDD.n914 VDD.n441 0.13325
R93004 VDD.n915 VDD.n440 0.13325
R93005 VDD.n916 VDD.n437 0.13325
R93006 VDD.n928 VDD.n422 0.13325
R93007 VDD.n945 VDD.n407 0.13325
R93008 VDD.n938 VDD.n413 0.13325
R93009 VDD.n937 VDD.n414 0.13325
R93010 VDD.n936 VDD.n415 0.13325
R93011 VDD.n926 VDD.n426 0.13325
R93012 VDD.n924 VDD.n430 0.13325
R93013 VDD.n947 VDD.n240 0.13325
R93014 VDD.n472 VDD.n471 0.133132
R93015 VDD.n444 VDD.n443 0.133132
R93016 VDD.n752 VDD.n670 0.13175
R93017 VDD.n765 VDD.n670 0.13175
R93018 VDD.n669 VDD.n668 0.13175
R93019 VDD.n765 VDD.n669 0.13175
R93020 VDD.n465 VDD.n462 0.114184
R93021 VDD.n439 VDD.n437 0.114184
R93022 VDD.n287 VDD.n280 0.113
R93023 VDD.n709 VDD.n401 0.110039
R93024 VDD.n695 VDD.n413 0.109447
R93025 VDD.n944 VDD.n408 0.0987895
R93026 VDD.n671 VDD.n436 0.0952368
R93027 VDD.n1130 VDD.n159 0.0905
R93028 VDD.n899 VDD.n488 0.0905
R93029 VDD.n901 VDD.n482 0.0905
R93030 VDD.n903 VDD.n474 0.0905
R93031 VDD.n908 VDD.n460 0.0905
R93032 VDD.n910 VDD.n454 0.0905
R93033 VDD.n912 VDD.n446 0.0905
R93034 VDD.n917 VDD.n436 0.0905
R93035 VDD.n927 VDD.n423 0.0905
R93036 VDD.n710 VDD.n709 0.0905
R93037 VDD.n948 VDD.n946 0.0905
R93038 VDD.n935 VDD.n416 0.0905
R93039 VDD.n925 VDD.n429 0.0905
R93040 VDD.n874 VDD.n873 0.0905
R93041 VDD.n1130 VDD.n160 0.0905
R93042 VDD.n172 VDD.n168 0.0781429
R93043 VDD.n176 VDD.n167 0.0781429
R93044 VDD.n180 VDD.n166 0.0781429
R93045 VDD.n184 VDD.n165 0.0781429
R93046 VDD.n188 VDD.n164 0.0781429
R93047 VDD.n192 VDD.n163 0.0781429
R93048 VDD.n196 VDD.n162 0.0781429
R93049 VDD.n200 VDD.n161 0.0781429
R93050 VDD.n1127 VDD.n168 0.0781429
R93051 VDD.n174 VDD.n167 0.0781429
R93052 VDD.n178 VDD.n166 0.0781429
R93053 VDD.n182 VDD.n165 0.0781429
R93054 VDD.n186 VDD.n164 0.0781429
R93055 VDD.n190 VDD.n163 0.0781429
R93056 VDD.n194 VDD.n162 0.0781429
R93057 VDD.n198 VDD.n161 0.0781429
R93058 VDD.n466 VDD.n465 0.0762895
R93059 VDD.n440 VDD.n439 0.0762895
R93060 VDD.n688 VDD.n416 0.0715526
R93061 VDD.n1067 VDD.n280 0.068
R93062 VDD.n488 VDD.n487 0.0668158
R93063 VDD.n460 VDD.n459 0.0668158
R93064 VDD.n876 VDD.n565 0.0645294
R93065 VDD.n878 VDD.n877 0.061
R93066 VDD.n851 VDD.n589 0.061
R93067 VDD.n1038 VDD.n1037 0.061
R93068 VDD.n499 VDD.n498 0.061
R93069 VDD.n260 VDD.n259 0.061
R93070 VDD.n798 VDD.n797 0.0596957
R93071 VDD.n980 VDD.n382 0.0596957
R93072 VDD.n471 VDD.n468 0.0573421
R93073 VDD.n443 VDD.n441 0.0573421
R93074 VDD.n1070 VDD.n1069 0.0539412
R93075 VDD.n1073 VDD.n1072 0.0539412
R93076 VDD.n768 VDD.n767 0.0526053
R93077 VDD.n711 VDD.n708 0.0526053
R93078 VDD.n693 VDD.n395 0.0526053
R93079 VDD.n717 VDD.n716 0.0526053
R93080 VDD.n691 VDD.n414 0.0526053
R93081 VDD.n723 VDD.n721 0.0526053
R93082 VDD.n730 VDD.n729 0.0526053
R93083 VDD.n404 VDD.n265 0.0526053
R93084 VDD.n1129 VDD.n161 0.0524286
R93085 VDD.n1129 VDD.n162 0.0524286
R93086 VDD.n1129 VDD.n163 0.0524286
R93087 VDD.n1129 VDD.n164 0.0524286
R93088 VDD.n1129 VDD.n165 0.0524286
R93089 VDD.n1129 VDD.n166 0.0524286
R93090 VDD.n1129 VDD.n167 0.0524286
R93091 VDD.n1129 VDD.n168 0.0524286
R93092 VDD.n752 VDD.n751 0.0478684
R93093 VDD.n477 VDD.n474 0.0478684
R93094 VDD.n668 VDD.n462 0.0478684
R93095 VDD.n449 VDD.n446 0.0478684
R93096 VDD.n429 VDD.n428 0.0407632
R93097 VDD.n1678 VDD.n1677 0.0362313
R93098 VDD.n1673 VDD.n0 0.0362313
R93099 VDD.n1674 VDD.n1673 0.0353837
R93100 VDD.n1672 VDD.n1671 0.0353837
R93101 VDD.n1415 VDD.n3 0.0353837
R93102 VDD.n1544 VDD.n4 0.0353837
R93103 VDD.n1414 VDD.n5 0.0353837
R93104 VDD.n1261 VDD.n1260 0.0353837
R93105 VDD.n1413 VDD.n8 0.0353837
R93106 VDD.n1262 VDD.n9 0.0353837
R93107 VDD.n1412 VDD.n10 0.0353837
R93108 VDD.n1264 VDD.n1263 0.0353837
R93109 VDD.n1411 VDD.n13 0.0353837
R93110 VDD.n1265 VDD.n14 0.0353837
R93111 VDD.n1410 VDD.n15 0.0353837
R93112 VDD.n1267 VDD.n1266 0.0353837
R93113 VDD.n1409 VDD.n18 0.0353837
R93114 VDD.n1268 VDD.n19 0.0353837
R93115 VDD.n1408 VDD.n20 0.0353837
R93116 VDD.n1270 VDD.n1269 0.0353837
R93117 VDD.n1407 VDD.n23 0.0353837
R93118 VDD.n1271 VDD.n24 0.0353837
R93119 VDD.n1406 VDD.n25 0.0353837
R93120 VDD.n1273 VDD.n1272 0.0353837
R93121 VDD.n1405 VDD.n28 0.0353837
R93122 VDD.n1274 VDD.n29 0.0353837
R93123 VDD.n1404 VDD.n30 0.0353837
R93124 VDD.n1276 VDD.n1275 0.0353837
R93125 VDD.n1403 VDD.n33 0.0353837
R93126 VDD.n1277 VDD.n34 0.0353837
R93127 VDD.n1402 VDD.n35 0.0353837
R93128 VDD.n1279 VDD.n1278 0.0353837
R93129 VDD.n1401 VDD.n38 0.0353837
R93130 VDD.n1280 VDD.n39 0.0353837
R93131 VDD.n1400 VDD.n40 0.0353837
R93132 VDD.n1282 VDD.n1281 0.0353837
R93133 VDD.n1399 VDD.n43 0.0353837
R93134 VDD.n1283 VDD.n44 0.0353837
R93135 VDD.n1398 VDD.n45 0.0353837
R93136 VDD.n1285 VDD.n1284 0.0353837
R93137 VDD.n1397 VDD.n48 0.0353837
R93138 VDD.n1286 VDD.n49 0.0353837
R93139 VDD.n1396 VDD.n50 0.0353837
R93140 VDD.n1288 VDD.n1287 0.0353837
R93141 VDD.n1395 VDD.n53 0.0353837
R93142 VDD.n1289 VDD.n54 0.0353837
R93143 VDD.n1394 VDD.n55 0.0353837
R93144 VDD.n1291 VDD.n1290 0.0353837
R93145 VDD.n1393 VDD.n58 0.0353837
R93146 VDD.n1292 VDD.n59 0.0353837
R93147 VDD.n1392 VDD.n60 0.0353837
R93148 VDD.n1294 VDD.n1293 0.0353837
R93149 VDD.n1391 VDD.n63 0.0353837
R93150 VDD.n1295 VDD.n64 0.0353837
R93151 VDD.n1390 VDD.n65 0.0353837
R93152 VDD.n1297 VDD.n1296 0.0353837
R93153 VDD.n1389 VDD.n68 0.0353837
R93154 VDD.n1298 VDD.n69 0.0353837
R93155 VDD.n1388 VDD.n70 0.0353837
R93156 VDD.n1300 VDD.n1299 0.0353837
R93157 VDD.n1387 VDD.n73 0.0353837
R93158 VDD.n1301 VDD.n74 0.0353837
R93159 VDD.n1386 VDD.n75 0.0353837
R93160 VDD.n1303 VDD.n1302 0.0353837
R93161 VDD.n1385 VDD.n78 0.0353837
R93162 VDD.n1304 VDD.n79 0.0353837
R93163 VDD.n1384 VDD.n80 0.0353837
R93164 VDD.n1306 VDD.n1305 0.0353837
R93165 VDD.n1383 VDD.n83 0.0353837
R93166 VDD.n1307 VDD.n84 0.0353837
R93167 VDD.n1382 VDD.n85 0.0353837
R93168 VDD.n1309 VDD.n1308 0.0353837
R93169 VDD.n1381 VDD.n88 0.0353837
R93170 VDD.n1310 VDD.n89 0.0353837
R93171 VDD.n1380 VDD.n90 0.0353837
R93172 VDD.n1312 VDD.n1311 0.0353837
R93173 VDD.n1379 VDD.n93 0.0353837
R93174 VDD.n1313 VDD.n94 0.0353837
R93175 VDD.n1378 VDD.n95 0.0353837
R93176 VDD.n1315 VDD.n1314 0.0353837
R93177 VDD.n1377 VDD.n98 0.0353837
R93178 VDD.n1316 VDD.n99 0.0353837
R93179 VDD.n1376 VDD.n100 0.0353837
R93180 VDD.n1318 VDD.n1317 0.0353837
R93181 VDD.n1375 VDD.n102 0.0353837
R93182 VDD.n1319 VDD.n103 0.0353837
R93183 VDD.n1374 VDD.n1373 0.0353837
R93184 VDD.n1320 VDD.n106 0.0353837
R93185 VDD.n1372 VDD.n107 0.0353837
R93186 VDD.n1321 VDD.n108 0.0353837
R93187 VDD.n1371 VDD.n1370 0.0353837
R93188 VDD.n1322 VDD.n111 0.0353837
R93189 VDD.n1369 VDD.n112 0.0353837
R93190 VDD.n1323 VDD.n113 0.0353837
R93191 VDD.n1368 VDD.n1367 0.0353837
R93192 VDD.n1324 VDD.n116 0.0353837
R93193 VDD.n1366 VDD.n117 0.0353837
R93194 VDD.n1325 VDD.n118 0.0353837
R93195 VDD.n1365 VDD.n1364 0.0353837
R93196 VDD.n1326 VDD.n121 0.0353837
R93197 VDD.n1363 VDD.n122 0.0353837
R93198 VDD.n1327 VDD.n123 0.0353837
R93199 VDD.n1362 VDD.n1361 0.0353837
R93200 VDD.n1328 VDD.n126 0.0353837
R93201 VDD.n1360 VDD.n127 0.0353837
R93202 VDD.n1329 VDD.n128 0.0353837
R93203 VDD.n1359 VDD.n1358 0.0353837
R93204 VDD.n1330 VDD.n131 0.0353837
R93205 VDD.n1357 VDD.n132 0.0353837
R93206 VDD.n1331 VDD.n133 0.0353837
R93207 VDD.n1356 VDD.n1355 0.0353837
R93208 VDD.n1332 VDD.n136 0.0353837
R93209 VDD.n1354 VDD.n137 0.0353837
R93210 VDD.n1333 VDD.n138 0.0353837
R93211 VDD.n1353 VDD.n1352 0.0353837
R93212 VDD.n1334 VDD.n141 0.0353837
R93213 VDD.n1351 VDD.n142 0.0353837
R93214 VDD.n1335 VDD.n143 0.0353837
R93215 VDD.n1350 VDD.n1349 0.0353837
R93216 VDD.n1336 VDD.n146 0.0353837
R93217 VDD.n1348 VDD.n147 0.0353837
R93218 VDD.n1337 VDD.n148 0.0353837
R93219 VDD.n1347 VDD.n1346 0.0353837
R93220 VDD.n1338 VDD.n151 0.0353837
R93221 VDD.n1345 VDD.n152 0.0353837
R93222 VDD.n1339 VDD.n153 0.0353837
R93223 VDD.n1344 VDD.n1343 0.0353837
R93224 VDD.n1340 VDD.n156 0.0353837
R93225 VDD.n1342 VDD.n157 0.0353837
R93226 VDD.n1341 VDD.n158 0.0353837
R93227 VDD.n1677 VDD.n1676 0.0353837
R93228 VDD.n1672 VDD.n2 0.0353837
R93229 VDD.n1866 VDD.n3 0.0353837
R93230 VDD.n1865 VDD.n4 0.0353837
R93231 VDD.n1864 VDD.n5 0.0353837
R93232 VDD.n1260 VDD.n6 0.0353837
R93233 VDD.n1860 VDD.n8 0.0353837
R93234 VDD.n1859 VDD.n9 0.0353837
R93235 VDD.n1858 VDD.n10 0.0353837
R93236 VDD.n1263 VDD.n11 0.0353837
R93237 VDD.n1854 VDD.n13 0.0353837
R93238 VDD.n1853 VDD.n14 0.0353837
R93239 VDD.n1852 VDD.n15 0.0353837
R93240 VDD.n1266 VDD.n16 0.0353837
R93241 VDD.n1848 VDD.n18 0.0353837
R93242 VDD.n1847 VDD.n19 0.0353837
R93243 VDD.n1846 VDD.n20 0.0353837
R93244 VDD.n1269 VDD.n21 0.0353837
R93245 VDD.n1842 VDD.n23 0.0353837
R93246 VDD.n1841 VDD.n24 0.0353837
R93247 VDD.n1840 VDD.n25 0.0353837
R93248 VDD.n1272 VDD.n26 0.0353837
R93249 VDD.n1836 VDD.n28 0.0353837
R93250 VDD.n1835 VDD.n29 0.0353837
R93251 VDD.n1834 VDD.n30 0.0353837
R93252 VDD.n1275 VDD.n31 0.0353837
R93253 VDD.n1830 VDD.n33 0.0353837
R93254 VDD.n1829 VDD.n34 0.0353837
R93255 VDD.n1828 VDD.n35 0.0353837
R93256 VDD.n1278 VDD.n36 0.0353837
R93257 VDD.n1824 VDD.n38 0.0353837
R93258 VDD.n1823 VDD.n39 0.0353837
R93259 VDD.n1822 VDD.n40 0.0353837
R93260 VDD.n1281 VDD.n41 0.0353837
R93261 VDD.n1818 VDD.n43 0.0353837
R93262 VDD.n1817 VDD.n44 0.0353837
R93263 VDD.n1816 VDD.n45 0.0353837
R93264 VDD.n1284 VDD.n46 0.0353837
R93265 VDD.n1812 VDD.n48 0.0353837
R93266 VDD.n1811 VDD.n49 0.0353837
R93267 VDD.n1810 VDD.n50 0.0353837
R93268 VDD.n1287 VDD.n51 0.0353837
R93269 VDD.n1806 VDD.n53 0.0353837
R93270 VDD.n1805 VDD.n54 0.0353837
R93271 VDD.n1804 VDD.n55 0.0353837
R93272 VDD.n1290 VDD.n56 0.0353837
R93273 VDD.n1800 VDD.n58 0.0353837
R93274 VDD.n1799 VDD.n59 0.0353837
R93275 VDD.n1798 VDD.n60 0.0353837
R93276 VDD.n1293 VDD.n61 0.0353837
R93277 VDD.n1794 VDD.n63 0.0353837
R93278 VDD.n1793 VDD.n64 0.0353837
R93279 VDD.n1792 VDD.n65 0.0353837
R93280 VDD.n1296 VDD.n66 0.0353837
R93281 VDD.n1788 VDD.n68 0.0353837
R93282 VDD.n1787 VDD.n69 0.0353837
R93283 VDD.n1786 VDD.n70 0.0353837
R93284 VDD.n1299 VDD.n71 0.0353837
R93285 VDD.n1782 VDD.n73 0.0353837
R93286 VDD.n1781 VDD.n74 0.0353837
R93287 VDD.n1780 VDD.n75 0.0353837
R93288 VDD.n1302 VDD.n76 0.0353837
R93289 VDD.n1776 VDD.n78 0.0353837
R93290 VDD.n1775 VDD.n79 0.0353837
R93291 VDD.n1774 VDD.n80 0.0353837
R93292 VDD.n1305 VDD.n81 0.0353837
R93293 VDD.n1770 VDD.n83 0.0353837
R93294 VDD.n1769 VDD.n84 0.0353837
R93295 VDD.n1768 VDD.n85 0.0353837
R93296 VDD.n1308 VDD.n86 0.0353837
R93297 VDD.n1764 VDD.n88 0.0353837
R93298 VDD.n1763 VDD.n89 0.0353837
R93299 VDD.n1762 VDD.n90 0.0353837
R93300 VDD.n1311 VDD.n91 0.0353837
R93301 VDD.n1758 VDD.n93 0.0353837
R93302 VDD.n1757 VDD.n94 0.0353837
R93303 VDD.n1756 VDD.n95 0.0353837
R93304 VDD.n1314 VDD.n96 0.0353837
R93305 VDD.n1752 VDD.n98 0.0353837
R93306 VDD.n1751 VDD.n99 0.0353837
R93307 VDD.n1750 VDD.n100 0.0353837
R93308 VDD.n1317 VDD.n101 0.0353837
R93309 VDD.n1746 VDD.n102 0.0353837
R93310 VDD.n1745 VDD.n103 0.0353837
R93311 VDD.n1373 VDD.n104 0.0353837
R93312 VDD.n1741 VDD.n106 0.0353837
R93313 VDD.n1740 VDD.n107 0.0353837
R93314 VDD.n1739 VDD.n108 0.0353837
R93315 VDD.n1370 VDD.n109 0.0353837
R93316 VDD.n1735 VDD.n111 0.0353837
R93317 VDD.n1734 VDD.n112 0.0353837
R93318 VDD.n1733 VDD.n113 0.0353837
R93319 VDD.n1367 VDD.n114 0.0353837
R93320 VDD.n1729 VDD.n116 0.0353837
R93321 VDD.n1728 VDD.n117 0.0353837
R93322 VDD.n1727 VDD.n118 0.0353837
R93323 VDD.n1364 VDD.n119 0.0353837
R93324 VDD.n1723 VDD.n121 0.0353837
R93325 VDD.n1722 VDD.n122 0.0353837
R93326 VDD.n1721 VDD.n123 0.0353837
R93327 VDD.n1361 VDD.n124 0.0353837
R93328 VDD.n1717 VDD.n126 0.0353837
R93329 VDD.n1716 VDD.n127 0.0353837
R93330 VDD.n1715 VDD.n128 0.0353837
R93331 VDD.n1358 VDD.n129 0.0353837
R93332 VDD.n1711 VDD.n131 0.0353837
R93333 VDD.n1710 VDD.n132 0.0353837
R93334 VDD.n1709 VDD.n133 0.0353837
R93335 VDD.n1355 VDD.n134 0.0353837
R93336 VDD.n1705 VDD.n136 0.0353837
R93337 VDD.n1704 VDD.n137 0.0353837
R93338 VDD.n1703 VDD.n138 0.0353837
R93339 VDD.n1352 VDD.n139 0.0353837
R93340 VDD.n1699 VDD.n141 0.0353837
R93341 VDD.n1698 VDD.n142 0.0353837
R93342 VDD.n1697 VDD.n143 0.0353837
R93343 VDD.n1349 VDD.n144 0.0353837
R93344 VDD.n1693 VDD.n146 0.0353837
R93345 VDD.n1692 VDD.n147 0.0353837
R93346 VDD.n1691 VDD.n148 0.0353837
R93347 VDD.n1346 VDD.n149 0.0353837
R93348 VDD.n1687 VDD.n151 0.0353837
R93349 VDD.n1686 VDD.n152 0.0353837
R93350 VDD.n1685 VDD.n153 0.0353837
R93351 VDD.n1343 VDD.n154 0.0353837
R93352 VDD.n1681 VDD.n156 0.0353837
R93353 VDD.n1680 VDD.n157 0.0353837
R93354 VDD.n1679 VDD.n158 0.0353837
R93355 VDD.n1867 VDD.n1866 0.0353837
R93356 VDD.n1865 VDD.n1 0.0353837
R93357 VDD.n1864 VDD.n1863 0.0353837
R93358 VDD.n1862 VDD.n6 0.0353837
R93359 VDD.n1861 VDD.n1860 0.0353837
R93360 VDD.n1859 VDD.n7 0.0353837
R93361 VDD.n1858 VDD.n1857 0.0353837
R93362 VDD.n1856 VDD.n11 0.0353837
R93363 VDD.n1855 VDD.n1854 0.0353837
R93364 VDD.n1853 VDD.n12 0.0353837
R93365 VDD.n1852 VDD.n1851 0.0353837
R93366 VDD.n1850 VDD.n16 0.0353837
R93367 VDD.n1849 VDD.n1848 0.0353837
R93368 VDD.n1847 VDD.n17 0.0353837
R93369 VDD.n1846 VDD.n1845 0.0353837
R93370 VDD.n1844 VDD.n21 0.0353837
R93371 VDD.n1843 VDD.n1842 0.0353837
R93372 VDD.n1841 VDD.n22 0.0353837
R93373 VDD.n1840 VDD.n1839 0.0353837
R93374 VDD.n1838 VDD.n26 0.0353837
R93375 VDD.n1837 VDD.n1836 0.0353837
R93376 VDD.n1835 VDD.n27 0.0353837
R93377 VDD.n1834 VDD.n1833 0.0353837
R93378 VDD.n1832 VDD.n31 0.0353837
R93379 VDD.n1831 VDD.n1830 0.0353837
R93380 VDD.n1829 VDD.n32 0.0353837
R93381 VDD.n1828 VDD.n1827 0.0353837
R93382 VDD.n1826 VDD.n36 0.0353837
R93383 VDD.n1825 VDD.n1824 0.0353837
R93384 VDD.n1823 VDD.n37 0.0353837
R93385 VDD.n1822 VDD.n1821 0.0353837
R93386 VDD.n1820 VDD.n41 0.0353837
R93387 VDD.n1819 VDD.n1818 0.0353837
R93388 VDD.n1817 VDD.n42 0.0353837
R93389 VDD.n1816 VDD.n1815 0.0353837
R93390 VDD.n1814 VDD.n46 0.0353837
R93391 VDD.n1813 VDD.n1812 0.0353837
R93392 VDD.n1811 VDD.n47 0.0353837
R93393 VDD.n1810 VDD.n1809 0.0353837
R93394 VDD.n1808 VDD.n51 0.0353837
R93395 VDD.n1807 VDD.n1806 0.0353837
R93396 VDD.n1805 VDD.n52 0.0353837
R93397 VDD.n1804 VDD.n1803 0.0353837
R93398 VDD.n1802 VDD.n56 0.0353837
R93399 VDD.n1801 VDD.n1800 0.0353837
R93400 VDD.n1799 VDD.n57 0.0353837
R93401 VDD.n1798 VDD.n1797 0.0353837
R93402 VDD.n1796 VDD.n61 0.0353837
R93403 VDD.n1795 VDD.n1794 0.0353837
R93404 VDD.n1793 VDD.n62 0.0353837
R93405 VDD.n1792 VDD.n1791 0.0353837
R93406 VDD.n1790 VDD.n66 0.0353837
R93407 VDD.n1789 VDD.n1788 0.0353837
R93408 VDD.n1787 VDD.n67 0.0353837
R93409 VDD.n1786 VDD.n1785 0.0353837
R93410 VDD.n1784 VDD.n71 0.0353837
R93411 VDD.n1783 VDD.n1782 0.0353837
R93412 VDD.n1781 VDD.n72 0.0353837
R93413 VDD.n1780 VDD.n1779 0.0353837
R93414 VDD.n1778 VDD.n76 0.0353837
R93415 VDD.n1777 VDD.n1776 0.0353837
R93416 VDD.n1775 VDD.n77 0.0353837
R93417 VDD.n1774 VDD.n1773 0.0353837
R93418 VDD.n1772 VDD.n81 0.0353837
R93419 VDD.n1771 VDD.n1770 0.0353837
R93420 VDD.n1769 VDD.n82 0.0353837
R93421 VDD.n1768 VDD.n1767 0.0353837
R93422 VDD.n1766 VDD.n86 0.0353837
R93423 VDD.n1765 VDD.n1764 0.0353837
R93424 VDD.n1763 VDD.n87 0.0353837
R93425 VDD.n1762 VDD.n1761 0.0353837
R93426 VDD.n1760 VDD.n91 0.0353837
R93427 VDD.n1759 VDD.n1758 0.0353837
R93428 VDD.n1757 VDD.n92 0.0353837
R93429 VDD.n1756 VDD.n1755 0.0353837
R93430 VDD.n1754 VDD.n96 0.0353837
R93431 VDD.n1753 VDD.n1752 0.0353837
R93432 VDD.n1751 VDD.n97 0.0353837
R93433 VDD.n1750 VDD.n1749 0.0353837
R93434 VDD.n1748 VDD.n101 0.0353837
R93435 VDD.n1747 VDD.n1746 0.0353837
R93436 VDD.n1745 VDD.n1744 0.0353837
R93437 VDD.n1743 VDD.n104 0.0353837
R93438 VDD.n1742 VDD.n1741 0.0353837
R93439 VDD.n1740 VDD.n105 0.0353837
R93440 VDD.n1739 VDD.n1738 0.0353837
R93441 VDD.n1737 VDD.n109 0.0353837
R93442 VDD.n1736 VDD.n1735 0.0353837
R93443 VDD.n1734 VDD.n110 0.0353837
R93444 VDD.n1733 VDD.n1732 0.0353837
R93445 VDD.n1731 VDD.n114 0.0353837
R93446 VDD.n1730 VDD.n1729 0.0353837
R93447 VDD.n1728 VDD.n115 0.0353837
R93448 VDD.n1727 VDD.n1726 0.0353837
R93449 VDD.n1725 VDD.n119 0.0353837
R93450 VDD.n1724 VDD.n1723 0.0353837
R93451 VDD.n1722 VDD.n120 0.0353837
R93452 VDD.n1721 VDD.n1720 0.0353837
R93453 VDD.n1719 VDD.n124 0.0353837
R93454 VDD.n1718 VDD.n1717 0.0353837
R93455 VDD.n1716 VDD.n125 0.0353837
R93456 VDD.n1715 VDD.n1714 0.0353837
R93457 VDD.n1713 VDD.n129 0.0353837
R93458 VDD.n1712 VDD.n1711 0.0353837
R93459 VDD.n1710 VDD.n130 0.0353837
R93460 VDD.n1709 VDD.n1708 0.0353837
R93461 VDD.n1707 VDD.n134 0.0353837
R93462 VDD.n1706 VDD.n1705 0.0353837
R93463 VDD.n1704 VDD.n135 0.0353837
R93464 VDD.n1703 VDD.n1702 0.0353837
R93465 VDD.n1701 VDD.n139 0.0353837
R93466 VDD.n1700 VDD.n1699 0.0353837
R93467 VDD.n1698 VDD.n140 0.0353837
R93468 VDD.n1697 VDD.n1696 0.0353837
R93469 VDD.n1695 VDD.n144 0.0353837
R93470 VDD.n1694 VDD.n1693 0.0353837
R93471 VDD.n1692 VDD.n145 0.0353837
R93472 VDD.n1691 VDD.n1690 0.0353837
R93473 VDD.n1689 VDD.n149 0.0353837
R93474 VDD.n1688 VDD.n1687 0.0353837
R93475 VDD.n1686 VDD.n150 0.0353837
R93476 VDD.n1685 VDD.n1684 0.0353837
R93477 VDD.n1683 VDD.n154 0.0353837
R93478 VDD.n1682 VDD.n1681 0.0353837
R93479 VDD.n1680 VDD.n155 0.0353837
R93480 VDD.n285 VDD.n280 0.023
R93481 VDD.n1867 VDD.n0 0.0188497
R93482 VDD.n1678 VDD.n155 0.0188497
R93483 VDD.n425 VDD.n423 0.0158947
R93484 VDD.n949 VDD.n948 0.0147105
R93485 VDD.n482 VDD.n481 0.00997368
R93486 VDD.n454 VDD.n453 0.00997368
R93487 VDD.n706 VDD.n408 0.00523684
R93488 VDD.n1130 VDD.n1129 0.0023
R93489 VDD.n1480 VDD.n1195 0.00134872
R93490 VDD.n1670 VDD.n1416 0.00134872
R93491 VDD.n1482 VDD.n1196 0.00134872
R93492 VDD.n1669 VDD.n1193 0.00134872
R93493 VDD.n1483 VDD.n1197 0.00134872
R93494 VDD.n1668 VDD.n1192 0.00134872
R93495 VDD.n1484 VDD.n1198 0.00134872
R93496 VDD.n1667 VDD.n1191 0.00134872
R93497 VDD.n1485 VDD.n1199 0.00134872
R93498 VDD.n1666 VDD.n1190 0.00134872
R93499 VDD.n1486 VDD.n1200 0.00134872
R93500 VDD.n1665 VDD.n1189 0.00134872
R93501 VDD.n1487 VDD.n1201 0.00134872
R93502 VDD.n1664 VDD.n1188 0.00134872
R93503 VDD.n1488 VDD.n1202 0.00134872
R93504 VDD.n1663 VDD.n1187 0.00134872
R93505 VDD.n1489 VDD.n1203 0.00134872
R93506 VDD.n1662 VDD.n1186 0.00134872
R93507 VDD.n1490 VDD.n1204 0.00134872
R93508 VDD.n1661 VDD.n1185 0.00134872
R93509 VDD.n1491 VDD.n1205 0.00134872
R93510 VDD.n1660 VDD.n1184 0.00134872
R93511 VDD.n1492 VDD.n1206 0.00134872
R93512 VDD.n1659 VDD.n1183 0.00134872
R93513 VDD.n1493 VDD.n1207 0.00134872
R93514 VDD.n1658 VDD.n1182 0.00134872
R93515 VDD.n1494 VDD.n1208 0.00134872
R93516 VDD.n1657 VDD.n1181 0.00134872
R93517 VDD.n1495 VDD.n1209 0.00134872
R93518 VDD.n1656 VDD.n1180 0.00134872
R93519 VDD.n1496 VDD.n1210 0.00134872
R93520 VDD.n1655 VDD.n1179 0.00134872
R93521 VDD.n1497 VDD.n1211 0.00134872
R93522 VDD.n1654 VDD.n1178 0.00134872
R93523 VDD.n1498 VDD.n1212 0.00134872
R93524 VDD.n1653 VDD.n1177 0.00134872
R93525 VDD.n1499 VDD.n1213 0.00134872
R93526 VDD.n1652 VDD.n1176 0.00134872
R93527 VDD.n1500 VDD.n1214 0.00134872
R93528 VDD.n1651 VDD.n1175 0.00134872
R93529 VDD.n1501 VDD.n1215 0.00134872
R93530 VDD.n1650 VDD.n1174 0.00134872
R93531 VDD.n1502 VDD.n1216 0.00134872
R93532 VDD.n1649 VDD.n1173 0.00134872
R93533 VDD.n1503 VDD.n1217 0.00134872
R93534 VDD.n1648 VDD.n1172 0.00134872
R93535 VDD.n1504 VDD.n1218 0.00134872
R93536 VDD.n1647 VDD.n1171 0.00134872
R93537 VDD.n1505 VDD.n1219 0.00134872
R93538 VDD.n1646 VDD.n1170 0.00134872
R93539 VDD.n1506 VDD.n1220 0.00134872
R93540 VDD.n1645 VDD.n1169 0.00134872
R93541 VDD.n1507 VDD.n1221 0.00134872
R93542 VDD.n1644 VDD.n1168 0.00134872
R93543 VDD.n1508 VDD.n1222 0.00134872
R93544 VDD.n1643 VDD.n1167 0.00134872
R93545 VDD.n1509 VDD.n1223 0.00134872
R93546 VDD.n1642 VDD.n1166 0.00134872
R93547 VDD.n1510 VDD.n1224 0.00134872
R93548 VDD.n1641 VDD.n1165 0.00134872
R93549 VDD.n1511 VDD.n1225 0.00134872
R93550 VDD.n1640 VDD.n1164 0.00134872
R93551 VDD.n1512 VDD.n1226 0.00134872
R93552 VDD.n1639 VDD.n1163 0.00134872
R93553 VDD.n1513 VDD.n1227 0.00134872
R93554 VDD.n1638 VDD.n1162 0.00134872
R93555 VDD.n1514 VDD.n1228 0.00134872
R93556 VDD.n1637 VDD.n1161 0.00134872
R93557 VDD.n1515 VDD.n1229 0.00134872
R93558 VDD.n1636 VDD.n1160 0.00134872
R93559 VDD.n1516 VDD.n1230 0.00134872
R93560 VDD.n1635 VDD.n1159 0.00134872
R93561 VDD.n1517 VDD.n1231 0.00134872
R93562 VDD.n1634 VDD.n1158 0.00134872
R93563 VDD.n1518 VDD.n1232 0.00134872
R93564 VDD.n1633 VDD.n1157 0.00134872
R93565 VDD.n1519 VDD.n1233 0.00134872
R93566 VDD.n1632 VDD.n1156 0.00134872
R93567 VDD.n1520 VDD.n1234 0.00134872
R93568 VDD.n1631 VDD.n1155 0.00134872
R93569 VDD.n1521 VDD.n1235 0.00134872
R93570 VDD.n1630 VDD.n1154 0.00134872
R93571 VDD.n1522 VDD.n1236 0.00134872
R93572 VDD.n1629 VDD.n1153 0.00134872
R93573 VDD.n1523 VDD.n1237 0.00134872
R93574 VDD.n1628 VDD.n1152 0.00134872
R93575 VDD.n1524 VDD.n1238 0.00134872
R93576 VDD.n1627 VDD.n1151 0.00134872
R93577 VDD.n1525 VDD.n1239 0.00134872
R93578 VDD.n1626 VDD.n1150 0.00134872
R93579 VDD.n1526 VDD.n1240 0.00134872
R93580 VDD.n1625 VDD.n1149 0.00134872
R93581 VDD.n1527 VDD.n1241 0.00134872
R93582 VDD.n1624 VDD.n1148 0.00134872
R93583 VDD.n1528 VDD.n1242 0.00134872
R93584 VDD.n1623 VDD.n1147 0.00134872
R93585 VDD.n1529 VDD.n1243 0.00134872
R93586 VDD.n1622 VDD.n1146 0.00134872
R93587 VDD.n1530 VDD.n1244 0.00134872
R93588 VDD.n1621 VDD.n1145 0.00134872
R93589 VDD.n1531 VDD.n1245 0.00134872
R93590 VDD.n1620 VDD.n1144 0.00134872
R93591 VDD.n1532 VDD.n1246 0.00134872
R93592 VDD.n1619 VDD.n1143 0.00134872
R93593 VDD.n1533 VDD.n1247 0.00134872
R93594 VDD.n1618 VDD.n1142 0.00134872
R93595 VDD.n1534 VDD.n1248 0.00134872
R93596 VDD.n1617 VDD.n1141 0.00134872
R93597 VDD.n1535 VDD.n1249 0.00134872
R93598 VDD.n1616 VDD.n1140 0.00134872
R93599 VDD.n1536 VDD.n1250 0.00134872
R93600 VDD.n1615 VDD.n1139 0.00134872
R93601 VDD.n1537 VDD.n1251 0.00134872
R93602 VDD.n1614 VDD.n1138 0.00134872
R93603 VDD.n1538 VDD.n1252 0.00134872
R93604 VDD.n1613 VDD.n1137 0.00134872
R93605 VDD.n1539 VDD.n1253 0.00134872
R93606 VDD.n1612 VDD.n1136 0.00134872
R93607 VDD.n1540 VDD.n1254 0.00134872
R93608 VDD.n1611 VDD.n1135 0.00134872
R93609 VDD.n1541 VDD.n1255 0.00134872
R93610 VDD.n1610 VDD.n1134 0.00134872
R93611 VDD.n1542 VDD.n1256 0.00134872
R93612 VDD.n1609 VDD.n1133 0.00134872
R93613 VDD.n1543 VDD.n1257 0.00134872
R93614 VDD.n1608 VDD.n1132 0.00134872
R93615 VDD.n1675 VDD.n1258 0.00134872
R93616 VDD.n1259 VDD.n1131 0.00134872
R93617 VDD.n1674 VDD.n1417 0.00134872
R93618 VDD.n1481 VDD.n1415 0.00134872
R93619 VDD.n1545 VDD.n1544 0.00134872
R93620 VDD.n1418 VDD.n1414 0.00134872
R93621 VDD.n1546 VDD.n1261 0.00134872
R93622 VDD.n1419 VDD.n1413 0.00134872
R93623 VDD.n1547 VDD.n1262 0.00134872
R93624 VDD.n1420 VDD.n1412 0.00134872
R93625 VDD.n1548 VDD.n1264 0.00134872
R93626 VDD.n1421 VDD.n1411 0.00134872
R93627 VDD.n1549 VDD.n1265 0.00134872
R93628 VDD.n1422 VDD.n1410 0.00134872
R93629 VDD.n1550 VDD.n1267 0.00134872
R93630 VDD.n1423 VDD.n1409 0.00134872
R93631 VDD.n1551 VDD.n1268 0.00134872
R93632 VDD.n1424 VDD.n1408 0.00134872
R93633 VDD.n1552 VDD.n1270 0.00134872
R93634 VDD.n1425 VDD.n1407 0.00134872
R93635 VDD.n1553 VDD.n1271 0.00134872
R93636 VDD.n1426 VDD.n1406 0.00134872
R93637 VDD.n1554 VDD.n1273 0.00134872
R93638 VDD.n1427 VDD.n1405 0.00134872
R93639 VDD.n1555 VDD.n1274 0.00134872
R93640 VDD.n1428 VDD.n1404 0.00134872
R93641 VDD.n1556 VDD.n1276 0.00134872
R93642 VDD.n1429 VDD.n1403 0.00134872
R93643 VDD.n1557 VDD.n1277 0.00134872
R93644 VDD.n1430 VDD.n1402 0.00134872
R93645 VDD.n1558 VDD.n1279 0.00134872
R93646 VDD.n1431 VDD.n1401 0.00134872
R93647 VDD.n1559 VDD.n1280 0.00134872
R93648 VDD.n1432 VDD.n1400 0.00134872
R93649 VDD.n1560 VDD.n1282 0.00134872
R93650 VDD.n1433 VDD.n1399 0.00134872
R93651 VDD.n1561 VDD.n1283 0.00134872
R93652 VDD.n1434 VDD.n1398 0.00134872
R93653 VDD.n1562 VDD.n1285 0.00134872
R93654 VDD.n1435 VDD.n1397 0.00134872
R93655 VDD.n1563 VDD.n1286 0.00134872
R93656 VDD.n1436 VDD.n1396 0.00134872
R93657 VDD.n1564 VDD.n1288 0.00134872
R93658 VDD.n1437 VDD.n1395 0.00134872
R93659 VDD.n1565 VDD.n1289 0.00134872
R93660 VDD.n1438 VDD.n1394 0.00134872
R93661 VDD.n1566 VDD.n1291 0.00134872
R93662 VDD.n1439 VDD.n1393 0.00134872
R93663 VDD.n1567 VDD.n1292 0.00134872
R93664 VDD.n1440 VDD.n1392 0.00134872
R93665 VDD.n1568 VDD.n1294 0.00134872
R93666 VDD.n1441 VDD.n1391 0.00134872
R93667 VDD.n1569 VDD.n1295 0.00134872
R93668 VDD.n1442 VDD.n1390 0.00134872
R93669 VDD.n1570 VDD.n1297 0.00134872
R93670 VDD.n1443 VDD.n1389 0.00134872
R93671 VDD.n1571 VDD.n1298 0.00134872
R93672 VDD.n1444 VDD.n1388 0.00134872
R93673 VDD.n1572 VDD.n1300 0.00134872
R93674 VDD.n1445 VDD.n1387 0.00134872
R93675 VDD.n1573 VDD.n1301 0.00134872
R93676 VDD.n1446 VDD.n1386 0.00134872
R93677 VDD.n1574 VDD.n1303 0.00134872
R93678 VDD.n1447 VDD.n1385 0.00134872
R93679 VDD.n1575 VDD.n1304 0.00134872
R93680 VDD.n1448 VDD.n1384 0.00134872
R93681 VDD.n1576 VDD.n1306 0.00134872
R93682 VDD.n1449 VDD.n1383 0.00134872
R93683 VDD.n1577 VDD.n1307 0.00134872
R93684 VDD.n1450 VDD.n1382 0.00134872
R93685 VDD.n1578 VDD.n1309 0.00134872
R93686 VDD.n1451 VDD.n1381 0.00134872
R93687 VDD.n1579 VDD.n1310 0.00134872
R93688 VDD.n1452 VDD.n1380 0.00134872
R93689 VDD.n1580 VDD.n1312 0.00134872
R93690 VDD.n1453 VDD.n1379 0.00134872
R93691 VDD.n1581 VDD.n1313 0.00134872
R93692 VDD.n1454 VDD.n1378 0.00134872
R93693 VDD.n1582 VDD.n1315 0.00134872
R93694 VDD.n1455 VDD.n1377 0.00134872
R93695 VDD.n1583 VDD.n1316 0.00134872
R93696 VDD.n1456 VDD.n1376 0.00134872
R93697 VDD.n1584 VDD.n1318 0.00134872
R93698 VDD.n1457 VDD.n1375 0.00134872
R93699 VDD.n1585 VDD.n1319 0.00134872
R93700 VDD.n1458 VDD.n1374 0.00134872
R93701 VDD.n1586 VDD.n1320 0.00134872
R93702 VDD.n1459 VDD.n1372 0.00134872
R93703 VDD.n1587 VDD.n1321 0.00134872
R93704 VDD.n1460 VDD.n1371 0.00134872
R93705 VDD.n1588 VDD.n1322 0.00134872
R93706 VDD.n1461 VDD.n1369 0.00134872
R93707 VDD.n1589 VDD.n1323 0.00134872
R93708 VDD.n1462 VDD.n1368 0.00134872
R93709 VDD.n1590 VDD.n1324 0.00134872
R93710 VDD.n1463 VDD.n1366 0.00134872
R93711 VDD.n1591 VDD.n1325 0.00134872
R93712 VDD.n1464 VDD.n1365 0.00134872
R93713 VDD.n1592 VDD.n1326 0.00134872
R93714 VDD.n1465 VDD.n1363 0.00134872
R93715 VDD.n1593 VDD.n1327 0.00134872
R93716 VDD.n1466 VDD.n1362 0.00134872
R93717 VDD.n1594 VDD.n1328 0.00134872
R93718 VDD.n1467 VDD.n1360 0.00134872
R93719 VDD.n1595 VDD.n1329 0.00134872
R93720 VDD.n1468 VDD.n1359 0.00134872
R93721 VDD.n1596 VDD.n1330 0.00134872
R93722 VDD.n1469 VDD.n1357 0.00134872
R93723 VDD.n1597 VDD.n1331 0.00134872
R93724 VDD.n1470 VDD.n1356 0.00134872
R93725 VDD.n1598 VDD.n1332 0.00134872
R93726 VDD.n1471 VDD.n1354 0.00134872
R93727 VDD.n1599 VDD.n1333 0.00134872
R93728 VDD.n1472 VDD.n1353 0.00134872
R93729 VDD.n1600 VDD.n1334 0.00134872
R93730 VDD.n1473 VDD.n1351 0.00134872
R93731 VDD.n1601 VDD.n1335 0.00134872
R93732 VDD.n1474 VDD.n1350 0.00134872
R93733 VDD.n1602 VDD.n1336 0.00134872
R93734 VDD.n1475 VDD.n1348 0.00134872
R93735 VDD.n1603 VDD.n1337 0.00134872
R93736 VDD.n1476 VDD.n1347 0.00134872
R93737 VDD.n1604 VDD.n1338 0.00134872
R93738 VDD.n1477 VDD.n1345 0.00134872
R93739 VDD.n1605 VDD.n1339 0.00134872
R93740 VDD.n1478 VDD.n1344 0.00134872
R93741 VDD.n1606 VDD.n1340 0.00134872
R93742 VDD.n1479 VDD.n1342 0.00134872
R93743 VDD.n1341 VDD.n1194 0.00134872
R93744 VDD.n1479 VDD.n1341 0.00134872
R93745 VDD.n1478 VDD.n1340 0.00134872
R93746 VDD.n1477 VDD.n1339 0.00134872
R93747 VDD.n1476 VDD.n1338 0.00134872
R93748 VDD.n1475 VDD.n1337 0.00134872
R93749 VDD.n1474 VDD.n1336 0.00134872
R93750 VDD.n1473 VDD.n1335 0.00134872
R93751 VDD.n1472 VDD.n1334 0.00134872
R93752 VDD.n1471 VDD.n1333 0.00134872
R93753 VDD.n1470 VDD.n1332 0.00134872
R93754 VDD.n1469 VDD.n1331 0.00134872
R93755 VDD.n1468 VDD.n1330 0.00134872
R93756 VDD.n1467 VDD.n1329 0.00134872
R93757 VDD.n1466 VDD.n1328 0.00134872
R93758 VDD.n1465 VDD.n1327 0.00134872
R93759 VDD.n1464 VDD.n1326 0.00134872
R93760 VDD.n1463 VDD.n1325 0.00134872
R93761 VDD.n1462 VDD.n1324 0.00134872
R93762 VDD.n1461 VDD.n1323 0.00134872
R93763 VDD.n1460 VDD.n1322 0.00134872
R93764 VDD.n1459 VDD.n1321 0.00134872
R93765 VDD.n1458 VDD.n1320 0.00134872
R93766 VDD.n1457 VDD.n1319 0.00134872
R93767 VDD.n1456 VDD.n1318 0.00134872
R93768 VDD.n1455 VDD.n1316 0.00134872
R93769 VDD.n1454 VDD.n1315 0.00134872
R93770 VDD.n1453 VDD.n1313 0.00134872
R93771 VDD.n1452 VDD.n1312 0.00134872
R93772 VDD.n1451 VDD.n1310 0.00134872
R93773 VDD.n1450 VDD.n1309 0.00134872
R93774 VDD.n1449 VDD.n1307 0.00134872
R93775 VDD.n1448 VDD.n1306 0.00134872
R93776 VDD.n1447 VDD.n1304 0.00134872
R93777 VDD.n1446 VDD.n1303 0.00134872
R93778 VDD.n1445 VDD.n1301 0.00134872
R93779 VDD.n1444 VDD.n1300 0.00134872
R93780 VDD.n1443 VDD.n1298 0.00134872
R93781 VDD.n1442 VDD.n1297 0.00134872
R93782 VDD.n1441 VDD.n1295 0.00134872
R93783 VDD.n1440 VDD.n1294 0.00134872
R93784 VDD.n1439 VDD.n1292 0.00134872
R93785 VDD.n1438 VDD.n1291 0.00134872
R93786 VDD.n1437 VDD.n1289 0.00134872
R93787 VDD.n1436 VDD.n1288 0.00134872
R93788 VDD.n1435 VDD.n1286 0.00134872
R93789 VDD.n1434 VDD.n1285 0.00134872
R93790 VDD.n1433 VDD.n1283 0.00134872
R93791 VDD.n1432 VDD.n1282 0.00134872
R93792 VDD.n1431 VDD.n1280 0.00134872
R93793 VDD.n1430 VDD.n1279 0.00134872
R93794 VDD.n1429 VDD.n1277 0.00134872
R93795 VDD.n1428 VDD.n1276 0.00134872
R93796 VDD.n1427 VDD.n1274 0.00134872
R93797 VDD.n1426 VDD.n1273 0.00134872
R93798 VDD.n1425 VDD.n1271 0.00134872
R93799 VDD.n1424 VDD.n1270 0.00134872
R93800 VDD.n1423 VDD.n1268 0.00134872
R93801 VDD.n1422 VDD.n1267 0.00134872
R93802 VDD.n1421 VDD.n1265 0.00134872
R93803 VDD.n1420 VDD.n1264 0.00134872
R93804 VDD.n1419 VDD.n1262 0.00134872
R93805 VDD.n1418 VDD.n1261 0.00134872
R93806 VDD.n1544 VDD.n1481 0.00134872
R93807 VDD.n1671 VDD.n1417 0.00134872
R93808 VDD.n1607 VDD.n1195 0.00134872
R93809 VDD.n1606 VDD.n1342 0.00134872
R93810 VDD.n1605 VDD.n1344 0.00134872
R93811 VDD.n1604 VDD.n1345 0.00134872
R93812 VDD.n1603 VDD.n1347 0.00134872
R93813 VDD.n1602 VDD.n1348 0.00134872
R93814 VDD.n1601 VDD.n1350 0.00134872
R93815 VDD.n1600 VDD.n1351 0.00134872
R93816 VDD.n1599 VDD.n1353 0.00134872
R93817 VDD.n1598 VDD.n1354 0.00134872
R93818 VDD.n1597 VDD.n1356 0.00134872
R93819 VDD.n1596 VDD.n1357 0.00134872
R93820 VDD.n1595 VDD.n1359 0.00134872
R93821 VDD.n1594 VDD.n1360 0.00134872
R93822 VDD.n1593 VDD.n1362 0.00134872
R93823 VDD.n1592 VDD.n1363 0.00134872
R93824 VDD.n1591 VDD.n1365 0.00134872
R93825 VDD.n1590 VDD.n1366 0.00134872
R93826 VDD.n1589 VDD.n1368 0.00134872
R93827 VDD.n1588 VDD.n1369 0.00134872
R93828 VDD.n1587 VDD.n1371 0.00134872
R93829 VDD.n1586 VDD.n1372 0.00134872
R93830 VDD.n1585 VDD.n1374 0.00134872
R93831 VDD.n1584 VDD.n1375 0.00134872
R93832 VDD.n1583 VDD.n1376 0.00134872
R93833 VDD.n1582 VDD.n1377 0.00134872
R93834 VDD.n1581 VDD.n1378 0.00134872
R93835 VDD.n1580 VDD.n1379 0.00134872
R93836 VDD.n1579 VDD.n1380 0.00134872
R93837 VDD.n1578 VDD.n1381 0.00134872
R93838 VDD.n1577 VDD.n1382 0.00134872
R93839 VDD.n1576 VDD.n1383 0.00134872
R93840 VDD.n1575 VDD.n1384 0.00134872
R93841 VDD.n1574 VDD.n1385 0.00134872
R93842 VDD.n1573 VDD.n1386 0.00134872
R93843 VDD.n1572 VDD.n1387 0.00134872
R93844 VDD.n1571 VDD.n1388 0.00134872
R93845 VDD.n1570 VDD.n1389 0.00134872
R93846 VDD.n1569 VDD.n1390 0.00134872
R93847 VDD.n1568 VDD.n1391 0.00134872
R93848 VDD.n1567 VDD.n1392 0.00134872
R93849 VDD.n1566 VDD.n1393 0.00134872
R93850 VDD.n1565 VDD.n1394 0.00134872
R93851 VDD.n1564 VDD.n1395 0.00134872
R93852 VDD.n1563 VDD.n1396 0.00134872
R93853 VDD.n1562 VDD.n1397 0.00134872
R93854 VDD.n1561 VDD.n1398 0.00134872
R93855 VDD.n1560 VDD.n1399 0.00134872
R93856 VDD.n1559 VDD.n1400 0.00134872
R93857 VDD.n1558 VDD.n1401 0.00134872
R93858 VDD.n1557 VDD.n1402 0.00134872
R93859 VDD.n1556 VDD.n1403 0.00134872
R93860 VDD.n1555 VDD.n1404 0.00134872
R93861 VDD.n1554 VDD.n1405 0.00134872
R93862 VDD.n1553 VDD.n1406 0.00134872
R93863 VDD.n1552 VDD.n1407 0.00134872
R93864 VDD.n1551 VDD.n1408 0.00134872
R93865 VDD.n1550 VDD.n1409 0.00134872
R93866 VDD.n1549 VDD.n1410 0.00134872
R93867 VDD.n1548 VDD.n1411 0.00134872
R93868 VDD.n1547 VDD.n1412 0.00134872
R93869 VDD.n1546 VDD.n1413 0.00134872
R93870 VDD.n1545 VDD.n1414 0.00134872
R93871 VDD.n1670 VDD.n1607 0.00134872
R93872 VDD.n1676 VDD.n1194 0.00134872
R93873 VDD.n1482 VDD.n1416 0.00134872
R93874 VDD.n1669 VDD.n1196 0.00134872
R93875 VDD.n1483 VDD.n1193 0.00134872
R93876 VDD.n1668 VDD.n1197 0.00134872
R93877 VDD.n1484 VDD.n1192 0.00134872
R93878 VDD.n1667 VDD.n1198 0.00134872
R93879 VDD.n1485 VDD.n1191 0.00134872
R93880 VDD.n1666 VDD.n1199 0.00134872
R93881 VDD.n1486 VDD.n1190 0.00134872
R93882 VDD.n1665 VDD.n1200 0.00134872
R93883 VDD.n1487 VDD.n1189 0.00134872
R93884 VDD.n1664 VDD.n1201 0.00134872
R93885 VDD.n1488 VDD.n1188 0.00134872
R93886 VDD.n1663 VDD.n1202 0.00134872
R93887 VDD.n1489 VDD.n1187 0.00134872
R93888 VDD.n1662 VDD.n1203 0.00134872
R93889 VDD.n1490 VDD.n1186 0.00134872
R93890 VDD.n1661 VDD.n1204 0.00134872
R93891 VDD.n1491 VDD.n1185 0.00134872
R93892 VDD.n1660 VDD.n1205 0.00134872
R93893 VDD.n1492 VDD.n1184 0.00134872
R93894 VDD.n1659 VDD.n1206 0.00134872
R93895 VDD.n1493 VDD.n1183 0.00134872
R93896 VDD.n1658 VDD.n1207 0.00134872
R93897 VDD.n1494 VDD.n1182 0.00134872
R93898 VDD.n1657 VDD.n1208 0.00134872
R93899 VDD.n1495 VDD.n1181 0.00134872
R93900 VDD.n1656 VDD.n1209 0.00134872
R93901 VDD.n1496 VDD.n1180 0.00134872
R93902 VDD.n1655 VDD.n1210 0.00134872
R93903 VDD.n1497 VDD.n1179 0.00134872
R93904 VDD.n1654 VDD.n1211 0.00134872
R93905 VDD.n1498 VDD.n1178 0.00134872
R93906 VDD.n1653 VDD.n1212 0.00134872
R93907 VDD.n1499 VDD.n1177 0.00134872
R93908 VDD.n1652 VDD.n1213 0.00134872
R93909 VDD.n1500 VDD.n1176 0.00134872
R93910 VDD.n1651 VDD.n1214 0.00134872
R93911 VDD.n1501 VDD.n1175 0.00134872
R93912 VDD.n1650 VDD.n1215 0.00134872
R93913 VDD.n1502 VDD.n1174 0.00134872
R93914 VDD.n1649 VDD.n1216 0.00134872
R93915 VDD.n1503 VDD.n1173 0.00134872
R93916 VDD.n1648 VDD.n1217 0.00134872
R93917 VDD.n1504 VDD.n1172 0.00134872
R93918 VDD.n1647 VDD.n1218 0.00134872
R93919 VDD.n1505 VDD.n1171 0.00134872
R93920 VDD.n1646 VDD.n1219 0.00134872
R93921 VDD.n1506 VDD.n1170 0.00134872
R93922 VDD.n1645 VDD.n1220 0.00134872
R93923 VDD.n1507 VDD.n1169 0.00134872
R93924 VDD.n1644 VDD.n1221 0.00134872
R93925 VDD.n1508 VDD.n1168 0.00134872
R93926 VDD.n1643 VDD.n1222 0.00134872
R93927 VDD.n1509 VDD.n1167 0.00134872
R93928 VDD.n1642 VDD.n1223 0.00134872
R93929 VDD.n1510 VDD.n1166 0.00134872
R93930 VDD.n1641 VDD.n1224 0.00134872
R93931 VDD.n1511 VDD.n1165 0.00134872
R93932 VDD.n1640 VDD.n1225 0.00134872
R93933 VDD.n1512 VDD.n1164 0.00134872
R93934 VDD.n1639 VDD.n1226 0.00134872
R93935 VDD.n1513 VDD.n1163 0.00134872
R93936 VDD.n1638 VDD.n1227 0.00134872
R93937 VDD.n1514 VDD.n1162 0.00134872
R93938 VDD.n1637 VDD.n1228 0.00134872
R93939 VDD.n1515 VDD.n1161 0.00134872
R93940 VDD.n1636 VDD.n1229 0.00134872
R93941 VDD.n1516 VDD.n1160 0.00134872
R93942 VDD.n1635 VDD.n1230 0.00134872
R93943 VDD.n1517 VDD.n1159 0.00134872
R93944 VDD.n1634 VDD.n1231 0.00134872
R93945 VDD.n1518 VDD.n1158 0.00134872
R93946 VDD.n1633 VDD.n1232 0.00134872
R93947 VDD.n1519 VDD.n1157 0.00134872
R93948 VDD.n1632 VDD.n1233 0.00134872
R93949 VDD.n1520 VDD.n1156 0.00134872
R93950 VDD.n1631 VDD.n1234 0.00134872
R93951 VDD.n1521 VDD.n1155 0.00134872
R93952 VDD.n1630 VDD.n1235 0.00134872
R93953 VDD.n1522 VDD.n1154 0.00134872
R93954 VDD.n1629 VDD.n1236 0.00134872
R93955 VDD.n1523 VDD.n1153 0.00134872
R93956 VDD.n1628 VDD.n1237 0.00134872
R93957 VDD.n1524 VDD.n1152 0.00134872
R93958 VDD.n1627 VDD.n1238 0.00134872
R93959 VDD.n1525 VDD.n1151 0.00134872
R93960 VDD.n1626 VDD.n1239 0.00134872
R93961 VDD.n1526 VDD.n1150 0.00134872
R93962 VDD.n1625 VDD.n1240 0.00134872
R93963 VDD.n1527 VDD.n1149 0.00134872
R93964 VDD.n1624 VDD.n1241 0.00134872
R93965 VDD.n1528 VDD.n1148 0.00134872
R93966 VDD.n1623 VDD.n1242 0.00134872
R93967 VDD.n1529 VDD.n1147 0.00134872
R93968 VDD.n1622 VDD.n1243 0.00134872
R93969 VDD.n1530 VDD.n1146 0.00134872
R93970 VDD.n1621 VDD.n1244 0.00134872
R93971 VDD.n1531 VDD.n1145 0.00134872
R93972 VDD.n1620 VDD.n1245 0.00134872
R93973 VDD.n1532 VDD.n1144 0.00134872
R93974 VDD.n1619 VDD.n1246 0.00134872
R93975 VDD.n1533 VDD.n1143 0.00134872
R93976 VDD.n1618 VDD.n1247 0.00134872
R93977 VDD.n1534 VDD.n1142 0.00134872
R93978 VDD.n1617 VDD.n1248 0.00134872
R93979 VDD.n1535 VDD.n1141 0.00134872
R93980 VDD.n1616 VDD.n1249 0.00134872
R93981 VDD.n1536 VDD.n1140 0.00134872
R93982 VDD.n1615 VDD.n1250 0.00134872
R93983 VDD.n1537 VDD.n1139 0.00134872
R93984 VDD.n1614 VDD.n1251 0.00134872
R93985 VDD.n1538 VDD.n1138 0.00134872
R93986 VDD.n1613 VDD.n1252 0.00134872
R93987 VDD.n1539 VDD.n1137 0.00134872
R93988 VDD.n1612 VDD.n1253 0.00134872
R93989 VDD.n1540 VDD.n1136 0.00134872
R93990 VDD.n1611 VDD.n1254 0.00134872
R93991 VDD.n1541 VDD.n1135 0.00134872
R93992 VDD.n1610 VDD.n1255 0.00134872
R93993 VDD.n1542 VDD.n1134 0.00134872
R93994 VDD.n1609 VDD.n1256 0.00134872
R93995 VDD.n1543 VDD.n1133 0.00134872
R93996 VDD.n1608 VDD.n1257 0.00134872
R93997 VDD.n1258 VDD.n1132 0.00134872
R93998 VDD.n1675 VDD.n1259 0.00134872
R93999 VDD.n2 VDD.n0 0.00134303
R94000 VDD.n1679 VDD.n1678 0.00134303
R94001 VDD.n1671 VDD.n1415 0.0011975
R94002 VDD.n1673 VDD.n1672 0.0011975
R94003 VDD.n1672 VDD.n3 0.0011975
R94004 VDD.n4 VDD.n3 0.0011975
R94005 VDD.n5 VDD.n4 0.0011975
R94006 VDD.n1260 VDD.n5 0.0011975
R94007 VDD.n1260 VDD.n8 0.0011975
R94008 VDD.n9 VDD.n8 0.0011975
R94009 VDD.n10 VDD.n9 0.0011975
R94010 VDD.n1263 VDD.n10 0.0011975
R94011 VDD.n1263 VDD.n13 0.0011975
R94012 VDD.n14 VDD.n13 0.0011975
R94013 VDD.n15 VDD.n14 0.0011975
R94014 VDD.n1266 VDD.n15 0.0011975
R94015 VDD.n1266 VDD.n18 0.0011975
R94016 VDD.n19 VDD.n18 0.0011975
R94017 VDD.n20 VDD.n19 0.0011975
R94018 VDD.n1269 VDD.n20 0.0011975
R94019 VDD.n1269 VDD.n23 0.0011975
R94020 VDD.n24 VDD.n23 0.0011975
R94021 VDD.n25 VDD.n24 0.0011975
R94022 VDD.n1272 VDD.n25 0.0011975
R94023 VDD.n1272 VDD.n28 0.0011975
R94024 VDD.n29 VDD.n28 0.0011975
R94025 VDD.n30 VDD.n29 0.0011975
R94026 VDD.n1275 VDD.n30 0.0011975
R94027 VDD.n1275 VDD.n33 0.0011975
R94028 VDD.n34 VDD.n33 0.0011975
R94029 VDD.n35 VDD.n34 0.0011975
R94030 VDD.n1278 VDD.n35 0.0011975
R94031 VDD.n1278 VDD.n38 0.0011975
R94032 VDD.n39 VDD.n38 0.0011975
R94033 VDD.n40 VDD.n39 0.0011975
R94034 VDD.n1281 VDD.n40 0.0011975
R94035 VDD.n1281 VDD.n43 0.0011975
R94036 VDD.n44 VDD.n43 0.0011975
R94037 VDD.n45 VDD.n44 0.0011975
R94038 VDD.n1284 VDD.n45 0.0011975
R94039 VDD.n1284 VDD.n48 0.0011975
R94040 VDD.n49 VDD.n48 0.0011975
R94041 VDD.n50 VDD.n49 0.0011975
R94042 VDD.n1287 VDD.n50 0.0011975
R94043 VDD.n1287 VDD.n53 0.0011975
R94044 VDD.n54 VDD.n53 0.0011975
R94045 VDD.n55 VDD.n54 0.0011975
R94046 VDD.n1290 VDD.n55 0.0011975
R94047 VDD.n1290 VDD.n58 0.0011975
R94048 VDD.n59 VDD.n58 0.0011975
R94049 VDD.n60 VDD.n59 0.0011975
R94050 VDD.n1293 VDD.n60 0.0011975
R94051 VDD.n1293 VDD.n63 0.0011975
R94052 VDD.n64 VDD.n63 0.0011975
R94053 VDD.n65 VDD.n64 0.0011975
R94054 VDD.n1296 VDD.n65 0.0011975
R94055 VDD.n1296 VDD.n68 0.0011975
R94056 VDD.n69 VDD.n68 0.0011975
R94057 VDD.n70 VDD.n69 0.0011975
R94058 VDD.n1299 VDD.n70 0.0011975
R94059 VDD.n1299 VDD.n73 0.0011975
R94060 VDD.n74 VDD.n73 0.0011975
R94061 VDD.n75 VDD.n74 0.0011975
R94062 VDD.n1302 VDD.n75 0.0011975
R94063 VDD.n1302 VDD.n78 0.0011975
R94064 VDD.n79 VDD.n78 0.0011975
R94065 VDD.n80 VDD.n79 0.0011975
R94066 VDD.n1305 VDD.n80 0.0011975
R94067 VDD.n1305 VDD.n83 0.0011975
R94068 VDD.n84 VDD.n83 0.0011975
R94069 VDD.n85 VDD.n84 0.0011975
R94070 VDD.n1308 VDD.n85 0.0011975
R94071 VDD.n1308 VDD.n88 0.0011975
R94072 VDD.n89 VDD.n88 0.0011975
R94073 VDD.n90 VDD.n89 0.0011975
R94074 VDD.n1311 VDD.n90 0.0011975
R94075 VDD.n1311 VDD.n93 0.0011975
R94076 VDD.n94 VDD.n93 0.0011975
R94077 VDD.n95 VDD.n94 0.0011975
R94078 VDD.n1314 VDD.n95 0.0011975
R94079 VDD.n1314 VDD.n98 0.0011975
R94080 VDD.n99 VDD.n98 0.0011975
R94081 VDD.n100 VDD.n99 0.0011975
R94082 VDD.n1317 VDD.n100 0.0011975
R94083 VDD.n1317 VDD.n102 0.0011975
R94084 VDD.n103 VDD.n102 0.0011975
R94085 VDD.n1373 VDD.n103 0.0011975
R94086 VDD.n1373 VDD.n106 0.0011975
R94087 VDD.n107 VDD.n106 0.0011975
R94088 VDD.n108 VDD.n107 0.0011975
R94089 VDD.n1370 VDD.n108 0.0011975
R94090 VDD.n1370 VDD.n111 0.0011975
R94091 VDD.n112 VDD.n111 0.0011975
R94092 VDD.n113 VDD.n112 0.0011975
R94093 VDD.n1367 VDD.n113 0.0011975
R94094 VDD.n1367 VDD.n116 0.0011975
R94095 VDD.n117 VDD.n116 0.0011975
R94096 VDD.n118 VDD.n117 0.0011975
R94097 VDD.n1364 VDD.n118 0.0011975
R94098 VDD.n1364 VDD.n121 0.0011975
R94099 VDD.n122 VDD.n121 0.0011975
R94100 VDD.n123 VDD.n122 0.0011975
R94101 VDD.n1361 VDD.n123 0.0011975
R94102 VDD.n1361 VDD.n126 0.0011975
R94103 VDD.n127 VDD.n126 0.0011975
R94104 VDD.n128 VDD.n127 0.0011975
R94105 VDD.n1358 VDD.n128 0.0011975
R94106 VDD.n1358 VDD.n131 0.0011975
R94107 VDD.n132 VDD.n131 0.0011975
R94108 VDD.n133 VDD.n132 0.0011975
R94109 VDD.n1355 VDD.n133 0.0011975
R94110 VDD.n1355 VDD.n136 0.0011975
R94111 VDD.n137 VDD.n136 0.0011975
R94112 VDD.n138 VDD.n137 0.0011975
R94113 VDD.n1352 VDD.n138 0.0011975
R94114 VDD.n1352 VDD.n141 0.0011975
R94115 VDD.n142 VDD.n141 0.0011975
R94116 VDD.n143 VDD.n142 0.0011975
R94117 VDD.n1349 VDD.n143 0.0011975
R94118 VDD.n1349 VDD.n146 0.0011975
R94119 VDD.n147 VDD.n146 0.0011975
R94120 VDD.n148 VDD.n147 0.0011975
R94121 VDD.n1346 VDD.n148 0.0011975
R94122 VDD.n1346 VDD.n151 0.0011975
R94123 VDD.n152 VDD.n151 0.0011975
R94124 VDD.n153 VDD.n152 0.0011975
R94125 VDD.n1343 VDD.n153 0.0011975
R94126 VDD.n1343 VDD.n156 0.0011975
R94127 VDD.n157 VDD.n156 0.0011975
R94128 VDD.n158 VDD.n157 0.0011975
R94129 VDD.n1677 VDD.n158 0.0011975
R94130 VDD.n1866 VDD.n2 0.0011975
R94131 VDD.n1866 VDD.n1865 0.0011975
R94132 VDD.n1865 VDD.n1864 0.0011975
R94133 VDD.n1864 VDD.n6 0.0011975
R94134 VDD.n1860 VDD.n6 0.0011975
R94135 VDD.n1860 VDD.n1859 0.0011975
R94136 VDD.n1859 VDD.n1858 0.0011975
R94137 VDD.n1858 VDD.n11 0.0011975
R94138 VDD.n1854 VDD.n11 0.0011975
R94139 VDD.n1854 VDD.n1853 0.0011975
R94140 VDD.n1853 VDD.n1852 0.0011975
R94141 VDD.n1852 VDD.n16 0.0011975
R94142 VDD.n1848 VDD.n16 0.0011975
R94143 VDD.n1848 VDD.n1847 0.0011975
R94144 VDD.n1847 VDD.n1846 0.0011975
R94145 VDD.n1846 VDD.n21 0.0011975
R94146 VDD.n1842 VDD.n21 0.0011975
R94147 VDD.n1842 VDD.n1841 0.0011975
R94148 VDD.n1841 VDD.n1840 0.0011975
R94149 VDD.n1840 VDD.n26 0.0011975
R94150 VDD.n1836 VDD.n26 0.0011975
R94151 VDD.n1836 VDD.n1835 0.0011975
R94152 VDD.n1835 VDD.n1834 0.0011975
R94153 VDD.n1834 VDD.n31 0.0011975
R94154 VDD.n1830 VDD.n31 0.0011975
R94155 VDD.n1830 VDD.n1829 0.0011975
R94156 VDD.n1829 VDD.n1828 0.0011975
R94157 VDD.n1828 VDD.n36 0.0011975
R94158 VDD.n1824 VDD.n36 0.0011975
R94159 VDD.n1824 VDD.n1823 0.0011975
R94160 VDD.n1823 VDD.n1822 0.0011975
R94161 VDD.n1822 VDD.n41 0.0011975
R94162 VDD.n1818 VDD.n41 0.0011975
R94163 VDD.n1818 VDD.n1817 0.0011975
R94164 VDD.n1817 VDD.n1816 0.0011975
R94165 VDD.n1816 VDD.n46 0.0011975
R94166 VDD.n1812 VDD.n46 0.0011975
R94167 VDD.n1812 VDD.n1811 0.0011975
R94168 VDD.n1811 VDD.n1810 0.0011975
R94169 VDD.n1810 VDD.n51 0.0011975
R94170 VDD.n1806 VDD.n51 0.0011975
R94171 VDD.n1806 VDD.n1805 0.0011975
R94172 VDD.n1805 VDD.n1804 0.0011975
R94173 VDD.n1804 VDD.n56 0.0011975
R94174 VDD.n1800 VDD.n56 0.0011975
R94175 VDD.n1800 VDD.n1799 0.0011975
R94176 VDD.n1799 VDD.n1798 0.0011975
R94177 VDD.n1798 VDD.n61 0.0011975
R94178 VDD.n1794 VDD.n61 0.0011975
R94179 VDD.n1794 VDD.n1793 0.0011975
R94180 VDD.n1793 VDD.n1792 0.0011975
R94181 VDD.n1792 VDD.n66 0.0011975
R94182 VDD.n1788 VDD.n66 0.0011975
R94183 VDD.n1788 VDD.n1787 0.0011975
R94184 VDD.n1787 VDD.n1786 0.0011975
R94185 VDD.n1786 VDD.n71 0.0011975
R94186 VDD.n1782 VDD.n71 0.0011975
R94187 VDD.n1782 VDD.n1781 0.0011975
R94188 VDD.n1781 VDD.n1780 0.0011975
R94189 VDD.n1780 VDD.n76 0.0011975
R94190 VDD.n1776 VDD.n76 0.0011975
R94191 VDD.n1776 VDD.n1775 0.0011975
R94192 VDD.n1775 VDD.n1774 0.0011975
R94193 VDD.n1774 VDD.n81 0.0011975
R94194 VDD.n1770 VDD.n81 0.0011975
R94195 VDD.n1770 VDD.n1769 0.0011975
R94196 VDD.n1769 VDD.n1768 0.0011975
R94197 VDD.n1768 VDD.n86 0.0011975
R94198 VDD.n1764 VDD.n86 0.0011975
R94199 VDD.n1764 VDD.n1763 0.0011975
R94200 VDD.n1763 VDD.n1762 0.0011975
R94201 VDD.n1762 VDD.n91 0.0011975
R94202 VDD.n1758 VDD.n91 0.0011975
R94203 VDD.n1758 VDD.n1757 0.0011975
R94204 VDD.n1757 VDD.n1756 0.0011975
R94205 VDD.n1756 VDD.n96 0.0011975
R94206 VDD.n1752 VDD.n96 0.0011975
R94207 VDD.n1752 VDD.n1751 0.0011975
R94208 VDD.n1751 VDD.n1750 0.0011975
R94209 VDD.n1750 VDD.n101 0.0011975
R94210 VDD.n1746 VDD.n101 0.0011975
R94211 VDD.n1746 VDD.n1745 0.0011975
R94212 VDD.n1745 VDD.n104 0.0011975
R94213 VDD.n1741 VDD.n104 0.0011975
R94214 VDD.n1741 VDD.n1740 0.0011975
R94215 VDD.n1740 VDD.n1739 0.0011975
R94216 VDD.n1739 VDD.n109 0.0011975
R94217 VDD.n1735 VDD.n109 0.0011975
R94218 VDD.n1735 VDD.n1734 0.0011975
R94219 VDD.n1734 VDD.n1733 0.0011975
R94220 VDD.n1733 VDD.n114 0.0011975
R94221 VDD.n1729 VDD.n114 0.0011975
R94222 VDD.n1729 VDD.n1728 0.0011975
R94223 VDD.n1728 VDD.n1727 0.0011975
R94224 VDD.n1727 VDD.n119 0.0011975
R94225 VDD.n1723 VDD.n119 0.0011975
R94226 VDD.n1723 VDD.n1722 0.0011975
R94227 VDD.n1722 VDD.n1721 0.0011975
R94228 VDD.n1721 VDD.n124 0.0011975
R94229 VDD.n1717 VDD.n124 0.0011975
R94230 VDD.n1717 VDD.n1716 0.0011975
R94231 VDD.n1716 VDD.n1715 0.0011975
R94232 VDD.n1715 VDD.n129 0.0011975
R94233 VDD.n1711 VDD.n129 0.0011975
R94234 VDD.n1711 VDD.n1710 0.0011975
R94235 VDD.n1710 VDD.n1709 0.0011975
R94236 VDD.n1709 VDD.n134 0.0011975
R94237 VDD.n1705 VDD.n134 0.0011975
R94238 VDD.n1705 VDD.n1704 0.0011975
R94239 VDD.n1704 VDD.n1703 0.0011975
R94240 VDD.n1703 VDD.n139 0.0011975
R94241 VDD.n1699 VDD.n139 0.0011975
R94242 VDD.n1699 VDD.n1698 0.0011975
R94243 VDD.n1698 VDD.n1697 0.0011975
R94244 VDD.n1697 VDD.n144 0.0011975
R94245 VDD.n1693 VDD.n144 0.0011975
R94246 VDD.n1693 VDD.n1692 0.0011975
R94247 VDD.n1692 VDD.n1691 0.0011975
R94248 VDD.n1691 VDD.n149 0.0011975
R94249 VDD.n1687 VDD.n149 0.0011975
R94250 VDD.n1687 VDD.n1686 0.0011975
R94251 VDD.n1686 VDD.n1685 0.0011975
R94252 VDD.n1685 VDD.n154 0.0011975
R94253 VDD.n1681 VDD.n154 0.0011975
R94254 VDD.n1681 VDD.n1680 0.0011975
R94255 VDD.n1680 VDD.n1679 0.0011975
R94256 VDD.n1867 VDD.n1 0.000965
R94257 VDD.n1863 VDD.n1 0.000965
R94258 VDD.n1863 VDD.n1862 0.000965
R94259 VDD.n1862 VDD.n1861 0.000965
R94260 VDD.n1861 VDD.n7 0.000965
R94261 VDD.n1857 VDD.n7 0.000965
R94262 VDD.n1857 VDD.n1856 0.000965
R94263 VDD.n1856 VDD.n1855 0.000965
R94264 VDD.n1855 VDD.n12 0.000965
R94265 VDD.n1851 VDD.n12 0.000965
R94266 VDD.n1851 VDD.n1850 0.000965
R94267 VDD.n1850 VDD.n1849 0.000965
R94268 VDD.n1849 VDD.n17 0.000965
R94269 VDD.n1845 VDD.n17 0.000965
R94270 VDD.n1845 VDD.n1844 0.000965
R94271 VDD.n1844 VDD.n1843 0.000965
R94272 VDD.n1843 VDD.n22 0.000965
R94273 VDD.n1839 VDD.n22 0.000965
R94274 VDD.n1839 VDD.n1838 0.000965
R94275 VDD.n1838 VDD.n1837 0.000965
R94276 VDD.n1837 VDD.n27 0.000965
R94277 VDD.n1833 VDD.n27 0.000965
R94278 VDD.n1833 VDD.n1832 0.000965
R94279 VDD.n1832 VDD.n1831 0.000965
R94280 VDD.n1831 VDD.n32 0.000965
R94281 VDD.n1827 VDD.n32 0.000965
R94282 VDD.n1827 VDD.n1826 0.000965
R94283 VDD.n1826 VDD.n1825 0.000965
R94284 VDD.n1825 VDD.n37 0.000965
R94285 VDD.n1821 VDD.n37 0.000965
R94286 VDD.n1821 VDD.n1820 0.000965
R94287 VDD.n1820 VDD.n1819 0.000965
R94288 VDD.n1819 VDD.n42 0.000965
R94289 VDD.n1815 VDD.n42 0.000965
R94290 VDD.n1815 VDD.n1814 0.000965
R94291 VDD.n1814 VDD.n1813 0.000965
R94292 VDD.n1813 VDD.n47 0.000965
R94293 VDD.n1809 VDD.n47 0.000965
R94294 VDD.n1809 VDD.n1808 0.000965
R94295 VDD.n1808 VDD.n1807 0.000965
R94296 VDD.n1807 VDD.n52 0.000965
R94297 VDD.n1803 VDD.n52 0.000965
R94298 VDD.n1803 VDD.n1802 0.000965
R94299 VDD.n1802 VDD.n1801 0.000965
R94300 VDD.n1801 VDD.n57 0.000965
R94301 VDD.n1797 VDD.n57 0.000965
R94302 VDD.n1797 VDD.n1796 0.000965
R94303 VDD.n1796 VDD.n1795 0.000965
R94304 VDD.n1795 VDD.n62 0.000965
R94305 VDD.n1791 VDD.n62 0.000965
R94306 VDD.n1791 VDD.n1790 0.000965
R94307 VDD.n1790 VDD.n1789 0.000965
R94308 VDD.n1789 VDD.n67 0.000965
R94309 VDD.n1785 VDD.n67 0.000965
R94310 VDD.n1785 VDD.n1784 0.000965
R94311 VDD.n1784 VDD.n1783 0.000965
R94312 VDD.n1783 VDD.n72 0.000965
R94313 VDD.n1779 VDD.n72 0.000965
R94314 VDD.n1779 VDD.n1778 0.000965
R94315 VDD.n1778 VDD.n1777 0.000965
R94316 VDD.n1777 VDD.n77 0.000965
R94317 VDD.n1773 VDD.n77 0.000965
R94318 VDD.n1773 VDD.n1772 0.000965
R94319 VDD.n1772 VDD.n1771 0.000965
R94320 VDD.n1771 VDD.n82 0.000965
R94321 VDD.n1767 VDD.n82 0.000965
R94322 VDD.n1767 VDD.n1766 0.000965
R94323 VDD.n1766 VDD.n1765 0.000965
R94324 VDD.n1765 VDD.n87 0.000965
R94325 VDD.n1761 VDD.n87 0.000965
R94326 VDD.n1761 VDD.n1760 0.000965
R94327 VDD.n1760 VDD.n1759 0.000965
R94328 VDD.n1759 VDD.n92 0.000965
R94329 VDD.n1755 VDD.n92 0.000965
R94330 VDD.n1755 VDD.n1754 0.000965
R94331 VDD.n1754 VDD.n1753 0.000965
R94332 VDD.n1753 VDD.n97 0.000965
R94333 VDD.n1749 VDD.n97 0.000965
R94334 VDD.n1749 VDD.n1748 0.000965
R94335 VDD.n1748 VDD.n1747 0.000965
R94336 VDD.n1744 VDD.n1743 0.000965
R94337 VDD.n1743 VDD.n1742 0.000965
R94338 VDD.n1742 VDD.n105 0.000965
R94339 VDD.n1738 VDD.n105 0.000965
R94340 VDD.n1738 VDD.n1737 0.000965
R94341 VDD.n1737 VDD.n1736 0.000965
R94342 VDD.n1736 VDD.n110 0.000965
R94343 VDD.n1732 VDD.n110 0.000965
R94344 VDD.n1732 VDD.n1731 0.000965
R94345 VDD.n1731 VDD.n1730 0.000965
R94346 VDD.n1730 VDD.n115 0.000965
R94347 VDD.n1726 VDD.n115 0.000965
R94348 VDD.n1726 VDD.n1725 0.000965
R94349 VDD.n1725 VDD.n1724 0.000965
R94350 VDD.n1724 VDD.n120 0.000965
R94351 VDD.n1720 VDD.n120 0.000965
R94352 VDD.n1720 VDD.n1719 0.000965
R94353 VDD.n1719 VDD.n1718 0.000965
R94354 VDD.n1718 VDD.n125 0.000965
R94355 VDD.n1714 VDD.n125 0.000965
R94356 VDD.n1714 VDD.n1713 0.000965
R94357 VDD.n1713 VDD.n1712 0.000965
R94358 VDD.n1712 VDD.n130 0.000965
R94359 VDD.n1708 VDD.n130 0.000965
R94360 VDD.n1708 VDD.n1707 0.000965
R94361 VDD.n1707 VDD.n1706 0.000965
R94362 VDD.n1706 VDD.n135 0.000965
R94363 VDD.n1702 VDD.n135 0.000965
R94364 VDD.n1702 VDD.n1701 0.000965
R94365 VDD.n1701 VDD.n1700 0.000965
R94366 VDD.n1700 VDD.n140 0.000965
R94367 VDD.n1696 VDD.n140 0.000965
R94368 VDD.n1696 VDD.n1695 0.000965
R94369 VDD.n1695 VDD.n1694 0.000965
R94370 VDD.n1694 VDD.n145 0.000965
R94371 VDD.n1690 VDD.n145 0.000965
R94372 VDD.n1690 VDD.n1689 0.000965
R94373 VDD.n1689 VDD.n1688 0.000965
R94374 VDD.n1688 VDD.n150 0.000965
R94375 VDD.n1684 VDD.n150 0.000965
R94376 VDD.n1684 VDD.n1683 0.000965
R94377 VDD.n1683 VDD.n1682 0.000965
R94378 VDD.n1682 VDD.n155 0.000965
R94379 VDD.n1747 VDD 0.00089
R94380 VDD.n1744 VDD 0.000575
C0 m2_434_n43048 VDD 48.0842f
C1 VDD IB 11.054f
C2 m2_434_n43048 IB 2.82537f
C3 VDD VINN 0.324965f
C4 VSS OUT 6.66314f
C5 m2_434_n43048 VINN 1.7813f
C6 IB VINN 0.159398f
C7 VSS VINP 1.48414f
C8 OUT VINP 0.172917f
C9 m2_434_n43048 VSS 1.00695f
C10 VSS IB 0.142004f
C11 VDD OUT 4.85827f
C12 m2_434_n43048 OUT 1.01343f
C13 a_n1924_n46660 VSS 0.940194f
C14 VSS VINN 1.6342f
C15 IB OUT 2.86622f
C16 VDD VINP 0.224928f
C17 m2_434_n43048 VINP 0.835684f
C18 VINP a_n3166_n47928 0.101706p
C19 VINN a_n3166_n47928 0.101888p
C20 OUT a_n3166_n47928 87.6969f
C21 IB a_n3166_n47928 81.075f
C22 VSS a_n3166_n47928 0.523001p
C23 VDD a_n3166_n47928 0.348713p
C24 m2_434_n43048 a_n3166_n47928 15.489f $ **FLOATING
C25 a_n1924_n46660 a_n3166_n47928 1.48755f
C26 VDD.n0 a_n3166_n47928 0.107553f
C27 VDD.n1 a_n3166_n47928 0.101866f
C28 VDD.n2 a_n3166_n47928 0.101866f
C29 VDD.n3 a_n3166_n47928 0.101866f
C30 VDD.n4 a_n3166_n47928 0.101866f
C31 VDD.n5 a_n3166_n47928 0.101866f
C32 VDD.n6 a_n3166_n47928 0.101866f
C33 VDD.n7 a_n3166_n47928 0.101866f
C34 VDD.n8 a_n3166_n47928 0.101866f
C35 VDD.n9 a_n3166_n47928 0.101866f
C36 VDD.n10 a_n3166_n47928 0.101866f
C37 VDD.n11 a_n3166_n47928 0.101866f
C38 VDD.n12 a_n3166_n47928 0.101866f
C39 VDD.n13 a_n3166_n47928 0.101866f
C40 VDD.n14 a_n3166_n47928 0.101866f
C41 VDD.n15 a_n3166_n47928 0.101866f
C42 VDD.n16 a_n3166_n47928 0.101866f
C43 VDD.n17 a_n3166_n47928 0.101866f
C44 VDD.n18 a_n3166_n47928 0.101866f
C45 VDD.n19 a_n3166_n47928 0.101866f
C46 VDD.n20 a_n3166_n47928 0.101866f
C47 VDD.n21 a_n3166_n47928 0.101866f
C48 VDD.n22 a_n3166_n47928 0.101866f
C49 VDD.n23 a_n3166_n47928 0.101866f
C50 VDD.n24 a_n3166_n47928 0.101866f
C51 VDD.n25 a_n3166_n47928 0.101866f
C52 VDD.n26 a_n3166_n47928 0.101866f
C53 VDD.n27 a_n3166_n47928 0.101866f
C54 VDD.n28 a_n3166_n47928 0.101866f
C55 VDD.n29 a_n3166_n47928 0.101866f
C56 VDD.n30 a_n3166_n47928 0.101866f
C57 VDD.n31 a_n3166_n47928 0.101866f
C58 VDD.n32 a_n3166_n47928 0.101866f
C59 VDD.n33 a_n3166_n47928 0.101866f
C60 VDD.n34 a_n3166_n47928 0.101866f
C61 VDD.n35 a_n3166_n47928 0.101866f
C62 VDD.n36 a_n3166_n47928 0.101866f
C63 VDD.n37 a_n3166_n47928 0.101866f
C64 VDD.n38 a_n3166_n47928 0.101866f
C65 VDD.n39 a_n3166_n47928 0.101866f
C66 VDD.n40 a_n3166_n47928 0.101866f
C67 VDD.n41 a_n3166_n47928 0.101866f
C68 VDD.n42 a_n3166_n47928 0.101866f
C69 VDD.n43 a_n3166_n47928 0.101866f
C70 VDD.n44 a_n3166_n47928 0.101866f
C71 VDD.n45 a_n3166_n47928 0.101866f
C72 VDD.n46 a_n3166_n47928 0.101866f
C73 VDD.n47 a_n3166_n47928 0.101866f
C74 VDD.n48 a_n3166_n47928 0.101866f
C75 VDD.n49 a_n3166_n47928 0.101866f
C76 VDD.n50 a_n3166_n47928 0.101866f
C77 VDD.n51 a_n3166_n47928 0.101866f
C78 VDD.n52 a_n3166_n47928 0.101866f
C79 VDD.n53 a_n3166_n47928 0.101866f
C80 VDD.n54 a_n3166_n47928 0.101866f
C81 VDD.n55 a_n3166_n47928 0.101866f
C82 VDD.n56 a_n3166_n47928 0.101866f
C83 VDD.n57 a_n3166_n47928 0.101866f
C84 VDD.n58 a_n3166_n47928 0.101866f
C85 VDD.n59 a_n3166_n47928 0.101866f
C86 VDD.n60 a_n3166_n47928 0.101866f
C87 VDD.n61 a_n3166_n47928 0.101866f
C88 VDD.n62 a_n3166_n47928 0.101866f
C89 VDD.n63 a_n3166_n47928 0.101866f
C90 VDD.n64 a_n3166_n47928 0.101866f
C91 VDD.n65 a_n3166_n47928 0.101866f
C92 VDD.n66 a_n3166_n47928 0.101866f
C93 VDD.n67 a_n3166_n47928 0.101866f
C94 VDD.n68 a_n3166_n47928 0.101866f
C95 VDD.n69 a_n3166_n47928 0.101866f
C96 VDD.n70 a_n3166_n47928 0.101866f
C97 VDD.n71 a_n3166_n47928 0.101866f
C98 VDD.n72 a_n3166_n47928 0.101866f
C99 VDD.n73 a_n3166_n47928 0.101866f
C100 VDD.n74 a_n3166_n47928 0.101866f
C101 VDD.n75 a_n3166_n47928 0.101866f
C102 VDD.n76 a_n3166_n47928 0.101866f
C103 VDD.n77 a_n3166_n47928 0.101866f
C104 VDD.n78 a_n3166_n47928 0.101866f
C105 VDD.n79 a_n3166_n47928 0.101866f
C106 VDD.n80 a_n3166_n47928 0.101866f
C107 VDD.n81 a_n3166_n47928 0.101866f
C108 VDD.n82 a_n3166_n47928 0.101866f
C109 VDD.n83 a_n3166_n47928 0.101866f
C110 VDD.n84 a_n3166_n47928 0.101866f
C111 VDD.n85 a_n3166_n47928 0.101866f
C112 VDD.n86 a_n3166_n47928 0.101866f
C113 VDD.n87 a_n3166_n47928 0.101866f
C114 VDD.n88 a_n3166_n47928 0.101866f
C115 VDD.n89 a_n3166_n47928 0.101866f
C116 VDD.n90 a_n3166_n47928 0.101866f
C117 VDD.n91 a_n3166_n47928 0.101866f
C118 VDD.n92 a_n3166_n47928 0.101866f
C119 VDD.n93 a_n3166_n47928 0.101866f
C120 VDD.n94 a_n3166_n47928 0.101866f
C121 VDD.n95 a_n3166_n47928 0.101866f
C122 VDD.n96 a_n3166_n47928 0.101866f
C123 VDD.n97 a_n3166_n47928 0.101866f
C124 VDD.n98 a_n3166_n47928 0.101866f
C125 VDD.n99 a_n3166_n47928 0.101866f
C126 VDD.n100 a_n3166_n47928 0.101866f
C127 VDD.n101 a_n3166_n47928 0.101866f
C128 VDD.n102 a_n3166_n47928 0.101866f
C129 VDD.n103 a_n3166_n47928 0.101866f
C130 VDD.n104 a_n3166_n47928 0.101866f
C131 VDD.n105 a_n3166_n47928 0.101866f
C132 VDD.n106 a_n3166_n47928 0.101866f
C133 VDD.n107 a_n3166_n47928 0.101866f
C134 VDD.n108 a_n3166_n47928 0.101866f
C135 VDD.n109 a_n3166_n47928 0.101866f
C136 VDD.n110 a_n3166_n47928 0.101866f
C137 VDD.n111 a_n3166_n47928 0.101866f
C138 VDD.n112 a_n3166_n47928 0.101866f
C139 VDD.n113 a_n3166_n47928 0.101866f
C140 VDD.n114 a_n3166_n47928 0.101866f
C141 VDD.n115 a_n3166_n47928 0.101866f
C142 VDD.n116 a_n3166_n47928 0.101866f
C143 VDD.n117 a_n3166_n47928 0.101866f
C144 VDD.n118 a_n3166_n47928 0.101866f
C145 VDD.n119 a_n3166_n47928 0.101866f
C146 VDD.n120 a_n3166_n47928 0.101866f
C147 VDD.n121 a_n3166_n47928 0.101866f
C148 VDD.n122 a_n3166_n47928 0.101866f
C149 VDD.n123 a_n3166_n47928 0.101866f
C150 VDD.n124 a_n3166_n47928 0.101866f
C151 VDD.n125 a_n3166_n47928 0.101866f
C152 VDD.n126 a_n3166_n47928 0.101866f
C153 VDD.n127 a_n3166_n47928 0.101866f
C154 VDD.n128 a_n3166_n47928 0.101866f
C155 VDD.n129 a_n3166_n47928 0.101866f
C156 VDD.n130 a_n3166_n47928 0.101866f
C157 VDD.n131 a_n3166_n47928 0.101866f
C158 VDD.n132 a_n3166_n47928 0.101866f
C159 VDD.n133 a_n3166_n47928 0.101866f
C160 VDD.n134 a_n3166_n47928 0.101866f
C161 VDD.n135 a_n3166_n47928 0.101866f
C162 VDD.n136 a_n3166_n47928 0.101866f
C163 VDD.n137 a_n3166_n47928 0.101866f
C164 VDD.n138 a_n3166_n47928 0.101866f
C165 VDD.n139 a_n3166_n47928 0.101866f
C166 VDD.n140 a_n3166_n47928 0.101866f
C167 VDD.n141 a_n3166_n47928 0.101866f
C168 VDD.n142 a_n3166_n47928 0.101866f
C169 VDD.n143 a_n3166_n47928 0.101866f
C170 VDD.n144 a_n3166_n47928 0.101866f
C171 VDD.n145 a_n3166_n47928 0.101866f
C172 VDD.n146 a_n3166_n47928 0.101866f
C173 VDD.n147 a_n3166_n47928 0.101866f
C174 VDD.n148 a_n3166_n47928 0.101866f
C175 VDD.n149 a_n3166_n47928 0.101866f
C176 VDD.n150 a_n3166_n47928 0.101866f
C177 VDD.n151 a_n3166_n47928 0.101866f
C178 VDD.n152 a_n3166_n47928 0.101866f
C179 VDD.n153 a_n3166_n47928 0.101866f
C180 VDD.n154 a_n3166_n47928 0.101866f
C181 VDD.n155 a_n3166_n47928 0.300709f
C182 VDD.n156 a_n3166_n47928 0.101866f
C183 VDD.n157 a_n3166_n47928 0.101866f
C184 VDD.n158 a_n3166_n47928 0.101866f
C185 VDD.n403 a_n3166_n47928 0.025309f
C186 VDD.n405 a_n3166_n47928 0.025309f
C187 VDD.t28 a_n3166_n47928 0.014879f
C188 VDD.n669 a_n3166_n47928 0.011112f
C189 VDD.n670 a_n3166_n47928 0.011112f
C190 VDD.n718 a_n3166_n47928 0.025309f
C191 VDD.t16 a_n3166_n47928 0.014879f
C192 VDD.t30 a_n3166_n47928 0.014879f
C193 VDD.n720 a_n3166_n47928 0.025309f
C194 VDD.n731 a_n3166_n47928 0.026181f
C195 VDD.t14 a_n3166_n47928 0.018416f
C196 VDD.t38 a_n3166_n47928 0.010613f
C197 VDD.t44 a_n3166_n47928 0.010613f
C198 VDD.t2 a_n3166_n47928 0.018416f
C199 VDD.n733 a_n3166_n47928 0.026181f
C200 VDD.n764 a_n3166_n47928 0.032995f
C201 VDD.t46 a_n3166_n47928 0.018416f
C202 VDD.t54 a_n3166_n47928 0.014151f
C203 VDD.t34 a_n3166_n47928 0.014151f
C204 VDD.t20 a_n3166_n47928 0.014151f
C205 VDD.t48 a_n3166_n47928 0.014151f
C206 VDD.t18 a_n3166_n47928 0.014151f
C207 VDD.t36 a_n3166_n47928 0.014151f
C208 VDD.t12 a_n3166_n47928 0.014151f
C209 VDD.t8 a_n3166_n47928 0.014151f
C210 VDD.t24 a_n3166_n47928 0.010613f
C211 VDD.t6 a_n3166_n47928 0.010613f
C212 VDD.t22 a_n3166_n47928 0.014151f
C213 VDD.t32 a_n3166_n47928 0.014151f
C214 VDD.t50 a_n3166_n47928 0.014151f
C215 VDD.t4 a_n3166_n47928 0.014151f
C216 VDD.t40 a_n3166_n47928 0.014151f
C217 VDD.t0 a_n3166_n47928 0.014151f
C218 VDD.t10 a_n3166_n47928 0.014151f
C219 VDD.t26 a_n3166_n47928 0.014151f
C220 VDD.t42 a_n3166_n47928 0.018416f
C221 VDD.n766 a_n3166_n47928 0.032995f
C222 VDD.t52 a_n3166_n47928 0.014879f
C223 VDD.n1129 a_n3166_n47928 0.013801f
C224 VDD.n1130 a_n3166_n47928 0.808283f
C225 VDD.n1131 a_n3166_n47928 0.898875f
C226 VDD.n1132 a_n3166_n47928 0.101866f
C227 VDD.n1133 a_n3166_n47928 0.101866f
C228 VDD.n1134 a_n3166_n47928 0.101866f
C229 VDD.n1135 a_n3166_n47928 0.101866f
C230 VDD.n1136 a_n3166_n47928 0.101866f
C231 VDD.n1137 a_n3166_n47928 0.101866f
C232 VDD.n1138 a_n3166_n47928 0.101866f
C233 VDD.n1139 a_n3166_n47928 0.101866f
C234 VDD.n1140 a_n3166_n47928 0.101866f
C235 VDD.n1141 a_n3166_n47928 0.101866f
C236 VDD.n1142 a_n3166_n47928 0.101866f
C237 VDD.n1143 a_n3166_n47928 0.101866f
C238 VDD.n1144 a_n3166_n47928 0.101866f
C239 VDD.n1145 a_n3166_n47928 0.101866f
C240 VDD.n1146 a_n3166_n47928 0.101866f
C241 VDD.n1147 a_n3166_n47928 0.101866f
C242 VDD.n1148 a_n3166_n47928 0.101866f
C243 VDD.n1149 a_n3166_n47928 0.101866f
C244 VDD.n1150 a_n3166_n47928 0.101866f
C245 VDD.n1151 a_n3166_n47928 0.101866f
C246 VDD.n1152 a_n3166_n47928 0.101866f
C247 VDD.n1153 a_n3166_n47928 0.101866f
C248 VDD.n1154 a_n3166_n47928 0.101866f
C249 VDD.n1155 a_n3166_n47928 0.101866f
C250 VDD.n1156 a_n3166_n47928 0.101866f
C251 VDD.n1157 a_n3166_n47928 0.101866f
C252 VDD.n1158 a_n3166_n47928 0.101866f
C253 VDD.n1159 a_n3166_n47928 0.101866f
C254 VDD.n1160 a_n3166_n47928 0.101866f
C255 VDD.n1161 a_n3166_n47928 0.101866f
C256 VDD.n1162 a_n3166_n47928 0.101866f
C257 VDD.n1163 a_n3166_n47928 0.101866f
C258 VDD.n1164 a_n3166_n47928 0.101866f
C259 VDD.n1165 a_n3166_n47928 0.101866f
C260 VDD.n1166 a_n3166_n47928 0.101866f
C261 VDD.n1167 a_n3166_n47928 0.101866f
C262 VDD.n1168 a_n3166_n47928 0.101866f
C263 VDD.n1169 a_n3166_n47928 0.101866f
C264 VDD.n1170 a_n3166_n47928 0.101866f
C265 VDD.n1171 a_n3166_n47928 0.101866f
C266 VDD.n1172 a_n3166_n47928 0.101866f
C267 VDD.n1173 a_n3166_n47928 0.101866f
C268 VDD.n1174 a_n3166_n47928 0.101866f
C269 VDD.n1175 a_n3166_n47928 0.101866f
C270 VDD.n1176 a_n3166_n47928 0.101866f
C271 VDD.n1177 a_n3166_n47928 0.101866f
C272 VDD.n1178 a_n3166_n47928 0.101866f
C273 VDD.n1179 a_n3166_n47928 0.101866f
C274 VDD.n1180 a_n3166_n47928 0.101866f
C275 VDD.n1181 a_n3166_n47928 0.101866f
C276 VDD.n1182 a_n3166_n47928 0.101866f
C277 VDD.n1183 a_n3166_n47928 0.101866f
C278 VDD.n1184 a_n3166_n47928 0.101866f
C279 VDD.n1185 a_n3166_n47928 0.101866f
C280 VDD.n1186 a_n3166_n47928 0.101866f
C281 VDD.n1187 a_n3166_n47928 0.101866f
C282 VDD.n1188 a_n3166_n47928 0.101866f
C283 VDD.n1189 a_n3166_n47928 0.101866f
C284 VDD.n1190 a_n3166_n47928 0.101866f
C285 VDD.n1191 a_n3166_n47928 0.101866f
C286 VDD.n1192 a_n3166_n47928 0.101866f
C287 VDD.n1193 a_n3166_n47928 0.101866f
C288 VDD.n1196 a_n3166_n47928 0.101866f
C289 VDD.n1197 a_n3166_n47928 0.101866f
C290 VDD.n1198 a_n3166_n47928 0.101866f
C291 VDD.n1199 a_n3166_n47928 0.101866f
C292 VDD.n1200 a_n3166_n47928 0.101866f
C293 VDD.n1201 a_n3166_n47928 0.101866f
C294 VDD.n1202 a_n3166_n47928 0.101866f
C295 VDD.n1203 a_n3166_n47928 0.101866f
C296 VDD.n1204 a_n3166_n47928 0.101866f
C297 VDD.n1205 a_n3166_n47928 0.101866f
C298 VDD.n1206 a_n3166_n47928 0.101866f
C299 VDD.n1207 a_n3166_n47928 0.101866f
C300 VDD.n1208 a_n3166_n47928 0.101866f
C301 VDD.n1209 a_n3166_n47928 0.101866f
C302 VDD.n1210 a_n3166_n47928 0.101866f
C303 VDD.n1211 a_n3166_n47928 0.101866f
C304 VDD.n1212 a_n3166_n47928 0.101866f
C305 VDD.n1213 a_n3166_n47928 0.101866f
C306 VDD.n1214 a_n3166_n47928 0.101866f
C307 VDD.n1215 a_n3166_n47928 0.101866f
C308 VDD.n1216 a_n3166_n47928 0.101866f
C309 VDD.n1217 a_n3166_n47928 0.101866f
C310 VDD.n1218 a_n3166_n47928 0.101866f
C311 VDD.n1219 a_n3166_n47928 0.101866f
C312 VDD.n1220 a_n3166_n47928 0.101866f
C313 VDD.n1221 a_n3166_n47928 0.101866f
C314 VDD.n1222 a_n3166_n47928 0.101866f
C315 VDD.n1223 a_n3166_n47928 0.101866f
C316 VDD.n1224 a_n3166_n47928 0.101866f
C317 VDD.n1225 a_n3166_n47928 0.101866f
C318 VDD.n1226 a_n3166_n47928 0.101866f
C319 VDD.n1227 a_n3166_n47928 0.101866f
C320 VDD.n1228 a_n3166_n47928 0.101866f
C321 VDD.n1229 a_n3166_n47928 0.101866f
C322 VDD.n1230 a_n3166_n47928 0.101866f
C323 VDD.n1231 a_n3166_n47928 0.101866f
C324 VDD.n1232 a_n3166_n47928 0.101866f
C325 VDD.n1233 a_n3166_n47928 0.101866f
C326 VDD.n1234 a_n3166_n47928 0.101866f
C327 VDD.n1235 a_n3166_n47928 0.101866f
C328 VDD.n1236 a_n3166_n47928 0.101866f
C329 VDD.n1237 a_n3166_n47928 0.101866f
C330 VDD.n1238 a_n3166_n47928 0.101866f
C331 VDD.n1239 a_n3166_n47928 0.101866f
C332 VDD.n1240 a_n3166_n47928 0.101866f
C333 VDD.n1241 a_n3166_n47928 0.101866f
C334 VDD.n1242 a_n3166_n47928 0.101866f
C335 VDD.n1243 a_n3166_n47928 0.101866f
C336 VDD.n1244 a_n3166_n47928 0.101866f
C337 VDD.n1245 a_n3166_n47928 0.101866f
C338 VDD.n1246 a_n3166_n47928 0.101866f
C339 VDD.n1247 a_n3166_n47928 0.101866f
C340 VDD.n1248 a_n3166_n47928 0.101866f
C341 VDD.n1249 a_n3166_n47928 0.101866f
C342 VDD.n1250 a_n3166_n47928 0.101866f
C343 VDD.n1251 a_n3166_n47928 0.101866f
C344 VDD.n1252 a_n3166_n47928 0.101866f
C345 VDD.n1253 a_n3166_n47928 0.101866f
C346 VDD.n1254 a_n3166_n47928 0.101866f
C347 VDD.n1255 a_n3166_n47928 0.101866f
C348 VDD.n1256 a_n3166_n47928 0.101866f
C349 VDD.n1257 a_n3166_n47928 0.101866f
C350 VDD.n1260 a_n3166_n47928 0.101866f
C351 VDD.n1261 a_n3166_n47928 0.101866f
C352 VDD.n1262 a_n3166_n47928 0.101866f
C353 VDD.n1263 a_n3166_n47928 0.101866f
C354 VDD.n1264 a_n3166_n47928 0.101866f
C355 VDD.n1265 a_n3166_n47928 0.101866f
C356 VDD.n1266 a_n3166_n47928 0.101866f
C357 VDD.n1267 a_n3166_n47928 0.101866f
C358 VDD.n1268 a_n3166_n47928 0.101866f
C359 VDD.n1269 a_n3166_n47928 0.101866f
C360 VDD.n1270 a_n3166_n47928 0.101866f
C361 VDD.n1271 a_n3166_n47928 0.101866f
C362 VDD.n1272 a_n3166_n47928 0.101866f
C363 VDD.n1273 a_n3166_n47928 0.101866f
C364 VDD.n1274 a_n3166_n47928 0.101866f
C365 VDD.n1275 a_n3166_n47928 0.101866f
C366 VDD.n1276 a_n3166_n47928 0.101866f
C367 VDD.n1277 a_n3166_n47928 0.101866f
C368 VDD.n1278 a_n3166_n47928 0.101866f
C369 VDD.n1279 a_n3166_n47928 0.101866f
C370 VDD.n1280 a_n3166_n47928 0.101866f
C371 VDD.n1281 a_n3166_n47928 0.101866f
C372 VDD.n1282 a_n3166_n47928 0.101866f
C373 VDD.n1283 a_n3166_n47928 0.101866f
C374 VDD.n1284 a_n3166_n47928 0.101866f
C375 VDD.n1285 a_n3166_n47928 0.101866f
C376 VDD.n1286 a_n3166_n47928 0.101866f
C377 VDD.n1287 a_n3166_n47928 0.101866f
C378 VDD.n1288 a_n3166_n47928 0.101866f
C379 VDD.n1289 a_n3166_n47928 0.101866f
C380 VDD.n1290 a_n3166_n47928 0.101866f
C381 VDD.n1291 a_n3166_n47928 0.101866f
C382 VDD.n1292 a_n3166_n47928 0.101866f
C383 VDD.n1293 a_n3166_n47928 0.101866f
C384 VDD.n1294 a_n3166_n47928 0.101866f
C385 VDD.n1295 a_n3166_n47928 0.101866f
C386 VDD.n1296 a_n3166_n47928 0.101866f
C387 VDD.n1297 a_n3166_n47928 0.101866f
C388 VDD.n1298 a_n3166_n47928 0.101866f
C389 VDD.n1299 a_n3166_n47928 0.101866f
C390 VDD.n1300 a_n3166_n47928 0.101866f
C391 VDD.n1301 a_n3166_n47928 0.101866f
C392 VDD.n1302 a_n3166_n47928 0.101866f
C393 VDD.n1303 a_n3166_n47928 0.101866f
C394 VDD.n1304 a_n3166_n47928 0.101866f
C395 VDD.n1305 a_n3166_n47928 0.101866f
C396 VDD.n1306 a_n3166_n47928 0.101866f
C397 VDD.n1307 a_n3166_n47928 0.101866f
C398 VDD.n1308 a_n3166_n47928 0.101866f
C399 VDD.n1309 a_n3166_n47928 0.101866f
C400 VDD.n1310 a_n3166_n47928 0.101866f
C401 VDD.n1311 a_n3166_n47928 0.101866f
C402 VDD.n1312 a_n3166_n47928 0.101866f
C403 VDD.n1313 a_n3166_n47928 0.101866f
C404 VDD.n1314 a_n3166_n47928 0.101866f
C405 VDD.n1315 a_n3166_n47928 0.101866f
C406 VDD.n1316 a_n3166_n47928 0.101866f
C407 VDD.n1317 a_n3166_n47928 0.101866f
C408 VDD.n1318 a_n3166_n47928 0.101866f
C409 VDD.n1319 a_n3166_n47928 0.101866f
C410 VDD.n1320 a_n3166_n47928 0.101866f
C411 VDD.n1321 a_n3166_n47928 0.101866f
C412 VDD.n1322 a_n3166_n47928 0.101866f
C413 VDD.n1323 a_n3166_n47928 0.101866f
C414 VDD.n1324 a_n3166_n47928 0.101866f
C415 VDD.n1325 a_n3166_n47928 0.101866f
C416 VDD.n1326 a_n3166_n47928 0.101866f
C417 VDD.n1327 a_n3166_n47928 0.101866f
C418 VDD.n1328 a_n3166_n47928 0.101866f
C419 VDD.n1329 a_n3166_n47928 0.101866f
C420 VDD.n1330 a_n3166_n47928 0.101866f
C421 VDD.n1331 a_n3166_n47928 0.101866f
C422 VDD.n1332 a_n3166_n47928 0.101866f
C423 VDD.n1333 a_n3166_n47928 0.101866f
C424 VDD.n1334 a_n3166_n47928 0.101866f
C425 VDD.n1335 a_n3166_n47928 0.101866f
C426 VDD.n1336 a_n3166_n47928 0.101866f
C427 VDD.n1337 a_n3166_n47928 0.101866f
C428 VDD.n1338 a_n3166_n47928 0.101866f
C429 VDD.n1339 a_n3166_n47928 0.101866f
C430 VDD.n1340 a_n3166_n47928 0.101866f
C431 VDD.n1341 a_n3166_n47928 0.101866f
C432 VDD.n1342 a_n3166_n47928 0.101866f
C433 VDD.n1343 a_n3166_n47928 0.101866f
C434 VDD.n1344 a_n3166_n47928 0.101866f
C435 VDD.n1345 a_n3166_n47928 0.101866f
C436 VDD.n1346 a_n3166_n47928 0.101866f
C437 VDD.n1347 a_n3166_n47928 0.101866f
C438 VDD.n1348 a_n3166_n47928 0.101866f
C439 VDD.n1349 a_n3166_n47928 0.101866f
C440 VDD.n1350 a_n3166_n47928 0.101866f
C441 VDD.n1351 a_n3166_n47928 0.101866f
C442 VDD.n1352 a_n3166_n47928 0.101866f
C443 VDD.n1353 a_n3166_n47928 0.101866f
C444 VDD.n1354 a_n3166_n47928 0.101866f
C445 VDD.n1355 a_n3166_n47928 0.101866f
C446 VDD.n1356 a_n3166_n47928 0.101866f
C447 VDD.n1357 a_n3166_n47928 0.101866f
C448 VDD.n1358 a_n3166_n47928 0.101866f
C449 VDD.n1359 a_n3166_n47928 0.101866f
C450 VDD.n1360 a_n3166_n47928 0.101866f
C451 VDD.n1361 a_n3166_n47928 0.101866f
C452 VDD.n1362 a_n3166_n47928 0.101866f
C453 VDD.n1363 a_n3166_n47928 0.101866f
C454 VDD.n1364 a_n3166_n47928 0.101866f
C455 VDD.n1365 a_n3166_n47928 0.101866f
C456 VDD.n1366 a_n3166_n47928 0.101866f
C457 VDD.n1367 a_n3166_n47928 0.101866f
C458 VDD.n1368 a_n3166_n47928 0.101866f
C459 VDD.n1369 a_n3166_n47928 0.101866f
C460 VDD.n1370 a_n3166_n47928 0.101866f
C461 VDD.n1371 a_n3166_n47928 0.101866f
C462 VDD.n1372 a_n3166_n47928 0.101866f
C463 VDD.n1373 a_n3166_n47928 0.101866f
C464 VDD.n1374 a_n3166_n47928 0.101866f
C465 VDD.n1375 a_n3166_n47928 0.101866f
C466 VDD.n1376 a_n3166_n47928 0.101866f
C467 VDD.n1377 a_n3166_n47928 0.101866f
C468 VDD.n1378 a_n3166_n47928 0.101866f
C469 VDD.n1379 a_n3166_n47928 0.101866f
C470 VDD.n1380 a_n3166_n47928 0.101866f
C471 VDD.n1381 a_n3166_n47928 0.101866f
C472 VDD.n1382 a_n3166_n47928 0.101866f
C473 VDD.n1383 a_n3166_n47928 0.101866f
C474 VDD.n1384 a_n3166_n47928 0.101866f
C475 VDD.n1385 a_n3166_n47928 0.101866f
C476 VDD.n1386 a_n3166_n47928 0.101866f
C477 VDD.n1387 a_n3166_n47928 0.101866f
C478 VDD.n1388 a_n3166_n47928 0.101866f
C479 VDD.n1389 a_n3166_n47928 0.101866f
C480 VDD.n1390 a_n3166_n47928 0.101866f
C481 VDD.n1391 a_n3166_n47928 0.101866f
C482 VDD.n1392 a_n3166_n47928 0.101866f
C483 VDD.n1393 a_n3166_n47928 0.101866f
C484 VDD.n1394 a_n3166_n47928 0.101866f
C485 VDD.n1395 a_n3166_n47928 0.101866f
C486 VDD.n1396 a_n3166_n47928 0.101866f
C487 VDD.n1397 a_n3166_n47928 0.101866f
C488 VDD.n1398 a_n3166_n47928 0.101866f
C489 VDD.n1399 a_n3166_n47928 0.101866f
C490 VDD.n1400 a_n3166_n47928 0.101866f
C491 VDD.n1401 a_n3166_n47928 0.101866f
C492 VDD.n1402 a_n3166_n47928 0.101866f
C493 VDD.n1403 a_n3166_n47928 0.101866f
C494 VDD.n1404 a_n3166_n47928 0.101866f
C495 VDD.n1405 a_n3166_n47928 0.101866f
C496 VDD.n1406 a_n3166_n47928 0.101866f
C497 VDD.n1407 a_n3166_n47928 0.101866f
C498 VDD.n1408 a_n3166_n47928 0.101866f
C499 VDD.n1409 a_n3166_n47928 0.101866f
C500 VDD.n1410 a_n3166_n47928 0.101866f
C501 VDD.n1411 a_n3166_n47928 0.101866f
C502 VDD.n1412 a_n3166_n47928 0.101866f
C503 VDD.n1413 a_n3166_n47928 0.101866f
C504 VDD.n1414 a_n3166_n47928 0.101866f
C505 VDD.n1415 a_n3166_n47928 0.101866f
C506 VDD.n1416 a_n3166_n47928 0.101866f
C507 VDD.n1480 a_n3166_n47928 0.103509f
C508 VDD.n1544 a_n3166_n47928 0.101866f
C509 VDD.n1607 a_n3166_n47928 0.101866f
C510 VDD.n1671 a_n3166_n47928 0.101866f
C511 VDD.n1672 a_n3166_n47928 0.101866f
C512 VDD.n1673 a_n3166_n47928 0.105997f
C513 VDD.n1674 a_n3166_n47928 0.103509f
C514 VDD.n1675 a_n3166_n47928 0.101866f
C515 VDD.n1676 a_n3166_n47928 0.103509f
C516 VDD.n1677 a_n3166_n47928 0.105997f
C517 VDD.n1678 a_n3166_n47928 0.107553f
C518 VDD.n1679 a_n3166_n47928 0.101866f
C519 VDD.n1680 a_n3166_n47928 0.101866f
C520 VDD.n1681 a_n3166_n47928 0.101866f
C521 VDD.n1682 a_n3166_n47928 0.101866f
C522 VDD.n1683 a_n3166_n47928 0.101866f
C523 VDD.n1684 a_n3166_n47928 0.101866f
C524 VDD.n1685 a_n3166_n47928 0.101866f
C525 VDD.n1686 a_n3166_n47928 0.101866f
C526 VDD.n1687 a_n3166_n47928 0.101866f
C527 VDD.n1688 a_n3166_n47928 0.101866f
C528 VDD.n1689 a_n3166_n47928 0.101866f
C529 VDD.n1690 a_n3166_n47928 0.101866f
C530 VDD.n1691 a_n3166_n47928 0.101866f
C531 VDD.n1692 a_n3166_n47928 0.101866f
C532 VDD.n1693 a_n3166_n47928 0.101866f
C533 VDD.n1694 a_n3166_n47928 0.101866f
C534 VDD.n1695 a_n3166_n47928 0.101866f
C535 VDD.n1696 a_n3166_n47928 0.101866f
C536 VDD.n1697 a_n3166_n47928 0.101866f
C537 VDD.n1698 a_n3166_n47928 0.101866f
C538 VDD.n1699 a_n3166_n47928 0.101866f
C539 VDD.n1700 a_n3166_n47928 0.101866f
C540 VDD.n1701 a_n3166_n47928 0.101866f
C541 VDD.n1702 a_n3166_n47928 0.101866f
C542 VDD.n1703 a_n3166_n47928 0.101866f
C543 VDD.n1704 a_n3166_n47928 0.101866f
C544 VDD.n1705 a_n3166_n47928 0.101866f
C545 VDD.n1706 a_n3166_n47928 0.101866f
C546 VDD.n1707 a_n3166_n47928 0.101866f
C547 VDD.n1708 a_n3166_n47928 0.101866f
C548 VDD.n1709 a_n3166_n47928 0.101866f
C549 VDD.n1710 a_n3166_n47928 0.101866f
C550 VDD.n1711 a_n3166_n47928 0.101866f
C551 VDD.n1712 a_n3166_n47928 0.101866f
C552 VDD.n1713 a_n3166_n47928 0.101866f
C553 VDD.n1714 a_n3166_n47928 0.101866f
C554 VDD.n1715 a_n3166_n47928 0.101866f
C555 VDD.n1716 a_n3166_n47928 0.101866f
C556 VDD.n1717 a_n3166_n47928 0.101866f
C557 VDD.n1718 a_n3166_n47928 0.101866f
C558 VDD.n1719 a_n3166_n47928 0.101866f
C559 VDD.n1720 a_n3166_n47928 0.101866f
C560 VDD.n1721 a_n3166_n47928 0.101866f
C561 VDD.n1722 a_n3166_n47928 0.101866f
C562 VDD.n1723 a_n3166_n47928 0.101866f
C563 VDD.n1724 a_n3166_n47928 0.101866f
C564 VDD.n1725 a_n3166_n47928 0.101866f
C565 VDD.n1726 a_n3166_n47928 0.101866f
C566 VDD.n1727 a_n3166_n47928 0.101866f
C567 VDD.n1728 a_n3166_n47928 0.101866f
C568 VDD.n1729 a_n3166_n47928 0.101866f
C569 VDD.n1730 a_n3166_n47928 0.101866f
C570 VDD.n1731 a_n3166_n47928 0.101866f
C571 VDD.n1732 a_n3166_n47928 0.101866f
C572 VDD.n1733 a_n3166_n47928 0.101866f
C573 VDD.n1734 a_n3166_n47928 0.101866f
C574 VDD.n1735 a_n3166_n47928 0.101866f
C575 VDD.n1736 a_n3166_n47928 0.101866f
C576 VDD.n1737 a_n3166_n47928 0.101866f
C577 VDD.n1738 a_n3166_n47928 0.101866f
C578 VDD.n1739 a_n3166_n47928 0.101866f
C579 VDD.n1740 a_n3166_n47928 0.101866f
C580 VDD.n1741 a_n3166_n47928 0.101866f
C581 VDD.n1742 a_n3166_n47928 0.101866f
C582 VDD.n1743 a_n3166_n47928 0.101866f
C583 VDD.n1744 a_n3166_n47928 0.059148f
C584 VDD.n1745 a_n3166_n47928 0.101866f
C585 VDD.n1746 a_n3166_n47928 0.101866f
C586 VDD.n1747 a_n3166_n47928 0.093651f
C587 VDD.n1748 a_n3166_n47928 0.101866f
C588 VDD.n1749 a_n3166_n47928 0.101866f
C589 VDD.n1750 a_n3166_n47928 0.101866f
C590 VDD.n1751 a_n3166_n47928 0.101866f
C591 VDD.n1752 a_n3166_n47928 0.101866f
C592 VDD.n1753 a_n3166_n47928 0.101866f
C593 VDD.n1754 a_n3166_n47928 0.101866f
C594 VDD.n1755 a_n3166_n47928 0.101866f
C595 VDD.n1756 a_n3166_n47928 0.101866f
C596 VDD.n1757 a_n3166_n47928 0.101866f
C597 VDD.n1758 a_n3166_n47928 0.101866f
C598 VDD.n1759 a_n3166_n47928 0.101866f
C599 VDD.n1760 a_n3166_n47928 0.101866f
C600 VDD.n1761 a_n3166_n47928 0.101866f
C601 VDD.n1762 a_n3166_n47928 0.101866f
C602 VDD.n1763 a_n3166_n47928 0.101866f
C603 VDD.n1764 a_n3166_n47928 0.101866f
C604 VDD.n1765 a_n3166_n47928 0.101866f
C605 VDD.n1766 a_n3166_n47928 0.101866f
C606 VDD.n1767 a_n3166_n47928 0.101866f
C607 VDD.n1768 a_n3166_n47928 0.101866f
C608 VDD.n1769 a_n3166_n47928 0.101866f
C609 VDD.n1770 a_n3166_n47928 0.101866f
C610 VDD.n1771 a_n3166_n47928 0.101866f
C611 VDD.n1772 a_n3166_n47928 0.101866f
C612 VDD.n1773 a_n3166_n47928 0.101866f
C613 VDD.n1774 a_n3166_n47928 0.101866f
C614 VDD.n1775 a_n3166_n47928 0.101866f
C615 VDD.n1776 a_n3166_n47928 0.101866f
C616 VDD.n1777 a_n3166_n47928 0.101866f
C617 VDD.n1778 a_n3166_n47928 0.101866f
C618 VDD.n1779 a_n3166_n47928 0.101866f
C619 VDD.n1780 a_n3166_n47928 0.101866f
C620 VDD.n1781 a_n3166_n47928 0.101866f
C621 VDD.n1782 a_n3166_n47928 0.101866f
C622 VDD.n1783 a_n3166_n47928 0.101866f
C623 VDD.n1784 a_n3166_n47928 0.101866f
C624 VDD.n1785 a_n3166_n47928 0.101866f
C625 VDD.n1786 a_n3166_n47928 0.101866f
C626 VDD.n1787 a_n3166_n47928 0.101866f
C627 VDD.n1788 a_n3166_n47928 0.101866f
C628 VDD.n1789 a_n3166_n47928 0.101866f
C629 VDD.n1790 a_n3166_n47928 0.101866f
C630 VDD.n1791 a_n3166_n47928 0.101866f
C631 VDD.n1792 a_n3166_n47928 0.101866f
C632 VDD.n1793 a_n3166_n47928 0.101866f
C633 VDD.n1794 a_n3166_n47928 0.101866f
C634 VDD.n1795 a_n3166_n47928 0.101866f
C635 VDD.n1796 a_n3166_n47928 0.101866f
C636 VDD.n1797 a_n3166_n47928 0.101866f
C637 VDD.n1798 a_n3166_n47928 0.101866f
C638 VDD.n1799 a_n3166_n47928 0.101866f
C639 VDD.n1800 a_n3166_n47928 0.101866f
C640 VDD.n1801 a_n3166_n47928 0.101866f
C641 VDD.n1802 a_n3166_n47928 0.101866f
C642 VDD.n1803 a_n3166_n47928 0.101866f
C643 VDD.n1804 a_n3166_n47928 0.101866f
C644 VDD.n1805 a_n3166_n47928 0.101866f
C645 VDD.n1806 a_n3166_n47928 0.101866f
C646 VDD.n1807 a_n3166_n47928 0.101866f
C647 VDD.n1808 a_n3166_n47928 0.101866f
C648 VDD.n1809 a_n3166_n47928 0.101866f
C649 VDD.n1810 a_n3166_n47928 0.101866f
C650 VDD.n1811 a_n3166_n47928 0.101866f
C651 VDD.n1812 a_n3166_n47928 0.101866f
C652 VDD.n1813 a_n3166_n47928 0.101866f
C653 VDD.n1814 a_n3166_n47928 0.101866f
C654 VDD.n1815 a_n3166_n47928 0.101866f
C655 VDD.n1816 a_n3166_n47928 0.101866f
C656 VDD.n1817 a_n3166_n47928 0.101866f
C657 VDD.n1818 a_n3166_n47928 0.101866f
C658 VDD.n1819 a_n3166_n47928 0.101866f
C659 VDD.n1820 a_n3166_n47928 0.101866f
C660 VDD.n1821 a_n3166_n47928 0.101866f
C661 VDD.n1822 a_n3166_n47928 0.101866f
C662 VDD.n1823 a_n3166_n47928 0.101866f
C663 VDD.n1824 a_n3166_n47928 0.101866f
C664 VDD.n1825 a_n3166_n47928 0.101866f
C665 VDD.n1826 a_n3166_n47928 0.101866f
C666 VDD.n1827 a_n3166_n47928 0.101866f
C667 VDD.n1828 a_n3166_n47928 0.101866f
C668 VDD.n1829 a_n3166_n47928 0.101866f
C669 VDD.n1830 a_n3166_n47928 0.101866f
C670 VDD.n1831 a_n3166_n47928 0.101866f
C671 VDD.n1832 a_n3166_n47928 0.101866f
C672 VDD.n1833 a_n3166_n47928 0.101866f
C673 VDD.n1834 a_n3166_n47928 0.101866f
C674 VDD.n1835 a_n3166_n47928 0.101866f
C675 VDD.n1836 a_n3166_n47928 0.101866f
C676 VDD.n1837 a_n3166_n47928 0.101866f
C677 VDD.n1838 a_n3166_n47928 0.101866f
C678 VDD.n1839 a_n3166_n47928 0.101866f
C679 VDD.n1840 a_n3166_n47928 0.101866f
C680 VDD.n1841 a_n3166_n47928 0.101866f
C681 VDD.n1842 a_n3166_n47928 0.101866f
C682 VDD.n1843 a_n3166_n47928 0.101866f
C683 VDD.n1844 a_n3166_n47928 0.101866f
C684 VDD.n1845 a_n3166_n47928 0.101866f
C685 VDD.n1846 a_n3166_n47928 0.101866f
C686 VDD.n1847 a_n3166_n47928 0.101866f
C687 VDD.n1848 a_n3166_n47928 0.101866f
C688 VDD.n1849 a_n3166_n47928 0.101866f
C689 VDD.n1850 a_n3166_n47928 0.101866f
C690 VDD.n1851 a_n3166_n47928 0.101866f
C691 VDD.n1852 a_n3166_n47928 0.101866f
C692 VDD.n1853 a_n3166_n47928 0.101866f
C693 VDD.n1854 a_n3166_n47928 0.101866f
C694 VDD.n1855 a_n3166_n47928 0.101866f
C695 VDD.n1856 a_n3166_n47928 0.101866f
C696 VDD.n1857 a_n3166_n47928 0.101866f
C697 VDD.n1858 a_n3166_n47928 0.101866f
C698 VDD.n1859 a_n3166_n47928 0.101866f
C699 VDD.n1860 a_n3166_n47928 0.101866f
C700 VDD.n1861 a_n3166_n47928 0.101866f
C701 VDD.n1862 a_n3166_n47928 0.101866f
C702 VDD.n1863 a_n3166_n47928 0.101866f
C703 VDD.n1864 a_n3166_n47928 0.101866f
C704 VDD.n1865 a_n3166_n47928 0.101866f
C705 VDD.n1866 a_n3166_n47928 0.101866f
C706 VDD.n1867 a_n3166_n47928 0.300709f
C707 IB.n18 a_n3166_n47928 0.016419f
C708 IB.n19 a_n3166_n47928 0.016419f
C709 IB.n22 a_n3166_n47928 0.016419f
C710 IB.n23 a_n3166_n47928 0.016419f
C711 IB.n24 a_n3166_n47928 0.015808f
C712 IB.n25 a_n3166_n47928 0.013916f
C713 IB.n28 a_n3166_n47928 0.273605f
C714 a_2044_n43060.n0 a_n3166_n47928 1.80114f
C715 a_2044_n43060.t10 a_n3166_n47928 0.034355f
C716 a_2044_n43060.t22 a_n3166_n47928 0.18159f
C717 a_2044_n43060.t1 a_n3166_n47928 0.280391f
C718 a_2044_n43060.t0 a_n3166_n47928 0.163334f
C719 a_2044_n43060.t4 a_n3166_n47928 0.271534f
C720 a_2044_n43060.n1 a_n3166_n47928 0.762311f
C721 a_2044_n43060.t16 a_n3166_n47928 0.034355f
C722 a_2044_n43060.t14 a_n3166_n47928 0.034355f
C723 a_2044_n43060.n2 a_n3166_n47928 0.170659f
C724 a_2044_n43060.n3 a_n3166_n47928 0.309174f
C725 a_2044_n43060.t8 a_n3166_n47928 0.034355f
C726 a_2044_n43060.t3 a_n3166_n47928 0.034355f
C727 a_2044_n43060.n4 a_n3166_n47928 0.170659f
C728 a_2044_n43060.n5 a_n3166_n47928 0.293318f
C729 a_2044_n43060.t12 a_n3166_n47928 0.034355f
C730 a_2044_n43060.t7 a_n3166_n47928 0.034355f
C731 a_2044_n43060.n6 a_n3166_n47928 0.170659f
C732 a_2044_n43060.n7 a_n3166_n47928 0.293318f
C733 a_2044_n43060.t20 a_n3166_n47928 0.034355f
C734 a_2044_n43060.t15 a_n3166_n47928 0.034355f
C735 a_2044_n43060.n8 a_n3166_n47928 0.170659f
C736 a_2044_n43060.n9 a_n3166_n47928 0.293318f
C737 a_2044_n43060.t11 a_n3166_n47928 0.034355f
C738 a_2044_n43060.t19 a_n3166_n47928 0.034355f
C739 a_2044_n43060.n10 a_n3166_n47928 0.170659f
C740 a_2044_n43060.n11 a_n3166_n47928 0.293318f
C741 a_2044_n43060.t5 a_n3166_n47928 0.276199f
C742 a_2044_n43060.t17 a_n3166_n47928 0.034355f
C743 a_2044_n43060.t13 a_n3166_n47928 0.034355f
C744 a_2044_n43060.n12 a_n3166_n47928 0.170659f
C745 a_2044_n43060.n13 a_n3166_n47928 0.546786f
C746 a_2044_n43060.t6 a_n3166_n47928 0.034355f
C747 a_2044_n43060.t9 a_n3166_n47928 0.034355f
C748 a_2044_n43060.n14 a_n3166_n47928 0.170659f
C749 a_2044_n43060.n15 a_n3166_n47928 0.293318f
C750 a_2044_n43060.t2 a_n3166_n47928 0.034355f
C751 a_2044_n43060.t18 a_n3166_n47928 0.034355f
C752 a_2044_n43060.n16 a_n3166_n47928 0.170659f
C753 a_2044_n43060.n17 a_n3166_n47928 0.293318f
C754 a_2044_n43060.n18 a_n3166_n47928 0.293318f
C755 a_2044_n43060.n19 a_n3166_n47928 0.170659f
C756 a_2044_n43060.t21 a_n3166_n47928 0.034355f
C757 VINN.n0 a_n3166_n47928 0.0274f
C758 VINN.n1 a_n3166_n47928 0.026615f
C759 VINN.n85 a_n3166_n47928 0.032685f
C760 VINN.n86 a_n3166_n47928 0.059161f
C761 VINN.n87 a_n3166_n47928 0.026615f
C762 VINN.n88 a_n3166_n47928 0.026615f
C763 VINN.n89 a_n3166_n47928 0.026615f
C764 VINN.n90 a_n3166_n47928 0.026615f
C765 VINN.n91 a_n3166_n47928 0.026615f
C766 VINN.n92 a_n3166_n47928 0.026615f
C767 VINN.n93 a_n3166_n47928 0.026615f
C768 VINN.n94 a_n3166_n47928 0.026615f
C769 VINN.n95 a_n3166_n47928 0.026615f
C770 VINN.n96 a_n3166_n47928 0.026615f
C771 VINN.n97 a_n3166_n47928 0.026615f
C772 VINN.n98 a_n3166_n47928 0.026615f
C773 VINN.n99 a_n3166_n47928 0.026615f
C774 VINN.n100 a_n3166_n47928 0.026615f
C775 VINN.n101 a_n3166_n47928 0.026615f
C776 VINN.n102 a_n3166_n47928 0.026615f
C777 VINN.n103 a_n3166_n47928 0.026615f
C778 VINN.n104 a_n3166_n47928 0.026615f
C779 VINN.n105 a_n3166_n47928 0.026615f
C780 VINN.n106 a_n3166_n47928 0.026615f
C781 VINN.n107 a_n3166_n47928 0.026615f
C782 VINN.n108 a_n3166_n47928 0.026615f
C783 VINN.n109 a_n3166_n47928 0.026615f
C784 VINN.n110 a_n3166_n47928 0.026615f
C785 VINN.n111 a_n3166_n47928 0.026615f
C786 VINN.n112 a_n3166_n47928 0.026615f
C787 VINN.n113 a_n3166_n47928 0.026615f
C788 VINN.n114 a_n3166_n47928 0.026615f
C789 VINN.n115 a_n3166_n47928 0.026615f
C790 VINN.n116 a_n3166_n47928 0.026615f
C791 VINN.n117 a_n3166_n47928 0.026615f
C792 VINN.n118 a_n3166_n47928 0.026615f
C793 VINN.n119 a_n3166_n47928 0.026615f
C794 VINN.n120 a_n3166_n47928 0.026615f
C795 VINN.n121 a_n3166_n47928 0.026615f
C796 VINN.n122 a_n3166_n47928 0.026615f
C797 VINN.n123 a_n3166_n47928 0.026615f
C798 VINN.n124 a_n3166_n47928 0.026615f
C799 VINN.n125 a_n3166_n47928 0.026615f
C800 VINN.n126 a_n3166_n47928 0.026615f
C801 VINN.n127 a_n3166_n47928 0.026615f
C802 VINN.n128 a_n3166_n47928 0.026615f
C803 VINN.n129 a_n3166_n47928 0.026615f
C804 VINN.n130 a_n3166_n47928 0.026615f
C805 VINN.n131 a_n3166_n47928 0.026615f
C806 VINN.n132 a_n3166_n47928 0.026615f
C807 VINN.n133 a_n3166_n47928 0.026615f
C808 VINN.n134 a_n3166_n47928 0.026615f
C809 VINN.n135 a_n3166_n47928 0.026615f
C810 VINN.n136 a_n3166_n47928 0.026615f
C811 VINN.n137 a_n3166_n47928 0.026615f
C812 VINN.n138 a_n3166_n47928 0.026615f
C813 VINN.n139 a_n3166_n47928 0.026615f
C814 VINN.n140 a_n3166_n47928 0.026615f
C815 VINN.n141 a_n3166_n47928 0.026615f
C816 VINN.n142 a_n3166_n47928 0.026615f
C817 VINN.n143 a_n3166_n47928 0.026615f
C818 VINN.n144 a_n3166_n47928 0.026615f
C819 VINN.n145 a_n3166_n47928 0.026615f
C820 VINN.n146 a_n3166_n47928 0.026615f
C821 VINN.n147 a_n3166_n47928 0.026615f
C822 VINN.n148 a_n3166_n47928 0.026615f
C823 VINN.n149 a_n3166_n47928 0.026615f
C824 VINN.n151 a_n3166_n47928 0.026615f
C825 VINN.n152 a_n3166_n47928 0.026615f
C826 VINN.n153 a_n3166_n47928 0.026615f
C827 VINN.n154 a_n3166_n47928 0.026615f
C828 VINN.n155 a_n3166_n47928 0.026615f
C829 VINN.n156 a_n3166_n47928 0.026615f
C830 VINN.n157 a_n3166_n47928 0.026615f
C831 VINN.n158 a_n3166_n47928 0.026615f
C832 VINN.n159 a_n3166_n47928 0.026615f
C833 VINN.n160 a_n3166_n47928 0.026615f
C834 VINN.n161 a_n3166_n47928 0.026615f
C835 VINN.n162 a_n3166_n47928 0.026615f
C836 VINN.n163 a_n3166_n47928 0.026615f
C837 VINN.n164 a_n3166_n47928 0.026615f
C838 VINN.n165 a_n3166_n47928 0.026615f
C839 VINN.n166 a_n3166_n47928 0.026615f
C840 VINN.n167 a_n3166_n47928 0.026615f
C841 VINN.n168 a_n3166_n47928 0.026615f
C842 VINN.n169 a_n3166_n47928 0.026615f
C843 VINN.n170 a_n3166_n47928 0.026615f
C844 VINN.n171 a_n3166_n47928 0.026615f
C845 VINN.n172 a_n3166_n47928 0.026615f
C846 VINN.n173 a_n3166_n47928 0.026615f
C847 VINN.n174 a_n3166_n47928 0.026615f
C848 VINN.n175 a_n3166_n47928 0.026615f
C849 VINN.n176 a_n3166_n47928 0.026615f
C850 VINN.n177 a_n3166_n47928 0.026615f
C851 VINN.n178 a_n3166_n47928 0.026615f
C852 VINN.n179 a_n3166_n47928 0.026615f
C853 VINN.n180 a_n3166_n47928 0.026615f
C854 VINN.n181 a_n3166_n47928 0.026615f
C855 VINN.n182 a_n3166_n47928 0.026615f
C856 VINN.n183 a_n3166_n47928 0.026615f
C857 VINN.n184 a_n3166_n47928 0.026615f
C858 VINN.n185 a_n3166_n47928 0.026615f
C859 VINN.n186 a_n3166_n47928 0.026615f
C860 VINN.n187 a_n3166_n47928 0.026615f
C861 VINN.n188 a_n3166_n47928 0.026615f
C862 VINN.n189 a_n3166_n47928 0.026615f
C863 VINN.n190 a_n3166_n47928 0.026615f
C864 VINN.n191 a_n3166_n47928 0.026615f
C865 VINN.n192 a_n3166_n47928 0.026615f
C866 VINN.n193 a_n3166_n47928 0.026615f
C867 VINN.n194 a_n3166_n47928 0.026615f
C868 VINN.n195 a_n3166_n47928 0.026615f
C869 VINN.n196 a_n3166_n47928 0.026615f
C870 VINN.n197 a_n3166_n47928 0.026615f
C871 VINN.n198 a_n3166_n47928 0.026615f
C872 VINN.n199 a_n3166_n47928 0.026615f
C873 VINN.n200 a_n3166_n47928 0.026615f
C874 VINN.n201 a_n3166_n47928 0.026615f
C875 VINN.n202 a_n3166_n47928 0.026615f
C876 VINN.n203 a_n3166_n47928 0.026615f
C877 VINN.n204 a_n3166_n47928 0.026615f
C878 VINN.n205 a_n3166_n47928 0.026615f
C879 VINN.n206 a_n3166_n47928 0.026615f
C880 VINN.n207 a_n3166_n47928 0.026615f
C881 VINN.n208 a_n3166_n47928 0.026615f
C882 VINN.n209 a_n3166_n47928 0.026615f
C883 VINN.n210 a_n3166_n47928 0.026615f
C884 VINN.n211 a_n3166_n47928 0.026615f
C885 VINN.n212 a_n3166_n47928 0.026615f
C886 VINN.n213 a_n3166_n47928 0.026615f
C887 VINN.n215 a_n3166_n47928 0.026615f
C888 VINN.n216 a_n3166_n47928 0.026615f
C889 VINN.n217 a_n3166_n47928 0.026615f
C890 VINN.n218 a_n3166_n47928 0.026615f
C891 VINN.n219 a_n3166_n47928 0.026615f
C892 VINN.n220 a_n3166_n47928 0.026615f
C893 VINN.n221 a_n3166_n47928 0.026615f
C894 VINN.n222 a_n3166_n47928 0.026615f
C895 VINN.n223 a_n3166_n47928 0.026615f
C896 VINN.n224 a_n3166_n47928 0.026615f
C897 VINN.n225 a_n3166_n47928 0.026615f
C898 VINN.n226 a_n3166_n47928 0.026615f
C899 VINN.n227 a_n3166_n47928 0.026615f
C900 VINN.n228 a_n3166_n47928 0.026615f
C901 VINN.n229 a_n3166_n47928 0.026615f
C902 VINN.n230 a_n3166_n47928 0.026615f
C903 VINN.n231 a_n3166_n47928 0.026615f
C904 VINN.n232 a_n3166_n47928 0.026615f
C905 VINN.n233 a_n3166_n47928 0.026615f
C906 VINN.n234 a_n3166_n47928 0.026615f
C907 VINN.n235 a_n3166_n47928 0.026615f
C908 VINN.n236 a_n3166_n47928 0.026615f
C909 VINN.n237 a_n3166_n47928 0.026615f
C910 VINN.n238 a_n3166_n47928 0.026615f
C911 VINN.n239 a_n3166_n47928 0.026615f
C912 VINN.n240 a_n3166_n47928 0.026615f
C913 VINN.n241 a_n3166_n47928 0.026615f
C914 VINN.n242 a_n3166_n47928 0.026615f
C915 VINN.n243 a_n3166_n47928 0.026615f
C916 VINN.n244 a_n3166_n47928 0.026615f
C917 VINN.n245 a_n3166_n47928 0.026615f
C918 VINN.n246 a_n3166_n47928 0.026615f
C919 VINN.n247 a_n3166_n47928 0.026615f
C920 VINN.n248 a_n3166_n47928 0.026615f
C921 VINN.n249 a_n3166_n47928 0.026615f
C922 VINN.n250 a_n3166_n47928 0.026615f
C923 VINN.n251 a_n3166_n47928 0.026615f
C924 VINN.n252 a_n3166_n47928 0.026615f
C925 VINN.n253 a_n3166_n47928 0.026615f
C926 VINN.n254 a_n3166_n47928 0.026615f
C927 VINN.n255 a_n3166_n47928 0.026615f
C928 VINN.n256 a_n3166_n47928 0.026615f
C929 VINN.n257 a_n3166_n47928 0.026615f
C930 VINN.n258 a_n3166_n47928 0.026615f
C931 VINN.n259 a_n3166_n47928 0.026615f
C932 VINN.n260 a_n3166_n47928 0.026615f
C933 VINN.n261 a_n3166_n47928 0.026615f
C934 VINN.n262 a_n3166_n47928 0.026615f
C935 VINN.n263 a_n3166_n47928 0.026615f
C936 VINN.n264 a_n3166_n47928 0.026615f
C937 VINN.n265 a_n3166_n47928 0.026615f
C938 VINN.n266 a_n3166_n47928 0.026615f
C939 VINN.n267 a_n3166_n47928 0.026615f
C940 VINN.n268 a_n3166_n47928 0.026615f
C941 VINN.n269 a_n3166_n47928 0.026615f
C942 VINN.n270 a_n3166_n47928 0.026615f
C943 VINN.n271 a_n3166_n47928 0.026615f
C944 VINN.n272 a_n3166_n47928 0.026615f
C945 VINN.n273 a_n3166_n47928 0.026615f
C946 VINN.n274 a_n3166_n47928 0.026615f
C947 VINN.n275 a_n3166_n47928 0.026615f
C948 VINN.n276 a_n3166_n47928 0.026615f
C949 VINN.n278 a_n3166_n47928 0.0274f
C950 VINN.n280 a_n3166_n47928 0.026615f
C951 VINN.n282 a_n3166_n47928 0.026615f
C952 VINN.n284 a_n3166_n47928 0.026615f
C953 VINN.n286 a_n3166_n47928 0.026615f
C954 VINN.n288 a_n3166_n47928 0.026615f
C955 VINN.n290 a_n3166_n47928 0.026615f
C956 VINN.n292 a_n3166_n47928 0.026615f
C957 VINN.n294 a_n3166_n47928 0.026615f
C958 VINN.n296 a_n3166_n47928 0.026615f
C959 VINN.n298 a_n3166_n47928 0.026615f
C960 VINN.n300 a_n3166_n47928 0.026615f
C961 VINN.n302 a_n3166_n47928 0.026615f
C962 VINN.n304 a_n3166_n47928 0.026615f
C963 VINN.n306 a_n3166_n47928 0.026615f
C964 VINN.n308 a_n3166_n47928 0.026615f
C965 VINN.n310 a_n3166_n47928 0.026615f
C966 VINN.n312 a_n3166_n47928 0.026615f
C967 VINN.n314 a_n3166_n47928 0.026615f
C968 VINN.n316 a_n3166_n47928 0.026615f
C969 VINN.n318 a_n3166_n47928 0.026615f
C970 VINN.n320 a_n3166_n47928 0.026615f
C971 VINN.n322 a_n3166_n47928 0.026615f
C972 VINN.n324 a_n3166_n47928 0.026615f
C973 VINN.n326 a_n3166_n47928 0.026615f
C974 VINN.n328 a_n3166_n47928 0.026615f
C975 VINN.n330 a_n3166_n47928 0.026615f
C976 VINN.n332 a_n3166_n47928 0.026615f
C977 VINN.n334 a_n3166_n47928 0.026615f
C978 VINN.n336 a_n3166_n47928 0.026615f
C979 VINN.n338 a_n3166_n47928 0.026615f
C980 VINN.n340 a_n3166_n47928 0.026615f
C981 VINN.n342 a_n3166_n47928 0.026615f
C982 VINN.n344 a_n3166_n47928 0.026615f
C983 VINN.n346 a_n3166_n47928 0.026615f
C984 VINN.n348 a_n3166_n47928 0.026615f
C985 VINN.n350 a_n3166_n47928 0.026615f
C986 VINN.n352 a_n3166_n47928 0.026615f
C987 VINN.n354 a_n3166_n47928 0.026615f
C988 VINN.n356 a_n3166_n47928 0.026615f
C989 VINN.n358 a_n3166_n47928 0.026615f
C990 VINN.n360 a_n3166_n47928 0.026615f
C991 VINN.n362 a_n3166_n47928 0.026615f
C992 VINN.n364 a_n3166_n47928 0.026615f
C993 VINN.n366 a_n3166_n47928 0.026615f
C994 VINN.n368 a_n3166_n47928 0.026615f
C995 VINN.n370 a_n3166_n47928 0.026615f
C996 VINN.n372 a_n3166_n47928 0.026615f
C997 VINN.n374 a_n3166_n47928 0.026615f
C998 VINN.n376 a_n3166_n47928 0.026615f
C999 VINN.n378 a_n3166_n47928 0.026615f
C1000 VINN.n380 a_n3166_n47928 0.026615f
C1001 VINN.n382 a_n3166_n47928 0.026615f
C1002 VINN.n384 a_n3166_n47928 0.026615f
C1003 VINN.n386 a_n3166_n47928 0.026615f
C1004 VINN.n388 a_n3166_n47928 0.026615f
C1005 VINN.n390 a_n3166_n47928 0.026615f
C1006 VINN.n392 a_n3166_n47928 0.026615f
C1007 VINN.n394 a_n3166_n47928 0.026615f
C1008 VINN.n396 a_n3166_n47928 0.026615f
C1009 VINN.n398 a_n3166_n47928 0.026615f
C1010 VINN.n400 a_n3166_n47928 0.026615f
C1011 VINN.n463 a_n3166_n47928 0.027044f
C1012 VINN.n528 a_n3166_n47928 0.026615f
C1013 VINN.n529 a_n3166_n47928 0.026615f
C1014 VINN.n530 a_n3166_n47928 0.053303f
C1015 VINN.n531 a_n3166_n47928 0.026615f
C1016 VINN.n532 a_n3166_n47928 0.026615f
C1017 VINN.n533 a_n3166_n47928 0.026615f
C1018 VINN.n534 a_n3166_n47928 0.026615f
C1019 VINN.n535 a_n3166_n47928 0.026615f
C1020 VINN.n536 a_n3166_n47928 0.026615f
C1021 VINN.n537 a_n3166_n47928 0.026615f
C1022 VINN.n538 a_n3166_n47928 0.026615f
C1023 VINN.n539 a_n3166_n47928 0.026615f
C1024 VINN.n540 a_n3166_n47928 0.026615f
C1025 VINN.n541 a_n3166_n47928 0.026615f
C1026 VINN.n542 a_n3166_n47928 0.026615f
C1027 VINN.n543 a_n3166_n47928 0.026615f
C1028 VINN.n544 a_n3166_n47928 0.026615f
C1029 VINN.n545 a_n3166_n47928 0.026615f
C1030 VINN.n546 a_n3166_n47928 0.026615f
C1031 VINN.n547 a_n3166_n47928 0.026615f
C1032 VINN.n548 a_n3166_n47928 0.026615f
C1033 VINN.n549 a_n3166_n47928 0.026615f
C1034 VINN.n550 a_n3166_n47928 0.026615f
C1035 VINN.n551 a_n3166_n47928 0.026615f
C1036 VINN.n552 a_n3166_n47928 0.026615f
C1037 VINN.n553 a_n3166_n47928 0.026615f
C1038 VINN.n554 a_n3166_n47928 0.026615f
C1039 VINN.n555 a_n3166_n47928 0.026615f
C1040 VINN.n556 a_n3166_n47928 0.026615f
C1041 VINN.n557 a_n3166_n47928 0.026615f
C1042 VINN.n558 a_n3166_n47928 0.026615f
C1043 VINN.n559 a_n3166_n47928 0.026615f
C1044 VINN.n560 a_n3166_n47928 0.026615f
C1045 VINN.n561 a_n3166_n47928 0.026615f
C1046 VINN.n562 a_n3166_n47928 0.026615f
C1047 VINN.n563 a_n3166_n47928 0.026615f
C1048 VINN.n564 a_n3166_n47928 0.026615f
C1049 VINN.n565 a_n3166_n47928 0.026615f
C1050 VINN.n566 a_n3166_n47928 0.026615f
C1051 VINN.n567 a_n3166_n47928 0.026615f
C1052 VINN.n568 a_n3166_n47928 0.026615f
C1053 VINN.n569 a_n3166_n47928 0.026615f
C1054 VINN.n570 a_n3166_n47928 0.026615f
C1055 VINN.n571 a_n3166_n47928 0.026615f
C1056 VINN.n572 a_n3166_n47928 0.026615f
C1057 VINN.n573 a_n3166_n47928 0.026615f
C1058 VINN.n574 a_n3166_n47928 0.015454f
C1059 VINN.n575 a_n3166_n47928 0.024469f
C1060 VINN.n576 a_n3166_n47928 0.026615f
C1061 VINN.n577 a_n3166_n47928 0.026615f
C1062 VINN.n578 a_n3166_n47928 0.026615f
C1063 VINN.n579 a_n3166_n47928 0.026615f
C1064 VINN.n580 a_n3166_n47928 0.026615f
C1065 VINN.n581 a_n3166_n47928 0.026615f
C1066 VINN.n582 a_n3166_n47928 0.026615f
C1067 VINN.n583 a_n3166_n47928 0.026615f
C1068 VINN.n584 a_n3166_n47928 0.026615f
C1069 VINN.n585 a_n3166_n47928 0.026615f
C1070 VINN.n586 a_n3166_n47928 0.026615f
C1071 VINN.n587 a_n3166_n47928 0.026615f
C1072 VINN.n588 a_n3166_n47928 0.026615f
C1073 VINN.n589 a_n3166_n47928 0.026615f
C1074 VINN.n590 a_n3166_n47928 0.026615f
C1075 VINN.n591 a_n3166_n47928 0.026615f
C1076 VINN.n592 a_n3166_n47928 0.026615f
C1077 VINN.n593 a_n3166_n47928 0.026615f
C1078 VINN.n594 a_n3166_n47928 0.026615f
C1079 VINN.n595 a_n3166_n47928 0.026615f
C1080 VINN.n596 a_n3166_n47928 0.026615f
C1081 VINN.n597 a_n3166_n47928 0.026615f
C1082 VINN.n598 a_n3166_n47928 0.026615f
C1083 VINN.n599 a_n3166_n47928 0.026615f
C1084 VINN.n600 a_n3166_n47928 0.026615f
C1085 VINN.n601 a_n3166_n47928 0.026615f
C1086 VINN.n602 a_n3166_n47928 0.026615f
C1087 VINN.n603 a_n3166_n47928 0.026615f
C1088 VINN.n604 a_n3166_n47928 0.026615f
C1089 VINN.n605 a_n3166_n47928 0.026615f
C1090 VINN.n606 a_n3166_n47928 0.026615f
C1091 VINN.n607 a_n3166_n47928 0.026615f
C1092 VINN.n608 a_n3166_n47928 0.026615f
C1093 VINN.n609 a_n3166_n47928 0.026615f
C1094 VINN.n610 a_n3166_n47928 0.026615f
C1095 VINN.n611 a_n3166_n47928 0.026615f
C1096 VINN.n612 a_n3166_n47928 0.026615f
C1097 VINN.n613 a_n3166_n47928 0.026615f
C1098 VINN.n614 a_n3166_n47928 0.026615f
C1099 VINN.n615 a_n3166_n47928 0.026615f
C1100 VINN.n616 a_n3166_n47928 0.026615f
C1101 VINN.n617 a_n3166_n47928 0.026615f
C1102 VINN.n618 a_n3166_n47928 0.026615f
C1103 VINN.n619 a_n3166_n47928 0.026615f
C1104 VINN.n620 a_n3166_n47928 0.026615f
C1105 VINN.n621 a_n3166_n47928 0.026615f
C1106 VINN.n622 a_n3166_n47928 0.026615f
C1107 VINN.n623 a_n3166_n47928 0.026615f
C1108 VINN.n624 a_n3166_n47928 0.026615f
C1109 VINN.n625 a_n3166_n47928 0.026615f
C1110 VINN.n626 a_n3166_n47928 0.026615f
C1111 VINN.n627 a_n3166_n47928 0.026615f
C1112 VINN.n628 a_n3166_n47928 0.026615f
C1113 VINN.n629 a_n3166_n47928 0.026615f
C1114 VINN.n630 a_n3166_n47928 0.026615f
C1115 VINN.n631 a_n3166_n47928 0.026615f
C1116 VINN.n632 a_n3166_n47928 0.026615f
C1117 VINN.n633 a_n3166_n47928 0.026615f
C1118 VINN.n634 a_n3166_n47928 0.026615f
C1119 VINN.n635 a_n3166_n47928 0.026615f
C1120 VINN.n636 a_n3166_n47928 0.026615f
C1121 VINN.n637 a_n3166_n47928 0.026615f
C1122 VINN.n638 a_n3166_n47928 0.026615f
C1123 VINN.n639 a_n3166_n47928 0.026615f
C1124 VINN.n640 a_n3166_n47928 0.026615f
C1125 VINN.n641 a_n3166_n47928 0.026615f
C1126 VINN.n642 a_n3166_n47928 0.026615f
C1127 VINN.n643 a_n3166_n47928 0.026615f
C1128 VINN.n644 a_n3166_n47928 0.026615f
C1129 VINN.n645 a_n3166_n47928 0.026615f
C1130 VINN.n646 a_n3166_n47928 0.026615f
C1131 VINN.n647 a_n3166_n47928 0.026615f
C1132 VINN.n648 a_n3166_n47928 0.026615f
C1133 VINN.n649 a_n3166_n47928 0.026615f
C1134 VINN.n650 a_n3166_n47928 0.026615f
C1135 VINN.n651 a_n3166_n47928 0.026615f
C1136 VINN.n652 a_n3166_n47928 0.026615f
C1137 VINN.n653 a_n3166_n47928 0.026615f
C1138 VINN.n654 a_n3166_n47928 0.026615f
C1139 VINN.n655 a_n3166_n47928 0.026615f
C1140 VINN.n656 a_n3166_n47928 0.026615f
C1141 VINN.n657 a_n3166_n47928 0.026615f
C1142 VINN.n658 a_n3166_n47928 0.053303f
C1143 w_1750_n43456.t12 a_n3166_n47928 0.022964f
C1144 w_1750_n43456.t32 a_n3166_n47928 0.022964f
C1145 w_1750_n43456.t22 a_n3166_n47928 0.022964f
C1146 w_1750_n43456.n0 a_n3166_n47928 0.10128f
C1147 w_1750_n43456.n1 a_n3166_n47928 0.242037f
C1148 w_1750_n43456.t2 a_n3166_n47928 0.184813f
C1149 w_1750_n43456.t0 a_n3166_n47928 0.022964f
C1150 w_1750_n43456.t1 a_n3166_n47928 0.022964f
C1151 w_1750_n43456.n2 a_n3166_n47928 0.114077f
C1152 w_1750_n43456.n3 a_n3166_n47928 0.32976f
C1153 w_1750_n43456.t43 a_n3166_n47928 0.181507f
C1154 w_1750_n43456.n4 a_n3166_n47928 0.689281f
C1155 w_1750_n43456.t79 a_n3166_n47928 0.022964f
C1156 w_1750_n43456.t55 a_n3166_n47928 0.022964f
C1157 w_1750_n43456.n5 a_n3166_n47928 0.10128f
C1158 w_1750_n43456.n6 a_n3166_n47928 0.247084f
C1159 w_1750_n43456.n7 a_n3166_n47928 0.310379f
C1160 w_1750_n43456.n8 a_n3166_n47928 0.341362f
C1161 w_1750_n43456.n9 a_n3166_n47928 0.341362f
C1162 w_1750_n43456.n10 a_n3166_n47928 0.341362f
C1163 w_1750_n43456.t59 a_n3166_n47928 0.022964f
C1164 w_1750_n43456.t71 a_n3166_n47928 0.022964f
C1165 w_1750_n43456.n11 a_n3166_n47928 0.10128f
C1166 w_1750_n43456.n12 a_n3166_n47928 0.242037f
C1167 w_1750_n43456.t81 a_n3166_n47928 0.022964f
C1168 w_1750_n43456.t63 a_n3166_n47928 0.022964f
C1169 w_1750_n43456.n13 a_n3166_n47928 0.10128f
C1170 w_1750_n43456.n14 a_n3166_n47928 0.242037f
C1171 w_1750_n43456.t73 a_n3166_n47928 0.022964f
C1172 w_1750_n43456.t47 a_n3166_n47928 0.022964f
C1173 w_1750_n43456.n15 a_n3166_n47928 0.10128f
C1174 w_1750_n43456.n16 a_n3166_n47928 0.242037f
C1175 w_1750_n43456.t57 a_n3166_n47928 0.022964f
C1176 w_1750_n43456.t65 a_n3166_n47928 0.022964f
C1177 w_1750_n43456.n17 a_n3166_n47928 0.10128f
C1178 w_1750_n43456.n18 a_n3166_n47928 0.242037f
C1179 w_1750_n43456.t49 a_n3166_n47928 0.022964f
C1180 w_1750_n43456.t45 a_n3166_n47928 0.022964f
C1181 w_1750_n43456.n19 a_n3166_n47928 0.10128f
C1182 w_1750_n43456.n20 a_n3166_n47928 0.242037f
C1183 w_1750_n43456.t67 a_n3166_n47928 0.022964f
C1184 w_1750_n43456.t83 a_n3166_n47928 0.022964f
C1185 w_1750_n43456.n21 a_n3166_n47928 0.10128f
C1186 w_1750_n43456.n22 a_n3166_n47928 0.242037f
C1187 w_1750_n43456.t51 a_n3166_n47928 0.022964f
C1188 w_1750_n43456.t75 a_n3166_n47928 0.022964f
C1189 w_1750_n43456.n23 a_n3166_n47928 0.10128f
C1190 w_1750_n43456.n24 a_n3166_n47928 0.242037f
C1191 w_1750_n43456.t69 a_n3166_n47928 0.022964f
C1192 w_1750_n43456.t53 a_n3166_n47928 0.022964f
C1193 w_1750_n43456.n25 a_n3166_n47928 0.10128f
C1194 w_1750_n43456.n26 a_n3166_n47928 0.242037f
C1195 w_1750_n43456.t61 a_n3166_n47928 0.022964f
C1196 w_1750_n43456.t77 a_n3166_n47928 0.022964f
C1197 w_1750_n43456.n27 a_n3166_n47928 0.10128f
C1198 w_1750_n43456.n28 a_n3166_n47928 0.400689f
C1199 w_1750_n43456.n29 a_n3166_n47928 0.188588f
C1200 w_1750_n43456.n30 a_n3166_n47928 0.189656f
C1201 w_1750_n43456.n31 a_n3166_n47928 1.01358f
C1202 w_1750_n43456.t76 a_n3166_n47928 0.565734f
C1203 w_1750_n43456.t60 a_n3166_n47928 0.434708f
C1204 w_1750_n43456.t52 a_n3166_n47928 0.434708f
C1205 w_1750_n43456.t68 a_n3166_n47928 0.434708f
C1206 w_1750_n43456.t74 a_n3166_n47928 0.434708f
C1207 w_1750_n43456.t50 a_n3166_n47928 0.434708f
C1208 w_1750_n43456.t82 a_n3166_n47928 0.434708f
C1209 w_1750_n43456.t66 a_n3166_n47928 0.434708f
C1210 w_1750_n43456.t44 a_n3166_n47928 0.434708f
C1211 w_1750_n43456.t48 a_n3166_n47928 0.326031f
C1212 w_1750_n43456.n32 a_n3166_n47928 0.217354f
C1213 w_1750_n43456.t64 a_n3166_n47928 0.326031f
C1214 w_1750_n43456.t56 a_n3166_n47928 0.434708f
C1215 w_1750_n43456.t46 a_n3166_n47928 0.434708f
C1216 w_1750_n43456.t72 a_n3166_n47928 0.434708f
C1217 w_1750_n43456.t62 a_n3166_n47928 0.434708f
C1218 w_1750_n43456.t80 a_n3166_n47928 0.434708f
C1219 w_1750_n43456.t70 a_n3166_n47928 0.434708f
C1220 w_1750_n43456.t58 a_n3166_n47928 0.434708f
C1221 w_1750_n43456.t54 a_n3166_n47928 0.434708f
C1222 w_1750_n43456.t78 a_n3166_n47928 0.565734f
C1223 w_1750_n43456.n33 a_n3166_n47928 1.01358f
C1224 w_1750_n43456.n34 a_n3166_n47928 0.189656f
C1225 w_1750_n43456.n35 a_n3166_n47928 0.18425f
C1226 w_1750_n43456.n36 a_n3166_n47928 0.324498f
C1227 w_1750_n43456.n37 a_n3166_n47928 0.868456f
C1228 w_1750_n43456.n38 a_n3166_n47928 0.18977f
C1229 w_1750_n43456.t30 a_n3166_n47928 0.022964f
C1230 w_1750_n43456.t4 a_n3166_n47928 0.022964f
C1231 w_1750_n43456.n39 a_n3166_n47928 0.10128f
C1232 w_1750_n43456.n40 a_n3166_n47928 0.400689f
C1233 w_1750_n43456.n41 a_n3166_n47928 0.188588f
C1234 w_1750_n43456.n42 a_n3166_n47928 1.01358f
C1235 w_1750_n43456.n43 a_n3166_n47928 1.01358f
C1236 w_1750_n43456.t29 a_n3166_n47928 0.565734f
C1237 w_1750_n43456.t3 a_n3166_n47928 0.434708f
C1238 w_1750_n43456.t31 a_n3166_n47928 0.434708f
C1239 w_1750_n43456.t21 a_n3166_n47928 0.434708f
C1240 w_1750_n43456.t11 a_n3166_n47928 0.434708f
C1241 w_1750_n43456.t41 a_n3166_n47928 0.434708f
C1242 w_1750_n43456.t17 a_n3166_n47928 0.434708f
C1243 w_1750_n43456.t5 a_n3166_n47928 0.434708f
C1244 w_1750_n43456.t37 a_n3166_n47928 0.434708f
C1245 w_1750_n43456.t27 a_n3166_n47928 0.326031f
C1246 w_1750_n43456.n44 a_n3166_n47928 0.189656f
C1247 w_1750_n43456.n45 a_n3166_n47928 0.341362f
C1248 w_1750_n43456.n46 a_n3166_n47928 0.341362f
C1249 w_1750_n43456.t13 a_n3166_n47928 0.565734f
C1250 w_1750_n43456.t23 a_n3166_n47928 0.434708f
C1251 w_1750_n43456.t7 a_n3166_n47928 0.434708f
C1252 w_1750_n43456.t39 a_n3166_n47928 0.434708f
C1253 w_1750_n43456.t25 a_n3166_n47928 0.434708f
C1254 w_1750_n43456.t35 a_n3166_n47928 0.434708f
C1255 w_1750_n43456.t9 a_n3166_n47928 0.434708f
C1256 w_1750_n43456.t19 a_n3166_n47928 0.434708f
C1257 w_1750_n43456.t33 a_n3166_n47928 0.434708f
C1258 w_1750_n43456.t15 a_n3166_n47928 0.326031f
C1259 w_1750_n43456.n47 a_n3166_n47928 0.217354f
C1260 w_1750_n43456.n48 a_n3166_n47928 0.341362f
C1261 w_1750_n43456.n49 a_n3166_n47928 0.310256f
C1262 w_1750_n43456.n50 a_n3166_n47928 0.184258f
C1263 w_1750_n43456.n51 a_n3166_n47928 0.309357f
C1264 w_1750_n43456.t24 a_n3166_n47928 0.022964f
C1265 w_1750_n43456.t14 a_n3166_n47928 0.022964f
C1266 w_1750_n43456.n52 a_n3166_n47928 0.10128f
C1267 w_1750_n43456.n53 a_n3166_n47928 0.247084f
C1268 w_1750_n43456.t40 a_n3166_n47928 0.022964f
C1269 w_1750_n43456.t8 a_n3166_n47928 0.022964f
C1270 w_1750_n43456.n54 a_n3166_n47928 0.10128f
C1271 w_1750_n43456.n55 a_n3166_n47928 0.242037f
C1272 w_1750_n43456.t36 a_n3166_n47928 0.022964f
C1273 w_1750_n43456.t26 a_n3166_n47928 0.022964f
C1274 w_1750_n43456.n56 a_n3166_n47928 0.10128f
C1275 w_1750_n43456.n57 a_n3166_n47928 0.242037f
C1276 w_1750_n43456.t20 a_n3166_n47928 0.022964f
C1277 w_1750_n43456.t10 a_n3166_n47928 0.022964f
C1278 w_1750_n43456.n58 a_n3166_n47928 0.10128f
C1279 w_1750_n43456.n59 a_n3166_n47928 0.242037f
C1280 w_1750_n43456.t16 a_n3166_n47928 0.022964f
C1281 w_1750_n43456.t34 a_n3166_n47928 0.022964f
C1282 w_1750_n43456.n60 a_n3166_n47928 0.10128f
C1283 w_1750_n43456.n61 a_n3166_n47928 0.242037f
C1284 w_1750_n43456.t38 a_n3166_n47928 0.022964f
C1285 w_1750_n43456.t28 a_n3166_n47928 0.022964f
C1286 w_1750_n43456.n62 a_n3166_n47928 0.10128f
C1287 w_1750_n43456.n63 a_n3166_n47928 0.242037f
C1288 w_1750_n43456.t18 a_n3166_n47928 0.022964f
C1289 w_1750_n43456.t6 a_n3166_n47928 0.022964f
C1290 w_1750_n43456.n64 a_n3166_n47928 0.10128f
C1291 w_1750_n43456.n65 a_n3166_n47928 0.242037f
C1292 w_1750_n43456.n66 a_n3166_n47928 0.242037f
C1293 w_1750_n43456.n67 a_n3166_n47928 0.10128f
C1294 w_1750_n43456.t42 a_n3166_n47928 0.022964f
C1295 VINP.n0 a_n3166_n47928 0.028463f
C1296 VINP.n1 a_n3166_n47928 0.027648f
C1297 VINP.n85 a_n3166_n47928 0.032056f
C1298 VINP.n86 a_n3166_n47928 0.059566f
C1299 VINP.n87 a_n3166_n47928 0.027648f
C1300 VINP.n88 a_n3166_n47928 0.027648f
C1301 VINP.n89 a_n3166_n47928 0.027648f
C1302 VINP.n90 a_n3166_n47928 0.027648f
C1303 VINP.n91 a_n3166_n47928 0.027648f
C1304 VINP.n92 a_n3166_n47928 0.027648f
C1305 VINP.n93 a_n3166_n47928 0.027648f
C1306 VINP.n94 a_n3166_n47928 0.027648f
C1307 VINP.n95 a_n3166_n47928 0.027648f
C1308 VINP.n96 a_n3166_n47928 0.027648f
C1309 VINP.n97 a_n3166_n47928 0.027648f
C1310 VINP.n98 a_n3166_n47928 0.027648f
C1311 VINP.n99 a_n3166_n47928 0.027648f
C1312 VINP.n100 a_n3166_n47928 0.027648f
C1313 VINP.n101 a_n3166_n47928 0.027648f
C1314 VINP.n102 a_n3166_n47928 0.027648f
C1315 VINP.n103 a_n3166_n47928 0.027648f
C1316 VINP.n104 a_n3166_n47928 0.027648f
C1317 VINP.n105 a_n3166_n47928 0.027648f
C1318 VINP.n106 a_n3166_n47928 0.027648f
C1319 VINP.n107 a_n3166_n47928 0.027648f
C1320 VINP.n108 a_n3166_n47928 0.027648f
C1321 VINP.n109 a_n3166_n47928 0.027648f
C1322 VINP.n110 a_n3166_n47928 0.027648f
C1323 VINP.n111 a_n3166_n47928 0.027648f
C1324 VINP.n112 a_n3166_n47928 0.027648f
C1325 VINP.n113 a_n3166_n47928 0.027648f
C1326 VINP.n114 a_n3166_n47928 0.027648f
C1327 VINP.n115 a_n3166_n47928 0.027648f
C1328 VINP.n116 a_n3166_n47928 0.027648f
C1329 VINP.n117 a_n3166_n47928 0.027648f
C1330 VINP.n118 a_n3166_n47928 0.027648f
C1331 VINP.n119 a_n3166_n47928 0.027648f
C1332 VINP.n120 a_n3166_n47928 0.027648f
C1333 VINP.n121 a_n3166_n47928 0.027648f
C1334 VINP.n122 a_n3166_n47928 0.027648f
C1335 VINP.n123 a_n3166_n47928 0.027648f
C1336 VINP.n124 a_n3166_n47928 0.027648f
C1337 VINP.n125 a_n3166_n47928 0.027648f
C1338 VINP.n126 a_n3166_n47928 0.027648f
C1339 VINP.n127 a_n3166_n47928 0.027648f
C1340 VINP.n128 a_n3166_n47928 0.027648f
C1341 VINP.n129 a_n3166_n47928 0.027648f
C1342 VINP.n130 a_n3166_n47928 0.027648f
C1343 VINP.n131 a_n3166_n47928 0.027648f
C1344 VINP.n132 a_n3166_n47928 0.027648f
C1345 VINP.n133 a_n3166_n47928 0.027648f
C1346 VINP.n134 a_n3166_n47928 0.027648f
C1347 VINP.n135 a_n3166_n47928 0.027648f
C1348 VINP.n136 a_n3166_n47928 0.027648f
C1349 VINP.n137 a_n3166_n47928 0.027648f
C1350 VINP.n138 a_n3166_n47928 0.027648f
C1351 VINP.n139 a_n3166_n47928 0.027648f
C1352 VINP.n140 a_n3166_n47928 0.027648f
C1353 VINP.n141 a_n3166_n47928 0.027648f
C1354 VINP.n142 a_n3166_n47928 0.027648f
C1355 VINP.n143 a_n3166_n47928 0.027648f
C1356 VINP.n144 a_n3166_n47928 0.027648f
C1357 VINP.n145 a_n3166_n47928 0.027648f
C1358 VINP.n146 a_n3166_n47928 0.027648f
C1359 VINP.n147 a_n3166_n47928 0.027648f
C1360 VINP.n148 a_n3166_n47928 0.027648f
C1361 VINP.n149 a_n3166_n47928 0.027648f
C1362 VINP.n151 a_n3166_n47928 0.027648f
C1363 VINP.n152 a_n3166_n47928 0.027648f
C1364 VINP.n153 a_n3166_n47928 0.027648f
C1365 VINP.n154 a_n3166_n47928 0.027648f
C1366 VINP.n155 a_n3166_n47928 0.027648f
C1367 VINP.n156 a_n3166_n47928 0.027648f
C1368 VINP.n157 a_n3166_n47928 0.027648f
C1369 VINP.n158 a_n3166_n47928 0.027648f
C1370 VINP.n159 a_n3166_n47928 0.027648f
C1371 VINP.n160 a_n3166_n47928 0.027648f
C1372 VINP.n161 a_n3166_n47928 0.027648f
C1373 VINP.n162 a_n3166_n47928 0.027648f
C1374 VINP.n163 a_n3166_n47928 0.027648f
C1375 VINP.n164 a_n3166_n47928 0.027648f
C1376 VINP.n165 a_n3166_n47928 0.027648f
C1377 VINP.n166 a_n3166_n47928 0.027648f
C1378 VINP.n167 a_n3166_n47928 0.027648f
C1379 VINP.n168 a_n3166_n47928 0.027648f
C1380 VINP.n169 a_n3166_n47928 0.027648f
C1381 VINP.n170 a_n3166_n47928 0.027648f
C1382 VINP.n171 a_n3166_n47928 0.027648f
C1383 VINP.n172 a_n3166_n47928 0.027648f
C1384 VINP.n173 a_n3166_n47928 0.027648f
C1385 VINP.n174 a_n3166_n47928 0.027648f
C1386 VINP.n175 a_n3166_n47928 0.027648f
C1387 VINP.n176 a_n3166_n47928 0.027648f
C1388 VINP.n177 a_n3166_n47928 0.027648f
C1389 VINP.n178 a_n3166_n47928 0.027648f
C1390 VINP.n179 a_n3166_n47928 0.027648f
C1391 VINP.n180 a_n3166_n47928 0.027648f
C1392 VINP.n181 a_n3166_n47928 0.027648f
C1393 VINP.n182 a_n3166_n47928 0.027648f
C1394 VINP.n183 a_n3166_n47928 0.027648f
C1395 VINP.n184 a_n3166_n47928 0.027648f
C1396 VINP.n185 a_n3166_n47928 0.027648f
C1397 VINP.n186 a_n3166_n47928 0.027648f
C1398 VINP.n187 a_n3166_n47928 0.027648f
C1399 VINP.n188 a_n3166_n47928 0.027648f
C1400 VINP.n189 a_n3166_n47928 0.027648f
C1401 VINP.n190 a_n3166_n47928 0.027648f
C1402 VINP.n191 a_n3166_n47928 0.027648f
C1403 VINP.n192 a_n3166_n47928 0.027648f
C1404 VINP.n193 a_n3166_n47928 0.027648f
C1405 VINP.n194 a_n3166_n47928 0.027648f
C1406 VINP.n195 a_n3166_n47928 0.027648f
C1407 VINP.n196 a_n3166_n47928 0.027648f
C1408 VINP.n197 a_n3166_n47928 0.027648f
C1409 VINP.n198 a_n3166_n47928 0.027648f
C1410 VINP.n199 a_n3166_n47928 0.027648f
C1411 VINP.n200 a_n3166_n47928 0.027648f
C1412 VINP.n201 a_n3166_n47928 0.027648f
C1413 VINP.n202 a_n3166_n47928 0.027648f
C1414 VINP.n203 a_n3166_n47928 0.027648f
C1415 VINP.n204 a_n3166_n47928 0.027648f
C1416 VINP.n205 a_n3166_n47928 0.027648f
C1417 VINP.n206 a_n3166_n47928 0.027648f
C1418 VINP.n207 a_n3166_n47928 0.027648f
C1419 VINP.n208 a_n3166_n47928 0.027648f
C1420 VINP.n209 a_n3166_n47928 0.027648f
C1421 VINP.n210 a_n3166_n47928 0.027648f
C1422 VINP.n211 a_n3166_n47928 0.027648f
C1423 VINP.n212 a_n3166_n47928 0.027648f
C1424 VINP.n213 a_n3166_n47928 0.027648f
C1425 VINP.n215 a_n3166_n47928 0.027648f
C1426 VINP.n216 a_n3166_n47928 0.027648f
C1427 VINP.n217 a_n3166_n47928 0.027648f
C1428 VINP.n218 a_n3166_n47928 0.027648f
C1429 VINP.n219 a_n3166_n47928 0.027648f
C1430 VINP.n220 a_n3166_n47928 0.027648f
C1431 VINP.n221 a_n3166_n47928 0.027648f
C1432 VINP.n222 a_n3166_n47928 0.027648f
C1433 VINP.n223 a_n3166_n47928 0.027648f
C1434 VINP.n224 a_n3166_n47928 0.027648f
C1435 VINP.n225 a_n3166_n47928 0.027648f
C1436 VINP.n226 a_n3166_n47928 0.027648f
C1437 VINP.n227 a_n3166_n47928 0.027648f
C1438 VINP.n228 a_n3166_n47928 0.027648f
C1439 VINP.n229 a_n3166_n47928 0.027648f
C1440 VINP.n230 a_n3166_n47928 0.027648f
C1441 VINP.n231 a_n3166_n47928 0.027648f
C1442 VINP.n232 a_n3166_n47928 0.027648f
C1443 VINP.n233 a_n3166_n47928 0.027648f
C1444 VINP.n234 a_n3166_n47928 0.027648f
C1445 VINP.n235 a_n3166_n47928 0.027648f
C1446 VINP.n236 a_n3166_n47928 0.027648f
C1447 VINP.n237 a_n3166_n47928 0.027648f
C1448 VINP.n238 a_n3166_n47928 0.027648f
C1449 VINP.n239 a_n3166_n47928 0.027648f
C1450 VINP.n240 a_n3166_n47928 0.027648f
C1451 VINP.n241 a_n3166_n47928 0.027648f
C1452 VINP.n242 a_n3166_n47928 0.027648f
C1453 VINP.n243 a_n3166_n47928 0.027648f
C1454 VINP.n244 a_n3166_n47928 0.027648f
C1455 VINP.n245 a_n3166_n47928 0.027648f
C1456 VINP.n246 a_n3166_n47928 0.027648f
C1457 VINP.n247 a_n3166_n47928 0.027648f
C1458 VINP.n248 a_n3166_n47928 0.027648f
C1459 VINP.n249 a_n3166_n47928 0.027648f
C1460 VINP.n250 a_n3166_n47928 0.027648f
C1461 VINP.n251 a_n3166_n47928 0.027648f
C1462 VINP.n252 a_n3166_n47928 0.027648f
C1463 VINP.n253 a_n3166_n47928 0.027648f
C1464 VINP.n254 a_n3166_n47928 0.027648f
C1465 VINP.n255 a_n3166_n47928 0.027648f
C1466 VINP.n256 a_n3166_n47928 0.027648f
C1467 VINP.n257 a_n3166_n47928 0.027648f
C1468 VINP.n258 a_n3166_n47928 0.027648f
C1469 VINP.n259 a_n3166_n47928 0.027648f
C1470 VINP.n260 a_n3166_n47928 0.027648f
C1471 VINP.n261 a_n3166_n47928 0.027648f
C1472 VINP.n262 a_n3166_n47928 0.027648f
C1473 VINP.n263 a_n3166_n47928 0.027648f
C1474 VINP.n264 a_n3166_n47928 0.027648f
C1475 VINP.n265 a_n3166_n47928 0.027648f
C1476 VINP.n266 a_n3166_n47928 0.027648f
C1477 VINP.n267 a_n3166_n47928 0.027648f
C1478 VINP.n268 a_n3166_n47928 0.027648f
C1479 VINP.n269 a_n3166_n47928 0.027648f
C1480 VINP.n270 a_n3166_n47928 0.027648f
C1481 VINP.n271 a_n3166_n47928 0.027648f
C1482 VINP.n272 a_n3166_n47928 0.027648f
C1483 VINP.n273 a_n3166_n47928 0.027648f
C1484 VINP.n274 a_n3166_n47928 0.027648f
C1485 VINP.n275 a_n3166_n47928 0.027648f
C1486 VINP.n276 a_n3166_n47928 0.027648f
C1487 VINP.n278 a_n3166_n47928 0.028463f
C1488 VINP.n280 a_n3166_n47928 0.027648f
C1489 VINP.n282 a_n3166_n47928 0.027648f
C1490 VINP.n284 a_n3166_n47928 0.027648f
C1491 VINP.n286 a_n3166_n47928 0.027648f
C1492 VINP.n288 a_n3166_n47928 0.027648f
C1493 VINP.n290 a_n3166_n47928 0.027648f
C1494 VINP.n292 a_n3166_n47928 0.027648f
C1495 VINP.n294 a_n3166_n47928 0.027648f
C1496 VINP.n296 a_n3166_n47928 0.027648f
C1497 VINP.n298 a_n3166_n47928 0.027648f
C1498 VINP.n300 a_n3166_n47928 0.027648f
C1499 VINP.n302 a_n3166_n47928 0.027648f
C1500 VINP.n304 a_n3166_n47928 0.027648f
C1501 VINP.n306 a_n3166_n47928 0.027648f
C1502 VINP.n308 a_n3166_n47928 0.027648f
C1503 VINP.n310 a_n3166_n47928 0.027648f
C1504 VINP.n312 a_n3166_n47928 0.027648f
C1505 VINP.n314 a_n3166_n47928 0.027648f
C1506 VINP.n316 a_n3166_n47928 0.027648f
C1507 VINP.n318 a_n3166_n47928 0.027648f
C1508 VINP.n320 a_n3166_n47928 0.027648f
C1509 VINP.n322 a_n3166_n47928 0.027648f
C1510 VINP.n324 a_n3166_n47928 0.027648f
C1511 VINP.n326 a_n3166_n47928 0.027648f
C1512 VINP.n328 a_n3166_n47928 0.027648f
C1513 VINP.n330 a_n3166_n47928 0.027648f
C1514 VINP.n332 a_n3166_n47928 0.027648f
C1515 VINP.n334 a_n3166_n47928 0.027648f
C1516 VINP.n336 a_n3166_n47928 0.027648f
C1517 VINP.n338 a_n3166_n47928 0.027648f
C1518 VINP.n340 a_n3166_n47928 0.027648f
C1519 VINP.n342 a_n3166_n47928 0.027648f
C1520 VINP.n344 a_n3166_n47928 0.027648f
C1521 VINP.n346 a_n3166_n47928 0.027648f
C1522 VINP.n348 a_n3166_n47928 0.027648f
C1523 VINP.n350 a_n3166_n47928 0.027648f
C1524 VINP.n352 a_n3166_n47928 0.027648f
C1525 VINP.n354 a_n3166_n47928 0.027648f
C1526 VINP.n356 a_n3166_n47928 0.027648f
C1527 VINP.n358 a_n3166_n47928 0.027648f
C1528 VINP.n360 a_n3166_n47928 0.027648f
C1529 VINP.n362 a_n3166_n47928 0.027648f
C1530 VINP.n364 a_n3166_n47928 0.027648f
C1531 VINP.n366 a_n3166_n47928 0.027648f
C1532 VINP.n368 a_n3166_n47928 0.027648f
C1533 VINP.n370 a_n3166_n47928 0.027648f
C1534 VINP.n372 a_n3166_n47928 0.027648f
C1535 VINP.n374 a_n3166_n47928 0.027648f
C1536 VINP.n376 a_n3166_n47928 0.027648f
C1537 VINP.n378 a_n3166_n47928 0.027648f
C1538 VINP.n380 a_n3166_n47928 0.027648f
C1539 VINP.n382 a_n3166_n47928 0.027648f
C1540 VINP.n384 a_n3166_n47928 0.027648f
C1541 VINP.n386 a_n3166_n47928 0.027648f
C1542 VINP.n388 a_n3166_n47928 0.027648f
C1543 VINP.n390 a_n3166_n47928 0.027648f
C1544 VINP.n392 a_n3166_n47928 0.027648f
C1545 VINP.n394 a_n3166_n47928 0.027648f
C1546 VINP.n396 a_n3166_n47928 0.027648f
C1547 VINP.n398 a_n3166_n47928 0.027648f
C1548 VINP.n400 a_n3166_n47928 0.027648f
C1549 VINP.n463 a_n3166_n47928 0.028094f
C1550 VINP.n528 a_n3166_n47928 0.027648f
C1551 VINP.n529 a_n3166_n47928 0.027648f
C1552 VINP.n530 a_n3166_n47928 0.055372f
C1553 VINP.n531 a_n3166_n47928 0.027648f
C1554 VINP.n532 a_n3166_n47928 0.027648f
C1555 VINP.n533 a_n3166_n47928 0.027648f
C1556 VINP.n534 a_n3166_n47928 0.027648f
C1557 VINP.n535 a_n3166_n47928 0.027648f
C1558 VINP.n536 a_n3166_n47928 0.027648f
C1559 VINP.n537 a_n3166_n47928 0.027648f
C1560 VINP.n538 a_n3166_n47928 0.027648f
C1561 VINP.n539 a_n3166_n47928 0.027648f
C1562 VINP.n540 a_n3166_n47928 0.027648f
C1563 VINP.n541 a_n3166_n47928 0.027648f
C1564 VINP.n542 a_n3166_n47928 0.027648f
C1565 VINP.n543 a_n3166_n47928 0.027648f
C1566 VINP.n544 a_n3166_n47928 0.027648f
C1567 VINP.n545 a_n3166_n47928 0.027648f
C1568 VINP.n546 a_n3166_n47928 0.027648f
C1569 VINP.n547 a_n3166_n47928 0.027648f
C1570 VINP.n548 a_n3166_n47928 0.027648f
C1571 VINP.n549 a_n3166_n47928 0.027648f
C1572 VINP.n550 a_n3166_n47928 0.027648f
C1573 VINP.n551 a_n3166_n47928 0.027648f
C1574 VINP.n552 a_n3166_n47928 0.027648f
C1575 VINP.n553 a_n3166_n47928 0.027648f
C1576 VINP.n554 a_n3166_n47928 0.027648f
C1577 VINP.n555 a_n3166_n47928 0.027648f
C1578 VINP.n556 a_n3166_n47928 0.027648f
C1579 VINP.n557 a_n3166_n47928 0.027648f
C1580 VINP.n558 a_n3166_n47928 0.027648f
C1581 VINP.n559 a_n3166_n47928 0.027648f
C1582 VINP.n560 a_n3166_n47928 0.027648f
C1583 VINP.n561 a_n3166_n47928 0.027648f
C1584 VINP.n562 a_n3166_n47928 0.027648f
C1585 VINP.n563 a_n3166_n47928 0.027648f
C1586 VINP.n564 a_n3166_n47928 0.027648f
C1587 VINP.n565 a_n3166_n47928 0.027648f
C1588 VINP.n566 a_n3166_n47928 0.027648f
C1589 VINP.n567 a_n3166_n47928 0.027648f
C1590 VINP.n568 a_n3166_n47928 0.027648f
C1591 VINP.n569 a_n3166_n47928 0.027648f
C1592 VINP.n570 a_n3166_n47928 0.027648f
C1593 VINP.n571 a_n3166_n47928 0.027648f
C1594 VINP.n572 a_n3166_n47928 0.027648f
C1595 VINP.n573 a_n3166_n47928 0.027648f
C1596 VINP.n574 a_n3166_n47928 0.016054f
C1597 VINP.n575 a_n3166_n47928 0.025418f
C1598 VINP.n576 a_n3166_n47928 0.027648f
C1599 VINP.n577 a_n3166_n47928 0.027648f
C1600 VINP.n578 a_n3166_n47928 0.027648f
C1601 VINP.n579 a_n3166_n47928 0.027648f
C1602 VINP.n580 a_n3166_n47928 0.027648f
C1603 VINP.n581 a_n3166_n47928 0.027648f
C1604 VINP.n582 a_n3166_n47928 0.027648f
C1605 VINP.n583 a_n3166_n47928 0.027648f
C1606 VINP.n584 a_n3166_n47928 0.027648f
C1607 VINP.n585 a_n3166_n47928 0.027648f
C1608 VINP.n586 a_n3166_n47928 0.027648f
C1609 VINP.n587 a_n3166_n47928 0.027648f
C1610 VINP.n588 a_n3166_n47928 0.027648f
C1611 VINP.n589 a_n3166_n47928 0.027648f
C1612 VINP.n590 a_n3166_n47928 0.027648f
C1613 VINP.n591 a_n3166_n47928 0.027648f
C1614 VINP.n592 a_n3166_n47928 0.027648f
C1615 VINP.n593 a_n3166_n47928 0.027648f
C1616 VINP.n594 a_n3166_n47928 0.027648f
C1617 VINP.n595 a_n3166_n47928 0.027648f
C1618 VINP.n596 a_n3166_n47928 0.027648f
C1619 VINP.n597 a_n3166_n47928 0.027648f
C1620 VINP.n598 a_n3166_n47928 0.027648f
C1621 VINP.n599 a_n3166_n47928 0.027648f
C1622 VINP.n600 a_n3166_n47928 0.027648f
C1623 VINP.n601 a_n3166_n47928 0.027648f
C1624 VINP.n602 a_n3166_n47928 0.027648f
C1625 VINP.n603 a_n3166_n47928 0.027648f
C1626 VINP.n604 a_n3166_n47928 0.027648f
C1627 VINP.n605 a_n3166_n47928 0.027648f
C1628 VINP.n606 a_n3166_n47928 0.027648f
C1629 VINP.n607 a_n3166_n47928 0.027648f
C1630 VINP.n608 a_n3166_n47928 0.027648f
C1631 VINP.n609 a_n3166_n47928 0.027648f
C1632 VINP.n610 a_n3166_n47928 0.027648f
C1633 VINP.n611 a_n3166_n47928 0.027648f
C1634 VINP.n612 a_n3166_n47928 0.027648f
C1635 VINP.n613 a_n3166_n47928 0.027648f
C1636 VINP.n614 a_n3166_n47928 0.027648f
C1637 VINP.n615 a_n3166_n47928 0.027648f
C1638 VINP.n616 a_n3166_n47928 0.027648f
C1639 VINP.n617 a_n3166_n47928 0.027648f
C1640 VINP.n618 a_n3166_n47928 0.027648f
C1641 VINP.n619 a_n3166_n47928 0.027648f
C1642 VINP.n620 a_n3166_n47928 0.027648f
C1643 VINP.n621 a_n3166_n47928 0.027648f
C1644 VINP.n622 a_n3166_n47928 0.027648f
C1645 VINP.n623 a_n3166_n47928 0.027648f
C1646 VINP.n624 a_n3166_n47928 0.027648f
C1647 VINP.n625 a_n3166_n47928 0.027648f
C1648 VINP.n626 a_n3166_n47928 0.027648f
C1649 VINP.n627 a_n3166_n47928 0.027648f
C1650 VINP.n628 a_n3166_n47928 0.027648f
C1651 VINP.n629 a_n3166_n47928 0.027648f
C1652 VINP.n630 a_n3166_n47928 0.027648f
C1653 VINP.n631 a_n3166_n47928 0.027648f
C1654 VINP.n632 a_n3166_n47928 0.027648f
C1655 VINP.n633 a_n3166_n47928 0.027648f
C1656 VINP.n634 a_n3166_n47928 0.027648f
C1657 VINP.n635 a_n3166_n47928 0.027648f
C1658 VINP.n636 a_n3166_n47928 0.027648f
C1659 VINP.n637 a_n3166_n47928 0.027648f
C1660 VINP.n638 a_n3166_n47928 0.027648f
C1661 VINP.n639 a_n3166_n47928 0.027648f
C1662 VINP.n640 a_n3166_n47928 0.027648f
C1663 VINP.n641 a_n3166_n47928 0.027648f
C1664 VINP.n642 a_n3166_n47928 0.027648f
C1665 VINP.n643 a_n3166_n47928 0.027648f
C1666 VINP.n644 a_n3166_n47928 0.027648f
C1667 VINP.n645 a_n3166_n47928 0.027648f
C1668 VINP.n646 a_n3166_n47928 0.027648f
C1669 VINP.n647 a_n3166_n47928 0.027648f
C1670 VINP.n648 a_n3166_n47928 0.027648f
C1671 VINP.n649 a_n3166_n47928 0.027648f
C1672 VINP.n650 a_n3166_n47928 0.027648f
C1673 VINP.n651 a_n3166_n47928 0.027648f
C1674 VINP.n652 a_n3166_n47928 0.027648f
C1675 VINP.n653 a_n3166_n47928 0.027648f
C1676 VINP.n654 a_n3166_n47928 0.027648f
C1677 VINP.n655 a_n3166_n47928 0.027648f
C1678 VINP.n656 a_n3166_n47928 0.027648f
C1679 VINP.n657 a_n3166_n47928 0.027648f
C1680 VINP.n658 a_n3166_n47928 0.055372f
C1681 a_16582_n43566.t0 a_n3166_n47928 0.045638f
C1682 a_16582_n43566.t1 a_n3166_n47928 0.046971f
C1683 a_16582_n43566.t2 a_n3166_n47928 1.2811f
C1684 a_16582_n43566.n0 a_n3166_n47928 0.626294f
C1685 a_n1924_n43526.n0 a_n3166_n47928 1.80049f
C1686 a_n1924_n43526.n1 a_n3166_n47928 1.14253f
C1687 a_n1924_n43526.t1 a_n3166_n47928 0.089578f
C1688 a_n1924_n43526.t3 a_n3166_n47928 0.090667f
C1689 a_n1924_n43526.t2 a_n3166_n47928 0.052808f
C1690 a_n1924_n43526.n2 a_n3166_n47928 0.524507f
C1691 a_n1924_n43526.t5 a_n3166_n47928 0.052995f
C1692 a_n1924_n43526.t7 a_n3166_n47928 0.052843f
C1693 a_n1924_n43526.t4 a_n3166_n47928 0.052985f
C1694 a_n1924_n43526.t6 a_n3166_n47928 0.052808f
C1695 a_n1924_n43526.t0 a_n3166_n47928 0.087791f
C1696 VSS.n457 a_n3166_n47928 3.80306f
C1697 VSS.t22 a_n3166_n47928 0.015535f
C1698 VSS.t34 a_n3166_n47928 0.01589f
C1699 VSS.t46 a_n3166_n47928 0.01589f
C1700 VSS.t24 a_n3166_n47928 0.01589f
C1701 VSS.t32 a_n3166_n47928 0.011492f
C1702 VSS.t38 a_n3166_n47928 0.01589f
C1703 VSS.t18 a_n3166_n47928 0.012343f
C1704 VSS.n707 a_n3166_n47928 0.025148f
C1705 VSS.n708 a_n3166_n47928 0.068597f
C1706 VSS.n774 a_n3166_n47928 0.019635f
C1707 VSS.n895 a_n3166_n47928 0.087068f
C1708 VSS.n1618 a_n3166_n47928 0.044194f
C1709 VSS.n1620 a_n3166_n47928 4.10856f
C1710 VSS.n1653 a_n3166_n47928 0.375855f
C1711 VSS.n1654 a_n3166_n47928 0.342108f
C1712 VSS.n1755 a_n3166_n47928 0.03732f
C1713 VSS.n2185 a_n3166_n47928 0.060581f
C1714 VSS.n2239 a_n3166_n47928 0.050011f
C1715 VSS.t4 a_n3166_n47928 0.035505f
C1716 VSS.n2242 a_n3166_n47928 0.024099f
C1717 VSS.n2727 a_n3166_n47928 0.011966f
C1718 VSS.n3049 a_n3166_n47928 0.011966f
C1719 VSS.n3053 a_n3166_n47928 0.132925f
C1720 VSS.n3054 a_n3166_n47928 0.127143f
C1721 VSS.n3422 a_n3166_n47928 0.020381f
C1722 VSS.t40 a_n3166_n47928 0.012698f
C1723 VSS.t20 a_n3166_n47928 0.010854f
C1724 VSS.t36 a_n3166_n47928 0.01589f
C1725 VSS.t16 a_n3166_n47928 0.014046f
C1726 VSS.n4027 a_n3166_n47928 0.024864f
C1727 VSS.n4028 a_n3166_n47928 0.037313f
C1728 VSS.t14 a_n3166_n47928 0.015039f
C1729 VSS.t12 a_n3166_n47928 0.018799f
C1730 VSS.n4160 a_n3166_n47928 0.054955f
C1731 VSS.n4188 a_n3166_n47928 0.119298f
C1732 VSS.n4412 a_n3166_n47928 0.011966f
C1733 VSS.n4499 a_n3166_n47928 0.011966f
C1734 VSS.n4503 a_n3166_n47928 0.124932f
C1735 OUT.n1 a_n3166_n47928 0.014657f
C1736 OUT.n18 a_n3166_n47928 0.044036f
C1737 OUT.t40 a_n3166_n47928 1.25476f
C1738 OUT.n19 a_n3166_n47928 1.52975f
C1739 OUT.n22 a_n3166_n47928 0.017449f
C1740 OUT.n38 a_n3166_n47928 0.193385f
C1741 OUT.n39 a_n3166_n47928 6.35792f
C1742 a_8360_n43060.n0 a_n3166_n47928 5.74752f
C1743 a_8360_n43060.n1 a_n3166_n47928 1.24635f
C1744 a_8360_n43060.n2 a_n3166_n47928 2.66138f
C1745 a_8360_n43060.t12 a_n3166_n47928 0.24864f
C1746 a_8360_n43060.t5 a_n3166_n47928 0.24864f
C1747 a_8360_n43060.t7 a_n3166_n47928 0.24864f
C1748 a_8360_n43060.t8 a_n3166_n47928 0.24864f
C1749 a_8360_n43060.t11 a_n3166_n47928 0.24864f
C1750 a_8360_n43060.t6 a_n3166_n47928 0.24864f
C1751 a_8360_n43060.t13 a_n3166_n47928 0.24864f
C1752 a_8360_n43060.t9 a_n3166_n47928 0.24864f
C1753 a_8360_n43060.t4 a_n3166_n47928 0.24864f
C1754 a_8360_n43060.t0 a_n3166_n47928 0.235766f
C1755 a_8360_n43060.n3 a_n3166_n47928 1.4279f
C1756 a_8360_n43060.t10 a_n3166_n47928 0.286989f
C1757 a_8360_n43060.t1 a_n3166_n47928 0.337431f
C1758 a_8360_n43060.t3 a_n3166_n47928 0.26955f
C1759 a_8360_n43060.t2 a_n3166_n47928 0.26321f
C1760 a_8360_n43060.t33 a_n3166_n47928 0.170043f
C1761 a_8360_n43060.t32 a_n3166_n47928 0.169661f
C1762 a_8360_n43060.t15 a_n3166_n47928 0.169661f
C1763 a_8360_n43060.t22 a_n3166_n47928 0.169661f
C1764 a_8360_n43060.t16 a_n3166_n47928 0.169661f
C1765 a_8360_n43060.t27 a_n3166_n47928 0.169661f
C1766 a_8360_n43060.t23 a_n3166_n47928 0.169661f
C1767 a_8360_n43060.t30 a_n3166_n47928 0.169661f
C1768 a_8360_n43060.t20 a_n3166_n47928 0.169661f
C1769 a_8360_n43060.t17 a_n3166_n47928 0.169661f
C1770 a_8360_n43060.t28 a_n3166_n47928 0.169661f
C1771 a_8360_n43060.t24 a_n3166_n47928 0.169661f
C1772 a_8360_n43060.t31 a_n3166_n47928 0.169661f
C1773 a_8360_n43060.t21 a_n3166_n47928 0.169661f
C1774 a_8360_n43060.t18 a_n3166_n47928 0.169661f
C1775 a_8360_n43060.t29 a_n3166_n47928 0.169661f
C1776 a_8360_n43060.t25 a_n3166_n47928 0.169661f
C1777 a_8360_n43060.t34 a_n3166_n47928 0.169661f
C1778 a_8360_n43060.t26 a_n3166_n47928 0.169661f
C1779 a_8360_n43060.t19 a_n3166_n47928 0.169661f
C1780 a_8360_n43060.n4 a_n3166_n47928 2.11049f
C1781 a_8360_n43060.t14 a_n3166_n47928 0.282053f
.ends

