magic
tech gf180mcuD
magscale 1 10
timestamp 1699608907
<< nwell >>
rect 1258 36416 78710 36934
rect 1258 34848 78710 35712
rect 1258 33280 78710 34144
rect 1258 31712 78710 32576
rect 1258 30144 78710 31008
rect 1258 28576 78710 29440
rect 1258 27008 78710 27872
rect 1258 25440 78710 26304
rect 1258 23872 78710 24736
rect 1258 22304 78710 23168
rect 1258 20736 78710 21600
rect 1258 19168 78710 20032
rect 1258 17600 78710 18464
rect 1258 16032 78710 16896
rect 1258 14464 78710 15328
rect 1258 12921 78710 13760
rect 1258 12896 10829 12921
rect 1258 12167 14413 12192
rect 1258 11353 78710 12167
rect 1258 11328 25320 11353
rect 1258 10599 10381 10624
rect 1258 9785 78710 10599
rect 1258 9760 16205 9785
rect 1258 9031 15800 9056
rect 1258 8217 78710 9031
rect 1258 8192 9933 8217
rect 1258 7463 36766 7488
rect 1258 6649 78710 7463
rect 1258 6624 7805 6649
rect 1258 5895 21736 5920
rect 1258 5081 78710 5895
rect 1258 5056 8968 5081
rect 1258 4327 12776 4352
rect 1258 3488 78710 4327
<< pwell >>
rect 1258 35712 78710 36416
rect 1258 34144 78710 34848
rect 1258 32576 78710 33280
rect 1258 31008 78710 31712
rect 1258 29440 78710 30144
rect 1258 27872 78710 28576
rect 1258 26304 78710 27008
rect 1258 24736 78710 25440
rect 1258 23168 78710 23872
rect 1258 21600 78710 22304
rect 1258 20032 78710 20736
rect 1258 18464 78710 19168
rect 1258 16896 78710 17600
rect 1258 15328 78710 16032
rect 1258 13760 78710 14464
rect 1258 12192 78710 12896
rect 1258 10624 78710 11328
rect 1258 9056 78710 9760
rect 1258 7488 78710 8192
rect 1258 5920 78710 6624
rect 1258 4352 78710 5056
rect 1258 3050 78710 3488
<< obsm1 >>
rect 1344 926 78784 36908
<< metal2 >>
rect 6272 0 6384 800
rect 6496 0 6608 800
rect 6720 0 6832 800
rect 6944 0 7056 800
rect 7168 0 7280 800
rect 7392 0 7504 800
rect 7616 0 7728 800
rect 7840 0 7952 800
rect 8064 0 8176 800
rect 8288 0 8400 800
rect 8512 0 8624 800
rect 8736 0 8848 800
rect 8960 0 9072 800
rect 9184 0 9296 800
rect 9408 0 9520 800
rect 9632 0 9744 800
rect 9856 0 9968 800
rect 10080 0 10192 800
rect 10304 0 10416 800
rect 10528 0 10640 800
rect 10752 0 10864 800
rect 10976 0 11088 800
rect 11200 0 11312 800
rect 11424 0 11536 800
rect 11648 0 11760 800
rect 11872 0 11984 800
rect 12096 0 12208 800
rect 12320 0 12432 800
rect 12544 0 12656 800
rect 12768 0 12880 800
rect 12992 0 13104 800
rect 13216 0 13328 800
rect 13440 0 13552 800
rect 13664 0 13776 800
rect 13888 0 14000 800
rect 14112 0 14224 800
rect 14336 0 14448 800
rect 14560 0 14672 800
rect 14784 0 14896 800
rect 15008 0 15120 800
rect 15232 0 15344 800
rect 15456 0 15568 800
rect 15680 0 15792 800
rect 15904 0 16016 800
rect 16128 0 16240 800
rect 16352 0 16464 800
rect 16576 0 16688 800
rect 16800 0 16912 800
rect 17024 0 17136 800
rect 17248 0 17360 800
rect 17472 0 17584 800
rect 17696 0 17808 800
rect 17920 0 18032 800
rect 18144 0 18256 800
rect 18368 0 18480 800
rect 18592 0 18704 800
rect 18816 0 18928 800
rect 19040 0 19152 800
rect 19264 0 19376 800
rect 19488 0 19600 800
rect 19712 0 19824 800
rect 19936 0 20048 800
rect 20160 0 20272 800
rect 20384 0 20496 800
rect 20608 0 20720 800
rect 20832 0 20944 800
rect 21056 0 21168 800
rect 21280 0 21392 800
rect 21504 0 21616 800
rect 21728 0 21840 800
rect 21952 0 22064 800
rect 22176 0 22288 800
rect 22400 0 22512 800
rect 22624 0 22736 800
rect 22848 0 22960 800
rect 23072 0 23184 800
rect 23296 0 23408 800
rect 23520 0 23632 800
rect 23744 0 23856 800
rect 23968 0 24080 800
rect 24192 0 24304 800
rect 24416 0 24528 800
rect 24640 0 24752 800
rect 24864 0 24976 800
rect 25088 0 25200 800
rect 25312 0 25424 800
rect 25536 0 25648 800
rect 25760 0 25872 800
rect 25984 0 26096 800
rect 26208 0 26320 800
rect 26432 0 26544 800
rect 26656 0 26768 800
rect 26880 0 26992 800
rect 27104 0 27216 800
rect 27328 0 27440 800
rect 27552 0 27664 800
rect 27776 0 27888 800
rect 28000 0 28112 800
rect 28224 0 28336 800
rect 28448 0 28560 800
rect 28672 0 28784 800
rect 28896 0 29008 800
rect 29120 0 29232 800
rect 29344 0 29456 800
rect 29568 0 29680 800
rect 29792 0 29904 800
rect 30016 0 30128 800
rect 30240 0 30352 800
rect 30464 0 30576 800
rect 30688 0 30800 800
rect 30912 0 31024 800
rect 31136 0 31248 800
rect 31360 0 31472 800
rect 31584 0 31696 800
rect 31808 0 31920 800
rect 32032 0 32144 800
rect 32256 0 32368 800
rect 32480 0 32592 800
rect 32704 0 32816 800
rect 32928 0 33040 800
rect 33152 0 33264 800
rect 33376 0 33488 800
rect 33600 0 33712 800
rect 33824 0 33936 800
rect 34048 0 34160 800
rect 34272 0 34384 800
rect 34496 0 34608 800
rect 34720 0 34832 800
rect 34944 0 35056 800
rect 35168 0 35280 800
rect 35392 0 35504 800
rect 35616 0 35728 800
rect 35840 0 35952 800
rect 36064 0 36176 800
rect 36288 0 36400 800
rect 36512 0 36624 800
rect 36736 0 36848 800
rect 36960 0 37072 800
rect 37184 0 37296 800
rect 37408 0 37520 800
rect 37632 0 37744 800
rect 37856 0 37968 800
rect 38080 0 38192 800
rect 38304 0 38416 800
rect 38528 0 38640 800
rect 38752 0 38864 800
rect 38976 0 39088 800
rect 39200 0 39312 800
rect 39424 0 39536 800
rect 39648 0 39760 800
rect 39872 0 39984 800
rect 40096 0 40208 800
rect 40320 0 40432 800
rect 40544 0 40656 800
rect 40768 0 40880 800
rect 40992 0 41104 800
rect 41216 0 41328 800
rect 41440 0 41552 800
rect 41664 0 41776 800
rect 41888 0 42000 800
rect 42112 0 42224 800
rect 42336 0 42448 800
rect 42560 0 42672 800
rect 42784 0 42896 800
rect 43008 0 43120 800
rect 43232 0 43344 800
rect 43456 0 43568 800
rect 43680 0 43792 800
rect 43904 0 44016 800
rect 44128 0 44240 800
rect 44352 0 44464 800
rect 44576 0 44688 800
rect 44800 0 44912 800
rect 45024 0 45136 800
rect 45248 0 45360 800
rect 45472 0 45584 800
rect 45696 0 45808 800
rect 45920 0 46032 800
rect 46144 0 46256 800
rect 46368 0 46480 800
rect 46592 0 46704 800
rect 46816 0 46928 800
rect 47040 0 47152 800
rect 47264 0 47376 800
rect 47488 0 47600 800
rect 47712 0 47824 800
rect 47936 0 48048 800
rect 48160 0 48272 800
rect 48384 0 48496 800
rect 48608 0 48720 800
rect 48832 0 48944 800
rect 49056 0 49168 800
rect 49280 0 49392 800
rect 49504 0 49616 800
rect 49728 0 49840 800
rect 49952 0 50064 800
rect 50176 0 50288 800
rect 50400 0 50512 800
rect 50624 0 50736 800
rect 50848 0 50960 800
rect 51072 0 51184 800
rect 51296 0 51408 800
rect 51520 0 51632 800
rect 51744 0 51856 800
rect 51968 0 52080 800
rect 52192 0 52304 800
rect 52416 0 52528 800
rect 52640 0 52752 800
rect 52864 0 52976 800
rect 53088 0 53200 800
rect 53312 0 53424 800
rect 53536 0 53648 800
rect 53760 0 53872 800
rect 53984 0 54096 800
rect 54208 0 54320 800
rect 54432 0 54544 800
rect 54656 0 54768 800
rect 54880 0 54992 800
rect 55104 0 55216 800
rect 55328 0 55440 800
rect 55552 0 55664 800
rect 55776 0 55888 800
rect 56000 0 56112 800
rect 56224 0 56336 800
rect 56448 0 56560 800
rect 56672 0 56784 800
rect 56896 0 57008 800
rect 57120 0 57232 800
rect 57344 0 57456 800
rect 57568 0 57680 800
rect 57792 0 57904 800
rect 58016 0 58128 800
rect 58240 0 58352 800
rect 58464 0 58576 800
rect 58688 0 58800 800
rect 58912 0 59024 800
rect 59136 0 59248 800
rect 59360 0 59472 800
rect 59584 0 59696 800
rect 59808 0 59920 800
rect 60032 0 60144 800
rect 60256 0 60368 800
rect 60480 0 60592 800
rect 60704 0 60816 800
rect 60928 0 61040 800
rect 61152 0 61264 800
rect 61376 0 61488 800
rect 61600 0 61712 800
rect 61824 0 61936 800
rect 62048 0 62160 800
rect 62272 0 62384 800
rect 62496 0 62608 800
rect 62720 0 62832 800
rect 62944 0 63056 800
rect 63168 0 63280 800
rect 63392 0 63504 800
rect 63616 0 63728 800
rect 63840 0 63952 800
rect 64064 0 64176 800
rect 64288 0 64400 800
rect 64512 0 64624 800
rect 64736 0 64848 800
rect 64960 0 65072 800
rect 65184 0 65296 800
rect 65408 0 65520 800
rect 65632 0 65744 800
rect 65856 0 65968 800
rect 66080 0 66192 800
rect 66304 0 66416 800
rect 66528 0 66640 800
rect 66752 0 66864 800
rect 66976 0 67088 800
rect 67200 0 67312 800
rect 67424 0 67536 800
rect 67648 0 67760 800
rect 67872 0 67984 800
rect 68096 0 68208 800
rect 68320 0 68432 800
rect 68544 0 68656 800
rect 68768 0 68880 800
rect 68992 0 69104 800
rect 69216 0 69328 800
rect 69440 0 69552 800
rect 69664 0 69776 800
rect 69888 0 70000 800
rect 70112 0 70224 800
rect 70336 0 70448 800
rect 70560 0 70672 800
rect 70784 0 70896 800
rect 71008 0 71120 800
rect 71232 0 71344 800
rect 71456 0 71568 800
rect 71680 0 71792 800
rect 71904 0 72016 800
rect 72128 0 72240 800
rect 72352 0 72464 800
rect 72576 0 72688 800
rect 72800 0 72912 800
rect 73024 0 73136 800
rect 73248 0 73360 800
rect 73472 0 73584 800
<< obsm2 >>
rect 1932 860 78756 36886
rect 1932 800 6212 860
rect 73644 800 78756 860
<< obsm3 >>
rect 1922 28 78766 36876
<< metal4 >>
rect 10844 3076 11164 36908
rect 20504 3076 20824 36908
rect 30164 3076 30484 36908
rect 39824 3076 40144 36908
rect 49484 3076 49804 36908
rect 59144 3076 59464 36908
rect 68804 3076 69124 36908
rect 78464 3076 78784 36908
<< labels >>
rlabel metal2 s 73024 0 73136 800 6 irq[0]
port 1 nsew signal output
rlabel metal2 s 73248 0 73360 800 6 irq[1]
port 2 nsew signal output
rlabel metal2 s 73472 0 73584 800 6 irq[2]
port 3 nsew signal output
rlabel metal2 s 30016 0 30128 800 6 la_data_in[0]
port 4 nsew signal input
rlabel metal2 s 36736 0 36848 800 6 la_data_in[10]
port 5 nsew signal input
rlabel metal2 s 37408 0 37520 800 6 la_data_in[11]
port 6 nsew signal input
rlabel metal2 s 38080 0 38192 800 6 la_data_in[12]
port 7 nsew signal input
rlabel metal2 s 38752 0 38864 800 6 la_data_in[13]
port 8 nsew signal input
rlabel metal2 s 39424 0 39536 800 6 la_data_in[14]
port 9 nsew signal input
rlabel metal2 s 40096 0 40208 800 6 la_data_in[15]
port 10 nsew signal input
rlabel metal2 s 40768 0 40880 800 6 la_data_in[16]
port 11 nsew signal input
rlabel metal2 s 41440 0 41552 800 6 la_data_in[17]
port 12 nsew signal input
rlabel metal2 s 42112 0 42224 800 6 la_data_in[18]
port 13 nsew signal input
rlabel metal2 s 42784 0 42896 800 6 la_data_in[19]
port 14 nsew signal input
rlabel metal2 s 30688 0 30800 800 6 la_data_in[1]
port 15 nsew signal input
rlabel metal2 s 43456 0 43568 800 6 la_data_in[20]
port 16 nsew signal input
rlabel metal2 s 44128 0 44240 800 6 la_data_in[21]
port 17 nsew signal input
rlabel metal2 s 44800 0 44912 800 6 la_data_in[22]
port 18 nsew signal input
rlabel metal2 s 45472 0 45584 800 6 la_data_in[23]
port 19 nsew signal input
rlabel metal2 s 46144 0 46256 800 6 la_data_in[24]
port 20 nsew signal input
rlabel metal2 s 46816 0 46928 800 6 la_data_in[25]
port 21 nsew signal input
rlabel metal2 s 47488 0 47600 800 6 la_data_in[26]
port 22 nsew signal input
rlabel metal2 s 48160 0 48272 800 6 la_data_in[27]
port 23 nsew signal input
rlabel metal2 s 48832 0 48944 800 6 la_data_in[28]
port 24 nsew signal input
rlabel metal2 s 49504 0 49616 800 6 la_data_in[29]
port 25 nsew signal input
rlabel metal2 s 31360 0 31472 800 6 la_data_in[2]
port 26 nsew signal input
rlabel metal2 s 50176 0 50288 800 6 la_data_in[30]
port 27 nsew signal input
rlabel metal2 s 50848 0 50960 800 6 la_data_in[31]
port 28 nsew signal input
rlabel metal2 s 51520 0 51632 800 6 la_data_in[32]
port 29 nsew signal input
rlabel metal2 s 52192 0 52304 800 6 la_data_in[33]
port 30 nsew signal input
rlabel metal2 s 52864 0 52976 800 6 la_data_in[34]
port 31 nsew signal input
rlabel metal2 s 53536 0 53648 800 6 la_data_in[35]
port 32 nsew signal input
rlabel metal2 s 54208 0 54320 800 6 la_data_in[36]
port 33 nsew signal input
rlabel metal2 s 54880 0 54992 800 6 la_data_in[37]
port 34 nsew signal input
rlabel metal2 s 55552 0 55664 800 6 la_data_in[38]
port 35 nsew signal input
rlabel metal2 s 56224 0 56336 800 6 la_data_in[39]
port 36 nsew signal input
rlabel metal2 s 32032 0 32144 800 6 la_data_in[3]
port 37 nsew signal input
rlabel metal2 s 56896 0 57008 800 6 la_data_in[40]
port 38 nsew signal input
rlabel metal2 s 57568 0 57680 800 6 la_data_in[41]
port 39 nsew signal input
rlabel metal2 s 58240 0 58352 800 6 la_data_in[42]
port 40 nsew signal input
rlabel metal2 s 58912 0 59024 800 6 la_data_in[43]
port 41 nsew signal input
rlabel metal2 s 59584 0 59696 800 6 la_data_in[44]
port 42 nsew signal input
rlabel metal2 s 60256 0 60368 800 6 la_data_in[45]
port 43 nsew signal input
rlabel metal2 s 60928 0 61040 800 6 la_data_in[46]
port 44 nsew signal input
rlabel metal2 s 61600 0 61712 800 6 la_data_in[47]
port 45 nsew signal input
rlabel metal2 s 62272 0 62384 800 6 la_data_in[48]
port 46 nsew signal input
rlabel metal2 s 62944 0 63056 800 6 la_data_in[49]
port 47 nsew signal input
rlabel metal2 s 32704 0 32816 800 6 la_data_in[4]
port 48 nsew signal input
rlabel metal2 s 63616 0 63728 800 6 la_data_in[50]
port 49 nsew signal input
rlabel metal2 s 64288 0 64400 800 6 la_data_in[51]
port 50 nsew signal input
rlabel metal2 s 64960 0 65072 800 6 la_data_in[52]
port 51 nsew signal input
rlabel metal2 s 65632 0 65744 800 6 la_data_in[53]
port 52 nsew signal input
rlabel metal2 s 66304 0 66416 800 6 la_data_in[54]
port 53 nsew signal input
rlabel metal2 s 66976 0 67088 800 6 la_data_in[55]
port 54 nsew signal input
rlabel metal2 s 67648 0 67760 800 6 la_data_in[56]
port 55 nsew signal input
rlabel metal2 s 68320 0 68432 800 6 la_data_in[57]
port 56 nsew signal input
rlabel metal2 s 68992 0 69104 800 6 la_data_in[58]
port 57 nsew signal input
rlabel metal2 s 69664 0 69776 800 6 la_data_in[59]
port 58 nsew signal input
rlabel metal2 s 33376 0 33488 800 6 la_data_in[5]
port 59 nsew signal input
rlabel metal2 s 70336 0 70448 800 6 la_data_in[60]
port 60 nsew signal input
rlabel metal2 s 71008 0 71120 800 6 la_data_in[61]
port 61 nsew signal input
rlabel metal2 s 71680 0 71792 800 6 la_data_in[62]
port 62 nsew signal input
rlabel metal2 s 72352 0 72464 800 6 la_data_in[63]
port 63 nsew signal input
rlabel metal2 s 34048 0 34160 800 6 la_data_in[6]
port 64 nsew signal input
rlabel metal2 s 34720 0 34832 800 6 la_data_in[7]
port 65 nsew signal input
rlabel metal2 s 35392 0 35504 800 6 la_data_in[8]
port 66 nsew signal input
rlabel metal2 s 36064 0 36176 800 6 la_data_in[9]
port 67 nsew signal input
rlabel metal2 s 30240 0 30352 800 6 la_data_out[0]
port 68 nsew signal output
rlabel metal2 s 36960 0 37072 800 6 la_data_out[10]
port 69 nsew signal output
rlabel metal2 s 37632 0 37744 800 6 la_data_out[11]
port 70 nsew signal output
rlabel metal2 s 38304 0 38416 800 6 la_data_out[12]
port 71 nsew signal output
rlabel metal2 s 38976 0 39088 800 6 la_data_out[13]
port 72 nsew signal output
rlabel metal2 s 39648 0 39760 800 6 la_data_out[14]
port 73 nsew signal output
rlabel metal2 s 40320 0 40432 800 6 la_data_out[15]
port 74 nsew signal output
rlabel metal2 s 40992 0 41104 800 6 la_data_out[16]
port 75 nsew signal output
rlabel metal2 s 41664 0 41776 800 6 la_data_out[17]
port 76 nsew signal output
rlabel metal2 s 42336 0 42448 800 6 la_data_out[18]
port 77 nsew signal output
rlabel metal2 s 43008 0 43120 800 6 la_data_out[19]
port 78 nsew signal output
rlabel metal2 s 30912 0 31024 800 6 la_data_out[1]
port 79 nsew signal output
rlabel metal2 s 43680 0 43792 800 6 la_data_out[20]
port 80 nsew signal output
rlabel metal2 s 44352 0 44464 800 6 la_data_out[21]
port 81 nsew signal output
rlabel metal2 s 45024 0 45136 800 6 la_data_out[22]
port 82 nsew signal output
rlabel metal2 s 45696 0 45808 800 6 la_data_out[23]
port 83 nsew signal output
rlabel metal2 s 46368 0 46480 800 6 la_data_out[24]
port 84 nsew signal output
rlabel metal2 s 47040 0 47152 800 6 la_data_out[25]
port 85 nsew signal output
rlabel metal2 s 47712 0 47824 800 6 la_data_out[26]
port 86 nsew signal output
rlabel metal2 s 48384 0 48496 800 6 la_data_out[27]
port 87 nsew signal output
rlabel metal2 s 49056 0 49168 800 6 la_data_out[28]
port 88 nsew signal output
rlabel metal2 s 49728 0 49840 800 6 la_data_out[29]
port 89 nsew signal output
rlabel metal2 s 31584 0 31696 800 6 la_data_out[2]
port 90 nsew signal output
rlabel metal2 s 50400 0 50512 800 6 la_data_out[30]
port 91 nsew signal output
rlabel metal2 s 51072 0 51184 800 6 la_data_out[31]
port 92 nsew signal output
rlabel metal2 s 51744 0 51856 800 6 la_data_out[32]
port 93 nsew signal output
rlabel metal2 s 52416 0 52528 800 6 la_data_out[33]
port 94 nsew signal output
rlabel metal2 s 53088 0 53200 800 6 la_data_out[34]
port 95 nsew signal output
rlabel metal2 s 53760 0 53872 800 6 la_data_out[35]
port 96 nsew signal output
rlabel metal2 s 54432 0 54544 800 6 la_data_out[36]
port 97 nsew signal output
rlabel metal2 s 55104 0 55216 800 6 la_data_out[37]
port 98 nsew signal output
rlabel metal2 s 55776 0 55888 800 6 la_data_out[38]
port 99 nsew signal output
rlabel metal2 s 56448 0 56560 800 6 la_data_out[39]
port 100 nsew signal output
rlabel metal2 s 32256 0 32368 800 6 la_data_out[3]
port 101 nsew signal output
rlabel metal2 s 57120 0 57232 800 6 la_data_out[40]
port 102 nsew signal output
rlabel metal2 s 57792 0 57904 800 6 la_data_out[41]
port 103 nsew signal output
rlabel metal2 s 58464 0 58576 800 6 la_data_out[42]
port 104 nsew signal output
rlabel metal2 s 59136 0 59248 800 6 la_data_out[43]
port 105 nsew signal output
rlabel metal2 s 59808 0 59920 800 6 la_data_out[44]
port 106 nsew signal output
rlabel metal2 s 60480 0 60592 800 6 la_data_out[45]
port 107 nsew signal output
rlabel metal2 s 61152 0 61264 800 6 la_data_out[46]
port 108 nsew signal output
rlabel metal2 s 61824 0 61936 800 6 la_data_out[47]
port 109 nsew signal output
rlabel metal2 s 62496 0 62608 800 6 la_data_out[48]
port 110 nsew signal output
rlabel metal2 s 63168 0 63280 800 6 la_data_out[49]
port 111 nsew signal output
rlabel metal2 s 32928 0 33040 800 6 la_data_out[4]
port 112 nsew signal output
rlabel metal2 s 63840 0 63952 800 6 la_data_out[50]
port 113 nsew signal output
rlabel metal2 s 64512 0 64624 800 6 la_data_out[51]
port 114 nsew signal output
rlabel metal2 s 65184 0 65296 800 6 la_data_out[52]
port 115 nsew signal output
rlabel metal2 s 65856 0 65968 800 6 la_data_out[53]
port 116 nsew signal output
rlabel metal2 s 66528 0 66640 800 6 la_data_out[54]
port 117 nsew signal output
rlabel metal2 s 67200 0 67312 800 6 la_data_out[55]
port 118 nsew signal output
rlabel metal2 s 67872 0 67984 800 6 la_data_out[56]
port 119 nsew signal output
rlabel metal2 s 68544 0 68656 800 6 la_data_out[57]
port 120 nsew signal output
rlabel metal2 s 69216 0 69328 800 6 la_data_out[58]
port 121 nsew signal output
rlabel metal2 s 69888 0 70000 800 6 la_data_out[59]
port 122 nsew signal output
rlabel metal2 s 33600 0 33712 800 6 la_data_out[5]
port 123 nsew signal output
rlabel metal2 s 70560 0 70672 800 6 la_data_out[60]
port 124 nsew signal output
rlabel metal2 s 71232 0 71344 800 6 la_data_out[61]
port 125 nsew signal output
rlabel metal2 s 71904 0 72016 800 6 la_data_out[62]
port 126 nsew signal output
rlabel metal2 s 72576 0 72688 800 6 la_data_out[63]
port 127 nsew signal output
rlabel metal2 s 34272 0 34384 800 6 la_data_out[6]
port 128 nsew signal output
rlabel metal2 s 34944 0 35056 800 6 la_data_out[7]
port 129 nsew signal output
rlabel metal2 s 35616 0 35728 800 6 la_data_out[8]
port 130 nsew signal output
rlabel metal2 s 36288 0 36400 800 6 la_data_out[9]
port 131 nsew signal output
rlabel metal2 s 30464 0 30576 800 6 la_oenb[0]
port 132 nsew signal input
rlabel metal2 s 37184 0 37296 800 6 la_oenb[10]
port 133 nsew signal input
rlabel metal2 s 37856 0 37968 800 6 la_oenb[11]
port 134 nsew signal input
rlabel metal2 s 38528 0 38640 800 6 la_oenb[12]
port 135 nsew signal input
rlabel metal2 s 39200 0 39312 800 6 la_oenb[13]
port 136 nsew signal input
rlabel metal2 s 39872 0 39984 800 6 la_oenb[14]
port 137 nsew signal input
rlabel metal2 s 40544 0 40656 800 6 la_oenb[15]
port 138 nsew signal input
rlabel metal2 s 41216 0 41328 800 6 la_oenb[16]
port 139 nsew signal input
rlabel metal2 s 41888 0 42000 800 6 la_oenb[17]
port 140 nsew signal input
rlabel metal2 s 42560 0 42672 800 6 la_oenb[18]
port 141 nsew signal input
rlabel metal2 s 43232 0 43344 800 6 la_oenb[19]
port 142 nsew signal input
rlabel metal2 s 31136 0 31248 800 6 la_oenb[1]
port 143 nsew signal input
rlabel metal2 s 43904 0 44016 800 6 la_oenb[20]
port 144 nsew signal input
rlabel metal2 s 44576 0 44688 800 6 la_oenb[21]
port 145 nsew signal input
rlabel metal2 s 45248 0 45360 800 6 la_oenb[22]
port 146 nsew signal input
rlabel metal2 s 45920 0 46032 800 6 la_oenb[23]
port 147 nsew signal input
rlabel metal2 s 46592 0 46704 800 6 la_oenb[24]
port 148 nsew signal input
rlabel metal2 s 47264 0 47376 800 6 la_oenb[25]
port 149 nsew signal input
rlabel metal2 s 47936 0 48048 800 6 la_oenb[26]
port 150 nsew signal input
rlabel metal2 s 48608 0 48720 800 6 la_oenb[27]
port 151 nsew signal input
rlabel metal2 s 49280 0 49392 800 6 la_oenb[28]
port 152 nsew signal input
rlabel metal2 s 49952 0 50064 800 6 la_oenb[29]
port 153 nsew signal input
rlabel metal2 s 31808 0 31920 800 6 la_oenb[2]
port 154 nsew signal input
rlabel metal2 s 50624 0 50736 800 6 la_oenb[30]
port 155 nsew signal input
rlabel metal2 s 51296 0 51408 800 6 la_oenb[31]
port 156 nsew signal input
rlabel metal2 s 51968 0 52080 800 6 la_oenb[32]
port 157 nsew signal input
rlabel metal2 s 52640 0 52752 800 6 la_oenb[33]
port 158 nsew signal input
rlabel metal2 s 53312 0 53424 800 6 la_oenb[34]
port 159 nsew signal input
rlabel metal2 s 53984 0 54096 800 6 la_oenb[35]
port 160 nsew signal input
rlabel metal2 s 54656 0 54768 800 6 la_oenb[36]
port 161 nsew signal input
rlabel metal2 s 55328 0 55440 800 6 la_oenb[37]
port 162 nsew signal input
rlabel metal2 s 56000 0 56112 800 6 la_oenb[38]
port 163 nsew signal input
rlabel metal2 s 56672 0 56784 800 6 la_oenb[39]
port 164 nsew signal input
rlabel metal2 s 32480 0 32592 800 6 la_oenb[3]
port 165 nsew signal input
rlabel metal2 s 57344 0 57456 800 6 la_oenb[40]
port 166 nsew signal input
rlabel metal2 s 58016 0 58128 800 6 la_oenb[41]
port 167 nsew signal input
rlabel metal2 s 58688 0 58800 800 6 la_oenb[42]
port 168 nsew signal input
rlabel metal2 s 59360 0 59472 800 6 la_oenb[43]
port 169 nsew signal input
rlabel metal2 s 60032 0 60144 800 6 la_oenb[44]
port 170 nsew signal input
rlabel metal2 s 60704 0 60816 800 6 la_oenb[45]
port 171 nsew signal input
rlabel metal2 s 61376 0 61488 800 6 la_oenb[46]
port 172 nsew signal input
rlabel metal2 s 62048 0 62160 800 6 la_oenb[47]
port 173 nsew signal input
rlabel metal2 s 62720 0 62832 800 6 la_oenb[48]
port 174 nsew signal input
rlabel metal2 s 63392 0 63504 800 6 la_oenb[49]
port 175 nsew signal input
rlabel metal2 s 33152 0 33264 800 6 la_oenb[4]
port 176 nsew signal input
rlabel metal2 s 64064 0 64176 800 6 la_oenb[50]
port 177 nsew signal input
rlabel metal2 s 64736 0 64848 800 6 la_oenb[51]
port 178 nsew signal input
rlabel metal2 s 65408 0 65520 800 6 la_oenb[52]
port 179 nsew signal input
rlabel metal2 s 66080 0 66192 800 6 la_oenb[53]
port 180 nsew signal input
rlabel metal2 s 66752 0 66864 800 6 la_oenb[54]
port 181 nsew signal input
rlabel metal2 s 67424 0 67536 800 6 la_oenb[55]
port 182 nsew signal input
rlabel metal2 s 68096 0 68208 800 6 la_oenb[56]
port 183 nsew signal input
rlabel metal2 s 68768 0 68880 800 6 la_oenb[57]
port 184 nsew signal input
rlabel metal2 s 69440 0 69552 800 6 la_oenb[58]
port 185 nsew signal input
rlabel metal2 s 70112 0 70224 800 6 la_oenb[59]
port 186 nsew signal input
rlabel metal2 s 33824 0 33936 800 6 la_oenb[5]
port 187 nsew signal input
rlabel metal2 s 70784 0 70896 800 6 la_oenb[60]
port 188 nsew signal input
rlabel metal2 s 71456 0 71568 800 6 la_oenb[61]
port 189 nsew signal input
rlabel metal2 s 72128 0 72240 800 6 la_oenb[62]
port 190 nsew signal input
rlabel metal2 s 72800 0 72912 800 6 la_oenb[63]
port 191 nsew signal input
rlabel metal2 s 34496 0 34608 800 6 la_oenb[6]
port 192 nsew signal input
rlabel metal2 s 35168 0 35280 800 6 la_oenb[7]
port 193 nsew signal input
rlabel metal2 s 35840 0 35952 800 6 la_oenb[8]
port 194 nsew signal input
rlabel metal2 s 36512 0 36624 800 6 la_oenb[9]
port 195 nsew signal input
rlabel metal4 s 10844 3076 11164 36908 6 vdd
port 196 nsew power bidirectional
rlabel metal4 s 30164 3076 30484 36908 6 vdd
port 196 nsew power bidirectional
rlabel metal4 s 49484 3076 49804 36908 6 vdd
port 196 nsew power bidirectional
rlabel metal4 s 68804 3076 69124 36908 6 vdd
port 196 nsew power bidirectional
rlabel metal4 s 20504 3076 20824 36908 6 vss
port 197 nsew ground bidirectional
rlabel metal4 s 39824 3076 40144 36908 6 vss
port 197 nsew ground bidirectional
rlabel metal4 s 59144 3076 59464 36908 6 vss
port 197 nsew ground bidirectional
rlabel metal4 s 78464 3076 78784 36908 6 vss
port 197 nsew ground bidirectional
rlabel metal2 s 6272 0 6384 800 6 wb_clk_i
port 198 nsew signal input
rlabel metal2 s 6496 0 6608 800 6 wb_rst_i
port 199 nsew signal input
rlabel metal2 s 6720 0 6832 800 6 wbs_ack_o
port 200 nsew signal output
rlabel metal2 s 7616 0 7728 800 6 wbs_adr_i[0]
port 201 nsew signal input
rlabel metal2 s 15232 0 15344 800 6 wbs_adr_i[10]
port 202 nsew signal input
rlabel metal2 s 15904 0 16016 800 6 wbs_adr_i[11]
port 203 nsew signal input
rlabel metal2 s 16576 0 16688 800 6 wbs_adr_i[12]
port 204 nsew signal input
rlabel metal2 s 17248 0 17360 800 6 wbs_adr_i[13]
port 205 nsew signal input
rlabel metal2 s 17920 0 18032 800 6 wbs_adr_i[14]
port 206 nsew signal input
rlabel metal2 s 18592 0 18704 800 6 wbs_adr_i[15]
port 207 nsew signal input
rlabel metal2 s 19264 0 19376 800 6 wbs_adr_i[16]
port 208 nsew signal input
rlabel metal2 s 19936 0 20048 800 6 wbs_adr_i[17]
port 209 nsew signal input
rlabel metal2 s 20608 0 20720 800 6 wbs_adr_i[18]
port 210 nsew signal input
rlabel metal2 s 21280 0 21392 800 6 wbs_adr_i[19]
port 211 nsew signal input
rlabel metal2 s 8512 0 8624 800 6 wbs_adr_i[1]
port 212 nsew signal input
rlabel metal2 s 21952 0 22064 800 6 wbs_adr_i[20]
port 213 nsew signal input
rlabel metal2 s 22624 0 22736 800 6 wbs_adr_i[21]
port 214 nsew signal input
rlabel metal2 s 23296 0 23408 800 6 wbs_adr_i[22]
port 215 nsew signal input
rlabel metal2 s 23968 0 24080 800 6 wbs_adr_i[23]
port 216 nsew signal input
rlabel metal2 s 24640 0 24752 800 6 wbs_adr_i[24]
port 217 nsew signal input
rlabel metal2 s 25312 0 25424 800 6 wbs_adr_i[25]
port 218 nsew signal input
rlabel metal2 s 25984 0 26096 800 6 wbs_adr_i[26]
port 219 nsew signal input
rlabel metal2 s 26656 0 26768 800 6 wbs_adr_i[27]
port 220 nsew signal input
rlabel metal2 s 27328 0 27440 800 6 wbs_adr_i[28]
port 221 nsew signal input
rlabel metal2 s 28000 0 28112 800 6 wbs_adr_i[29]
port 222 nsew signal input
rlabel metal2 s 9408 0 9520 800 6 wbs_adr_i[2]
port 223 nsew signal input
rlabel metal2 s 28672 0 28784 800 6 wbs_adr_i[30]
port 224 nsew signal input
rlabel metal2 s 29344 0 29456 800 6 wbs_adr_i[31]
port 225 nsew signal input
rlabel metal2 s 10304 0 10416 800 6 wbs_adr_i[3]
port 226 nsew signal input
rlabel metal2 s 11200 0 11312 800 6 wbs_adr_i[4]
port 227 nsew signal input
rlabel metal2 s 11872 0 11984 800 6 wbs_adr_i[5]
port 228 nsew signal input
rlabel metal2 s 12544 0 12656 800 6 wbs_adr_i[6]
port 229 nsew signal input
rlabel metal2 s 13216 0 13328 800 6 wbs_adr_i[7]
port 230 nsew signal input
rlabel metal2 s 13888 0 14000 800 6 wbs_adr_i[8]
port 231 nsew signal input
rlabel metal2 s 14560 0 14672 800 6 wbs_adr_i[9]
port 232 nsew signal input
rlabel metal2 s 6944 0 7056 800 6 wbs_cyc_i
port 233 nsew signal input
rlabel metal2 s 7840 0 7952 800 6 wbs_dat_i[0]
port 234 nsew signal input
rlabel metal2 s 15456 0 15568 800 6 wbs_dat_i[10]
port 235 nsew signal input
rlabel metal2 s 16128 0 16240 800 6 wbs_dat_i[11]
port 236 nsew signal input
rlabel metal2 s 16800 0 16912 800 6 wbs_dat_i[12]
port 237 nsew signal input
rlabel metal2 s 17472 0 17584 800 6 wbs_dat_i[13]
port 238 nsew signal input
rlabel metal2 s 18144 0 18256 800 6 wbs_dat_i[14]
port 239 nsew signal input
rlabel metal2 s 18816 0 18928 800 6 wbs_dat_i[15]
port 240 nsew signal input
rlabel metal2 s 19488 0 19600 800 6 wbs_dat_i[16]
port 241 nsew signal input
rlabel metal2 s 20160 0 20272 800 6 wbs_dat_i[17]
port 242 nsew signal input
rlabel metal2 s 20832 0 20944 800 6 wbs_dat_i[18]
port 243 nsew signal input
rlabel metal2 s 21504 0 21616 800 6 wbs_dat_i[19]
port 244 nsew signal input
rlabel metal2 s 8736 0 8848 800 6 wbs_dat_i[1]
port 245 nsew signal input
rlabel metal2 s 22176 0 22288 800 6 wbs_dat_i[20]
port 246 nsew signal input
rlabel metal2 s 22848 0 22960 800 6 wbs_dat_i[21]
port 247 nsew signal input
rlabel metal2 s 23520 0 23632 800 6 wbs_dat_i[22]
port 248 nsew signal input
rlabel metal2 s 24192 0 24304 800 6 wbs_dat_i[23]
port 249 nsew signal input
rlabel metal2 s 24864 0 24976 800 6 wbs_dat_i[24]
port 250 nsew signal input
rlabel metal2 s 25536 0 25648 800 6 wbs_dat_i[25]
port 251 nsew signal input
rlabel metal2 s 26208 0 26320 800 6 wbs_dat_i[26]
port 252 nsew signal input
rlabel metal2 s 26880 0 26992 800 6 wbs_dat_i[27]
port 253 nsew signal input
rlabel metal2 s 27552 0 27664 800 6 wbs_dat_i[28]
port 254 nsew signal input
rlabel metal2 s 28224 0 28336 800 6 wbs_dat_i[29]
port 255 nsew signal input
rlabel metal2 s 9632 0 9744 800 6 wbs_dat_i[2]
port 256 nsew signal input
rlabel metal2 s 28896 0 29008 800 6 wbs_dat_i[30]
port 257 nsew signal input
rlabel metal2 s 29568 0 29680 800 6 wbs_dat_i[31]
port 258 nsew signal input
rlabel metal2 s 10528 0 10640 800 6 wbs_dat_i[3]
port 259 nsew signal input
rlabel metal2 s 11424 0 11536 800 6 wbs_dat_i[4]
port 260 nsew signal input
rlabel metal2 s 12096 0 12208 800 6 wbs_dat_i[5]
port 261 nsew signal input
rlabel metal2 s 12768 0 12880 800 6 wbs_dat_i[6]
port 262 nsew signal input
rlabel metal2 s 13440 0 13552 800 6 wbs_dat_i[7]
port 263 nsew signal input
rlabel metal2 s 14112 0 14224 800 6 wbs_dat_i[8]
port 264 nsew signal input
rlabel metal2 s 14784 0 14896 800 6 wbs_dat_i[9]
port 265 nsew signal input
rlabel metal2 s 8064 0 8176 800 6 wbs_dat_o[0]
port 266 nsew signal output
rlabel metal2 s 15680 0 15792 800 6 wbs_dat_o[10]
port 267 nsew signal output
rlabel metal2 s 16352 0 16464 800 6 wbs_dat_o[11]
port 268 nsew signal output
rlabel metal2 s 17024 0 17136 800 6 wbs_dat_o[12]
port 269 nsew signal output
rlabel metal2 s 17696 0 17808 800 6 wbs_dat_o[13]
port 270 nsew signal output
rlabel metal2 s 18368 0 18480 800 6 wbs_dat_o[14]
port 271 nsew signal output
rlabel metal2 s 19040 0 19152 800 6 wbs_dat_o[15]
port 272 nsew signal output
rlabel metal2 s 19712 0 19824 800 6 wbs_dat_o[16]
port 273 nsew signal output
rlabel metal2 s 20384 0 20496 800 6 wbs_dat_o[17]
port 274 nsew signal output
rlabel metal2 s 21056 0 21168 800 6 wbs_dat_o[18]
port 275 nsew signal output
rlabel metal2 s 21728 0 21840 800 6 wbs_dat_o[19]
port 276 nsew signal output
rlabel metal2 s 8960 0 9072 800 6 wbs_dat_o[1]
port 277 nsew signal output
rlabel metal2 s 22400 0 22512 800 6 wbs_dat_o[20]
port 278 nsew signal output
rlabel metal2 s 23072 0 23184 800 6 wbs_dat_o[21]
port 279 nsew signal output
rlabel metal2 s 23744 0 23856 800 6 wbs_dat_o[22]
port 280 nsew signal output
rlabel metal2 s 24416 0 24528 800 6 wbs_dat_o[23]
port 281 nsew signal output
rlabel metal2 s 25088 0 25200 800 6 wbs_dat_o[24]
port 282 nsew signal output
rlabel metal2 s 25760 0 25872 800 6 wbs_dat_o[25]
port 283 nsew signal output
rlabel metal2 s 26432 0 26544 800 6 wbs_dat_o[26]
port 284 nsew signal output
rlabel metal2 s 27104 0 27216 800 6 wbs_dat_o[27]
port 285 nsew signal output
rlabel metal2 s 27776 0 27888 800 6 wbs_dat_o[28]
port 286 nsew signal output
rlabel metal2 s 28448 0 28560 800 6 wbs_dat_o[29]
port 287 nsew signal output
rlabel metal2 s 9856 0 9968 800 6 wbs_dat_o[2]
port 288 nsew signal output
rlabel metal2 s 29120 0 29232 800 6 wbs_dat_o[30]
port 289 nsew signal output
rlabel metal2 s 29792 0 29904 800 6 wbs_dat_o[31]
port 290 nsew signal output
rlabel metal2 s 10752 0 10864 800 6 wbs_dat_o[3]
port 291 nsew signal output
rlabel metal2 s 11648 0 11760 800 6 wbs_dat_o[4]
port 292 nsew signal output
rlabel metal2 s 12320 0 12432 800 6 wbs_dat_o[5]
port 293 nsew signal output
rlabel metal2 s 12992 0 13104 800 6 wbs_dat_o[6]
port 294 nsew signal output
rlabel metal2 s 13664 0 13776 800 6 wbs_dat_o[7]
port 295 nsew signal output
rlabel metal2 s 14336 0 14448 800 6 wbs_dat_o[8]
port 296 nsew signal output
rlabel metal2 s 15008 0 15120 800 6 wbs_dat_o[9]
port 297 nsew signal output
rlabel metal2 s 8288 0 8400 800 6 wbs_sel_i[0]
port 298 nsew signal input
rlabel metal2 s 9184 0 9296 800 6 wbs_sel_i[1]
port 299 nsew signal input
rlabel metal2 s 10080 0 10192 800 6 wbs_sel_i[2]
port 300 nsew signal input
rlabel metal2 s 10976 0 11088 800 6 wbs_sel_i[3]
port 301 nsew signal input
rlabel metal2 s 7168 0 7280 800 6 wbs_stb_i
port 302 nsew signal input
rlabel metal2 s 7392 0 7504 800 6 wbs_we_i
port 303 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1250738
string GDS_FILE /home/ishi-kai/test/caravel_user_project-gfmpw-1c/openlane/user_proj_example/runs/23_11_10_17_53/results/signoff/user_proj_example.magic.gds
string GDS_START 207420
<< end >>

