* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD GND A6 Q7
X0 Q7.t8 A6.t0 VDD.t11 VDD.t10 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.6u
X1 Q7.t0 A6.t1 GND.t5 GND.t4 nfet_06v0 ad=0.876p pd=3.86u as=0.312p ps=1.72u w=1.2u l=0.6u
X2 Q7.t7 A6.t2 VDD.t9 VDD.t8 pfet_06v0 ad=0.312p pd=1.72u as=0.924p ps=3.94u w=1.2u l=0.6u
X3 Q7.t6 A6.t3 VDD.t7 VDD.t6 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.6u
X4 GND.t3 A6.t4 Q7.t1 GND.t2 nfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.6u
X5 VDD.t5 A6.t5 Q7.t5 VDD.t4 pfet_06v0 ad=0.924p pd=3.94u as=0.312p ps=1.72u w=1.2u l=0.6u
X6 Q7.t2 A6.t6 GND.t1 GND.t0 nfet_06v0 ad=0.312p pd=1.72u as=0.876p ps=3.86u w=1.2u l=0.6u
X7 VDD.t3 A6.t7 Q7.t4 VDD.t2 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.6u
X8 VDD.t1 A6.t8 Q7.t3 VDD.t0 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.6u
R0 A6.n0 A6.t5 21.2634
R1 A6.n7 A6.t2 21.2622
R2 A6.n6 A6.t8 21.2622
R3 A6.n5 A6.t3 21.2622
R4 A6.n3 A6.t7 21.2622
R5 A6.n1 A6.t0 21.2622
R6 A6.n4 A6.t6 21.1405
R7 A6.n2 A6.t4 21.1405
R8 A6.n0 A6.t1 21.1405
R9 A6 A6.n7 0.813264
R10 A6.n6 A6.n5 0.0279659
R11 A6.n7 A6.n6 0.0279659
R12 A6.n1 A6.n0 0.0267398
R13 A6.n3 A6.n2 0.0267398
R14 A6.n5 A6.n4 0.0267398
R15 A6.n2 A6.n1 0.00172616
R16 A6.n4 A6.n3 0.00172616
R17 VDD.n0 VDD.t8 614.89
R18 VDD.t10 VDD.t4 434.11
R19 VDD.t2 VDD.t10 434.11
R20 VDD.t6 VDD.t2 434.11
R21 VDD.t0 VDD.t6 434.11
R22 VDD.t8 VDD.t0 434.11
R23 VDD.n2 VDD.t5 10.8957
R24 VDD.n4 VDD.n3 7.17866
R25 VDD.n2 VDD.n1 7.17866
R26 VDD.n0 VDD.t9 5.81367
R27 VDD.n5 VDD.n4 5.0675
R28 VDD.n3 VDD.t7 1.51717
R29 VDD.n3 VDD.t1 1.51717
R30 VDD.n1 VDD.t11 1.51717
R31 VDD.n1 VDD.t3 1.51717
R32 VDD VDD.n5 0.783131
R33 VDD.n4 VDD.n2 0.5045
R34 VDD.n5 VDD.n0 0.0213929
R35 Q7.n6 Q7.t0 14.9587
R36 Q7.n6 Q7.n5 12.7178
R37 Q7.n2 Q7.n0 12.1827
R38 Q7.n2 Q7.n1 11.6787
R39 Q7.n4 Q7.n3 11.6787
R40 Q7 Q7.n7 10.4064
R41 Q7.n0 Q7.t3 1.51717
R42 Q7.n0 Q7.t7 1.51717
R43 Q7.n1 Q7.t4 1.51717
R44 Q7.n1 Q7.t6 1.51717
R45 Q7.n3 Q7.t5 1.51717
R46 Q7.n3 Q7.t8 1.51717
R47 Q7.n5 Q7.t1 1.3655
R48 Q7.n5 Q7.t2 1.3655
R49 Q7.n7 Q7.n4 1.265
R50 Q7.n7 Q7.n6 0.91263
R51 Q7.n4 Q7.n2 0.5045
R52 GND.n0 GND.t4 13396.6
R53 GND.n0 GND.t0 430.147
R54 GND.t4 GND.t2 314.88
R55 GND.t2 GND.t0 314.88
R56 GND.n3 GND.n2 12.6805
R57 GND.n1 GND.t1 5.94194
R58 GND.n1 GND.n0 5.26194
R59 GND.n2 GND.t5 1.3655
R60 GND.n2 GND.t3 1.3655
R61 GND GND.n3 0.431818
R62 GND.n3 GND.n1 0.0225909
C0 A6 VDD 1.36314f
C1 Q7 VDD 0.795268f
C2 A6 Q7 0.821901f
C3 Q7 GND 3.302f
C4 A6 GND 4.64255f
C5 VDD GND 5.22904f
.ends

