* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VSS OUT VINP VDD VINN IB
X0 a_61329_n6784.t11 VINN.t0 dw_60815_n7004.t21 dw_60815_n7004.t25 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X1 OUT.t39 IB.t0 VDD.t45 VDD.t44 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X2 OUT.t38 IB.t1 VDD.t43 VDD.t42 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X3 VSS.t50 a_66329_n6784.t9 OUT.t15 VSS.t49 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X4 a_66329_n6784.t0 a_55035_n6784.t3 a_79287_n10784.t1 VSS.t0 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X5 OUT.t14 a_66329_n6784.t10 VSS.t48 VSS.t47 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X6 a_79287_n10784.t1 a_55035_n6784.t4 a_66329_n6784.t4 VSS.t2 nfet_06v0 ad=0.91p pd=4.02u as=2.555p ps=8.46u w=3.5u l=0.7u
X7 dw_60815_n7004.t9 VINP.t0 a_66329_n6784.t3 dw_60815_n7004.t8 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X8 OUT.t37 IB.t2 VDD.t41 VDD.t40 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X9 a_66329_n6784.t3 VINP.t1 dw_60815_n7004.t4 dw_60815_n7004.t3 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X10 VSS.t10 a_55043_n10784 a_55043_n10784 VSS.t9 nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X11 dw_60815_n7004.t1 VINP.t2 a_66329_n6784.t1 dw_60815_n7004.t0 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X12 OUT.t36 IB.t3 VDD.t39 VDD.t38 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X13 a_66329_n6784.t7 a_55035_n6784.t5 a_79287_n10784.t0 VSS.t4 nfet_06v0 ad=2.555p pd=8.46u as=0.91p ps=4.02u w=3.5u l=0.7u
X14 dw_60815_n7004.t6 VINP.t3 a_66329_n6784.t5 dw_60815_n7004.t5 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X15 a_66329_n6784.t8 a_61329_n6784.t12 VSS.t8 VSS.t7 nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X16 dw_60815_n7004.t28 IB.t4 VDD.t37 VDD.t36 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X17 a_61329_n6784.t10 VINN.t1 dw_60815_n7004.t15 dw_60815_n7004.t24 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X18 dw_60815_n7004.t13 VINN.t2 a_61329_n6784.t9 dw_60815_n7004.t23 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X19 dw_60815_n7004.t11 VINN.t3 a_61329_n6784.t8 dw_60815_n7004.t22 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X20 OUT.t19 a_66329_n6784.t11 VSS.t46 VSS.t45 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X21 VDD.t35 IB.t5 a_55035_n6784.t2 VDD.t34 pfet_06v0 ad=5.39p pd=15.539999u as=5.39p ps=15.539999u w=7u l=0.7u
X22 VSS.t44 a_66329_n6784.t12 OUT.t10 VSS.t43 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X23 VSS.t42 a_66329_n6784.t13 OUT.t4 VSS.t41 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X24 dw_60815_n7004.t21 VINN.t4 a_61329_n6784.t7 dw_60815_n7004.t20 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X25 OUT.t35 IB.t6 VDD.t33 VDD.t32 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X26 VDD.t31 IB.t7 OUT.t34 VDD.t30 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X27 OUT.t13 a_66329_n6784.t14 VSS.t40 VSS.t39 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X28 OUT.t7 a_66329_n6784.t15 VSS.t38 VSS.t37 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X29 VDD.t29 IB.t8 OUT.t33 VDD.t28 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X30 VSS.t6 a_61329_n6784.t0 a_61329_n6784.t1 VSS.t5 nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X31 VSS.t36 a_66329_n6784.t16 OUT.t9 VSS.t35 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X32 VDD.t27 IB.t9 OUT.t32 VDD.t26 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X33 VDD.t25 IB.t10 OUT.t31 VDD.t24 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X34 OUT.t5 a_66329_n6784.t17 VSS.t34 VSS.t33 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X35 VSS.t32 a_66329_n6784.t18 OUT.t3 VSS.t31 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X36 dw_60815_n7004.t27 VINP.t4 a_66329_n6784.t2 dw_60815_n7004.t26 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X37 OUT.t30 IB.t11 VDD.t3 VDD.t2 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X38 VSS.t30 a_66329_n6784.t19 OUT.t12 VSS.t29 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X39 VSS.t28 a_66329_n6784.t20 OUT.t11 VSS.t27 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X40 OUT.t2 a_66329_n6784.t21 VSS.t26 VSS.t25 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X41 a_66329_n6784.t5 VINP.t5 dw_60815_n7004.t31 dw_60815_n7004.t30 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X42 VDD.t23 IB.t12 OUT.t29 VDD.t22 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X43 a_66329_n6784.t1 VINP.t6 dw_60815_n7004.t9 dw_60815_n7004.t32 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X44 VDD.t21 IB.t13 OUT.t28 VDD.t20 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X46 dw_60815_n7004.t19 VINN.t5 a_61329_n6784.t6 dw_60815_n7004.t18 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X47 a_79287_n10784.t0 a_55035_n6784.t6 a_66329_n6784.t0 VSS.t1 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X48 a_61329_n6784.t5 VINN.t6 dw_60815_n7004.t17 dw_60815_n7004.t16 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X49 dw_60815_n7004.t4 VINP.t7 a_66329_n6784.t6 dw_60815_n7004.t7 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X50 OUT.t18 a_66329_n6784.t22 VSS.t24 VSS.t23 nfet_06v0 ad=0.91p pd=4.02u as=2.555p ps=8.46u w=3.5u l=0.7u
X51 a_61329_n6784.t4 VINN.t7 dw_60815_n7004.t13 dw_60815_n7004.t12 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X52 VDD.t5 IB.t14 OUT.t27 VDD.t4 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X53 OUT.t26 IB.t15 VDD.t19 VDD.t18 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X54 dw_60815_n7004.t15 VINN.t8 a_61329_n6784.t3 dw_60815_n7004.t14 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X55 OUT.t25 IB.t16 VDD.t17 VDD.t16 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X56 VDD.t9 IB.t17 OUT.t24 VDD.t8 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X57 VSS.t22 a_66329_n6784.t23 OUT.t0 VSS.t21 nfet_06v0 ad=2.555p pd=8.46u as=0.91p ps=4.02u w=3.5u l=0.7u
X58 a_66329_n6784.t2 VINP.t8 dw_60815_n7004.t1 dw_60815_n7004.t2 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X59 OUT.t23 IB.t18 VDD.t15 VDD.t14 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X60 VDD.t13 IB.t19 OUT.t22 VDD.t12 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X61 OUT.t17 a_66329_n6784.t24 VSS.t20 VSS.t19 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X62 OUT.t8 a_66329_n6784.t25 VSS.t18 VSS.t17 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X63 OUT.t21 IB.t20 VDD.t11 VDD.t10 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X64 a_66329_n6784.t6 VINP.t9 dw_60815_n7004.t6 dw_60815_n7004.t29 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X65 a_61329_n6784.t2 VINN.t9 dw_60815_n7004.t11 dw_60815_n7004.t10 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X66 VDD.t7 IB.t21 OUT.t20 VDD.t6 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X67 VSS.t16 a_66329_n6784.t26 OUT.t16 VSS.t15 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X68 VSS.t14 a_66329_n6784.t27 OUT.t6 VSS.t13 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X69 VDD.t1 IB.t22 dw_60815_n7004.t28 VDD.t0 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X70 a_55035_n6784.t1 a_55035_n6784.t0 a_55043_n10784 VSS.t3 nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X71 OUT.t1 a_66329_n6784.t28 VSS.t12 VSS.t11 nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
R0 VINN.n0 VINN.t5 49.8994
R1 VINN.n8 VINN.t6 49.6105
R2 VINN.n7 VINN.t4 49.6105
R3 VINN.n6 VINN.t0 49.6105
R4 VINN.n5 VINN.t8 49.6105
R5 VINN.n4 VINN.t1 49.6105
R6 VINN.n3 VINN.t2 49.6105
R7 VINN.n2 VINN.t7 49.6105
R8 VINN.n1 VINN.t3 49.6105
R9 VINN.n0 VINN.t9 49.6105
R10 VINN VINN.n8 19.0298
R11 VINN.n1 VINN.n0 0.289447
R12 VINN.n2 VINN.n1 0.289447
R13 VINN.n3 VINN.n2 0.289447
R14 VINN.n4 VINN.n3 0.289447
R15 VINN.n5 VINN.n4 0.289447
R16 VINN.n6 VINN.n5 0.289447
R17 VINN.n7 VINN.n6 0.289447
R18 VINN.n8 VINN.n7 0.176947
R19 dw_60815_n7004.n1 dw_60815_n7004.t26 201.668
R20 dw_60815_n7004.n0 dw_60815_n7004.t18 201.649
R21 dw_60815_n7004.t18 dw_60815_n7004.t10 148.78
R22 dw_60815_n7004.t10 dw_60815_n7004.t22 148.78
R23 dw_60815_n7004.t22 dw_60815_n7004.t12 148.78
R24 dw_60815_n7004.t12 dw_60815_n7004.t23 148.78
R25 dw_60815_n7004.t23 dw_60815_n7004.t24 148.78
R26 dw_60815_n7004.t24 dw_60815_n7004.t14 148.78
R27 dw_60815_n7004.t14 dw_60815_n7004.t25 148.78
R28 dw_60815_n7004.t25 dw_60815_n7004.t20 148.78
R29 dw_60815_n7004.t20 dw_60815_n7004.t16 148.78
R30 dw_60815_n7004.t26 dw_60815_n7004.t2 148.78
R31 dw_60815_n7004.t2 dw_60815_n7004.t0 148.78
R32 dw_60815_n7004.t0 dw_60815_n7004.t32 148.78
R33 dw_60815_n7004.t32 dw_60815_n7004.t8 148.78
R34 dw_60815_n7004.t8 dw_60815_n7004.t3 148.78
R35 dw_60815_n7004.t3 dw_60815_n7004.t7 148.78
R36 dw_60815_n7004.t7 dw_60815_n7004.t29 148.78
R37 dw_60815_n7004.t29 dw_60815_n7004.t5 148.78
R38 dw_60815_n7004.t5 dw_60815_n7004.t30 148.78
R39 dw_60815_n7004.n0 dw_60815_n7004.t17 4.10017
R40 dw_60815_n7004.n1 dw_60815_n7004.t27 4.10017
R41 dw_60815_n7004.n0 dw_60815_n7004.t31 4.10017
R42 dw_60815_n7004.n0 dw_60815_n7004.t19 4.10017
R43 dw_60815_n7004.n0 dw_60815_n7004.t28 3.91439
R44 dw_60815_n7004.n1 dw_60815_n7004.t9 3.56016
R45 dw_60815_n7004.n0 dw_60815_n7004.t4 3.56016
R46 dw_60815_n7004.n0 dw_60815_n7004.t6 3.56016
R47 dw_60815_n7004.t1 dw_60815_n7004.n1 3.55916
R48 dw_60815_n7004.n0 dw_60815_n7004.t11 3.55898
R49 dw_60815_n7004.n0 dw_60815_n7004.t13 3.55898
R50 dw_60815_n7004.n0 dw_60815_n7004.t15 3.55898
R51 dw_60815_n7004.n0 dw_60815_n7004.t21 3.55898
R52 dw_60815_n7004.n1 dw_60815_n7004.n0 0.992713
R53 a_61329_n6784.n2 a_61329_n6784.t12 46.1695
R54 a_61329_n6784.n2 a_61329_n6784.t0 44.9214
R55 a_61329_n6784.n3 a_61329_n6784.t1 16.544
R56 a_61329_n6784.n1 a_61329_n6784.n7 5.23275
R57 a_61329_n6784.n0 a_61329_n6784.n4 5.19973
R58 a_61329_n6784.n0 a_61329_n6784.n5 5.18121
R59 a_61329_n6784.n1 a_61329_n6784.n6 5.18121
R60 a_61329_n6784.n8 a_61329_n6784.n1 5.18099
R61 a_61329_n6784.n3 a_61329_n6784.n2 0.590649
R62 a_61329_n6784.n0 a_61329_n6784.n3 0.331645
R63 a_61329_n6784.n7 a_61329_n6784.t7 0.2605
R64 a_61329_n6784.n7 a_61329_n6784.t5 0.2605
R65 a_61329_n6784.n6 a_61329_n6784.t9 0.2605
R66 a_61329_n6784.n6 a_61329_n6784.t10 0.2605
R67 a_61329_n6784.n5 a_61329_n6784.t8 0.2605
R68 a_61329_n6784.n5 a_61329_n6784.t4 0.2605
R69 a_61329_n6784.n4 a_61329_n6784.t6 0.2605
R70 a_61329_n6784.n4 a_61329_n6784.t2 0.2605
R71 a_61329_n6784.n8 a_61329_n6784.t3 0.2605
R72 a_61329_n6784.t11 a_61329_n6784.n8 0.2605
R73 a_61329_n6784.n1 a_61329_n6784.n0 0.130746
R74 IB.n21 IB.t5 63.8429
R75 IB.n1 IB.t14 49.8719
R76 IB.n18 IB.t18 49.6432
R77 IB.n0 IB.t4 49.6105
R78 IB.n0 IB.t22 49.6105
R79 IB.n19 IB.t13 49.6105
R80 IB.n17 IB.t3 49.6105
R81 IB.n16 IB.t21 49.6105
R82 IB.n15 IB.t11 49.6105
R83 IB.n14 IB.t9 49.6105
R84 IB.n13 IB.t20 49.6105
R85 IB.n12 IB.t12 49.6105
R86 IB.n11 IB.t2 49.6105
R87 IB.n10 IB.t17 49.6105
R88 IB.n9 IB.t15 49.6105
R89 IB.n8 IB.t10 49.6105
R90 IB.n7 IB.t1 49.6105
R91 IB.n6 IB.t19 49.6105
R92 IB.n5 IB.t6 49.6105
R93 IB.n4 IB.t7 49.6105
R94 IB.n3 IB.t16 49.6105
R95 IB.n2 IB.t8 49.6105
R96 IB.n1 IB.t0 49.6105
R97 IB.n10 IB.n9 16.533
R98 IB.n20 IB.n19 15.2974
R99 IB.n20 IB.n0 13.7519
R100 IB IB.n21 2.039
R101 IB.n21 IB.n20 0.356306
R102 IB.n11 IB.n10 0.285695
R103 IB.n12 IB.n11 0.285695
R104 IB.n13 IB.n12 0.285695
R105 IB.n14 IB.n13 0.285695
R106 IB.n15 IB.n14 0.285695
R107 IB.n16 IB.n15 0.285695
R108 IB.n17 IB.n16 0.285695
R109 IB.n2 IB.n1 0.261929
R110 IB.n3 IB.n2 0.261929
R111 IB.n4 IB.n3 0.261929
R112 IB.n5 IB.n4 0.261929
R113 IB.n6 IB.n5 0.261929
R114 IB.n7 IB.n6 0.261929
R115 IB.n8 IB.n7 0.261929
R116 IB.n9 IB.n8 0.261929
R117 IB.n18 IB.n17 0.236604
R118 IB.n19 IB.n18 0.000848837
R119 VDD.n2 VDD.t0 203.292
R120 VDD.n12 VDD.t4 201.668
R121 VDD.n31 VDD.t8 201.649
R122 VDD.n10 VDD.t34 198.462
R123 VDD.t8 VDD.t40 148.78
R124 VDD.t40 VDD.t22 148.78
R125 VDD.t22 VDD.t10 148.78
R126 VDD.t10 VDD.t26 148.78
R127 VDD.t26 VDD.t2 148.78
R128 VDD.t2 VDD.t6 148.78
R129 VDD.t6 VDD.t38 148.78
R130 VDD.t38 VDD.t20 148.78
R131 VDD.t20 VDD.t14 148.78
R132 VDD.t4 VDD.t44 148.78
R133 VDD.t44 VDD.t28 148.78
R134 VDD.t28 VDD.t16 148.78
R135 VDD.t16 VDD.t30 148.78
R136 VDD.t30 VDD.t32 148.78
R137 VDD.t32 VDD.t12 148.78
R138 VDD.t12 VDD.t42 148.78
R139 VDD.t42 VDD.t24 148.78
R140 VDD.t24 VDD.t18 148.78
R141 VDD.t0 VDD.t36 148.78
R142 VDD.n9 VDD.n0 9.0005
R143 VDD.n9 VDD.n8 9.0005
R144 VDD.n8 VDD.n7 9.0005
R145 VDD.n11 VDD.n10 5.8128
R146 VDD.n3 VDD.t37 5.72121
R147 VDD.n2 VDD.t1 5.72002
R148 VDD.n6 VDD.n1 4.50853
R149 VDD.n5 VDD.n4 4.49348
R150 VDD.n7 VDD.n6 4.49348
R151 VDD.n23 VDD.t15 4.17154
R152 VDD.n12 VDD.t5 4.10017
R153 VDD.n21 VDD.t19 4.10017
R154 VDD.n30 VDD.t9 4.10017
R155 VDD.n33 VDD.n32 3.87873
R156 VDD.n14 VDD.n13 3.56016
R157 VDD.n16 VDD.n15 3.56016
R158 VDD.n18 VDD.n17 3.56016
R159 VDD.n20 VDD.n19 3.56016
R160 VDD.n29 VDD.n28 3.56016
R161 VDD.n27 VDD.n26 3.56016
R162 VDD.n25 VDD.n24 3.56016
R163 VDD.n23 VDD.n22 3.56016
R164 VDD.n10 VDD.t35 0.911929
R165 VDD VDD.n33 0.878874
R166 VDD.n33 VDD.n11 0.532701
R167 VDD.n11 VDD.n9 0.494214
R168 VDD.n22 VDD.t39 0.2605
R169 VDD.n22 VDD.t21 0.2605
R170 VDD.n24 VDD.t3 0.2605
R171 VDD.n24 VDD.t7 0.2605
R172 VDD.n26 VDD.t11 0.2605
R173 VDD.n26 VDD.t27 0.2605
R174 VDD.n28 VDD.t41 0.2605
R175 VDD.n28 VDD.t23 0.2605
R176 VDD.n19 VDD.t43 0.2605
R177 VDD.n19 VDD.t25 0.2605
R178 VDD.n17 VDD.t33 0.2605
R179 VDD.n17 VDD.t13 0.2605
R180 VDD.n15 VDD.t17 0.2605
R181 VDD.n15 VDD.t31 0.2605
R182 VDD.n13 VDD.t45 0.2605
R183 VDD.n13 VDD.t29 0.2605
R184 VDD.n8 VDD.n3 0.162259
R185 VDD.n32 VDD.n31 0.153411
R186 VDD.n32 VDD.n21 0.150525
R187 VDD.n3 VDD.n2 0.091103
R188 VDD.n21 VDD.n20 0.0720015
R189 VDD.n30 VDD.n29 0.0718703
R190 VDD.n14 VDD.n12 0.0717391
R191 VDD.n16 VDD.n14 0.0645233
R192 VDD.n18 VDD.n16 0.0645233
R193 VDD.n20 VDD.n18 0.0645233
R194 VDD.n29 VDD.n27 0.0645233
R195 VDD.n27 VDD.n25 0.0645233
R196 VDD.n25 VDD.n23 0.0645233
R197 VDD.n7 VDD.n5 0.0326429
R198 VDD.n31 VDD.n30 0.0196545
R199 VDD.n9 VDD.n1 0.0170428
R200 VDD.n5 VDD.n1 0.0170428
R201 VDD.n4 VDD.n0 0.0160502
R202 VDD.n8 VDD.n4 0.0160502
R203 VDD.n6 VDD.n0 0.0160502
R204 OUT.n2 OUT.n0 14.8246
R205 OUT.n2 OUT.n1 14.6677
R206 OUT.n4 OUT.n3 14.6677
R207 OUT.n6 OUT.n5 14.6677
R208 OUT.n8 OUT.n7 14.6677
R209 OUT.n10 OUT.n9 14.6677
R210 OUT.n12 OUT.n11 14.6677
R211 OUT.n14 OUT.n13 14.6677
R212 OUT.n16 OUT.n15 14.6677
R213 OUT.n18 OUT.n17 14.6677
R214 OUT OUT.n39 8.1668
R215 OUT.n21 OUT.n19 5.25392
R216 OUT.n28 OUT.n26 5.25392
R217 OUT.n21 OUT.n20 5.18121
R218 OUT.n23 OUT.n22 5.18121
R219 OUT.n25 OUT.n24 5.18121
R220 OUT.n36 OUT.n35 5.18121
R221 OUT.n34 OUT.n33 5.18121
R222 OUT.n32 OUT.n31 5.18121
R223 OUT.n30 OUT.n29 5.18121
R224 OUT.n28 OUT.n27 5.18121
R225 OUT.n39 OUT.t40 4.9497
R226 OUT.n39 OUT.n38 1.38146
R227 OUT.n38 OUT.n37 1.12455
R228 OUT.n0 OUT.t12 0.4685
R229 OUT.n0 OUT.t18 0.4685
R230 OUT.n1 OUT.t16 0.4685
R231 OUT.n1 OUT.t14 0.4685
R232 OUT.n3 OUT.t11 0.4685
R233 OUT.n3 OUT.t1 0.4685
R234 OUT.n5 OUT.t15 0.4685
R235 OUT.n5 OUT.t5 0.4685
R236 OUT.n7 OUT.t6 0.4685
R237 OUT.n7 OUT.t13 0.4685
R238 OUT.n9 OUT.t9 0.4685
R239 OUT.n9 OUT.t2 0.4685
R240 OUT.n11 OUT.t10 0.4685
R241 OUT.n11 OUT.t7 0.4685
R242 OUT.n13 OUT.t3 0.4685
R243 OUT.n13 OUT.t17 0.4685
R244 OUT.n15 OUT.t4 0.4685
R245 OUT.n15 OUT.t8 0.4685
R246 OUT.n17 OUT.t0 0.4685
R247 OUT.n17 OUT.t19 0.4685
R248 OUT.n36 OUT.n34 0.454672
R249 OUT.n26 OUT.t28 0.2605
R250 OUT.n26 OUT.t23 0.2605
R251 OUT.n27 OUT.t20 0.2605
R252 OUT.n27 OUT.t36 0.2605
R253 OUT.n29 OUT.t32 0.2605
R254 OUT.n29 OUT.t30 0.2605
R255 OUT.n31 OUT.t29 0.2605
R256 OUT.n31 OUT.t21 0.2605
R257 OUT.n33 OUT.t24 0.2605
R258 OUT.n33 OUT.t37 0.2605
R259 OUT.n35 OUT.t31 0.2605
R260 OUT.n35 OUT.t26 0.2605
R261 OUT.n24 OUT.t22 0.2605
R262 OUT.n24 OUT.t38 0.2605
R263 OUT.n22 OUT.t34 0.2605
R264 OUT.n22 OUT.t35 0.2605
R265 OUT.n20 OUT.t33 0.2605
R266 OUT.n20 OUT.t25 0.2605
R267 OUT.n19 OUT.t27 0.2605
R268 OUT.n19 OUT.t39 0.2605
R269 OUT.n38 OUT.n18 0.220357
R270 OUT.n18 OUT.n16 0.157357
R271 OUT.n16 OUT.n14 0.157357
R272 OUT.n14 OUT.n12 0.157357
R273 OUT.n12 OUT.n10 0.157357
R274 OUT.n10 OUT.n8 0.157357
R275 OUT.n8 OUT.n6 0.157357
R276 OUT.n6 OUT.n4 0.157357
R277 OUT.n4 OUT.n2 0.157357
R278 OUT.n23 OUT.n21 0.0732152
R279 OUT.n25 OUT.n23 0.0732152
R280 OUT.n34 OUT.n32 0.0732152
R281 OUT.n32 OUT.n30 0.0732152
R282 OUT.n30 OUT.n28 0.0732152
R283 OUT.n37 OUT.n25 0.0407318
R284 OUT.n37 OUT.n36 0.0329834
R285 a_66329_n6784.n5 a_66329_n6784.t23 31.5452
R286 a_66329_n6784.n6 a_66329_n6784.t22 31.2562
R287 a_66329_n6784.n6 a_66329_n6784.t19 31.2562
R288 a_66329_n6784.n6 a_66329_n6784.t10 31.2562
R289 a_66329_n6784.n6 a_66329_n6784.t26 31.2562
R290 a_66329_n6784.n3 a_66329_n6784.t28 31.2562
R291 a_66329_n6784.n3 a_66329_n6784.t20 31.2562
R292 a_66329_n6784.n3 a_66329_n6784.t17 31.2562
R293 a_66329_n6784.n3 a_66329_n6784.t9 31.2562
R294 a_66329_n6784.n2 a_66329_n6784.t14 31.2562
R295 a_66329_n6784.n2 a_66329_n6784.t27 31.2562
R296 a_66329_n6784.n2 a_66329_n6784.t21 31.2562
R297 a_66329_n6784.n2 a_66329_n6784.t16 31.2562
R298 a_66329_n6784.n4 a_66329_n6784.t15 31.2562
R299 a_66329_n6784.n4 a_66329_n6784.t12 31.2562
R300 a_66329_n6784.n4 a_66329_n6784.t24 31.2562
R301 a_66329_n6784.n4 a_66329_n6784.t18 31.2562
R302 a_66329_n6784.n5 a_66329_n6784.t25 31.2562
R303 a_66329_n6784.n5 a_66329_n6784.t13 31.2562
R304 a_66329_n6784.n5 a_66329_n6784.t11 31.2562
R305 a_66329_n6784.n1 a_66329_n6784.n8 16.5173
R306 a_66329_n6784.n0 a_66329_n6784.t8 16.349
R307 a_66329_n6784.n0 a_66329_n6784.n6 15.9887
R308 a_66329_n6784.n7 a_66329_n6784.t7 11.403
R309 a_66329_n6784.n7 a_66329_n6784.t0 10.2897
R310 a_66329_n6784.n8 a_66329_n6784.n7 9.4158
R311 a_66329_n6784.n1 a_66329_n6784.t2 5.25416
R312 a_66329_n6784.n1 a_66329_n6784.t5 5.25416
R313 a_66329_n6784.n1 a_66329_n6784.t3 5.18121
R314 a_66329_n6784.n1 a_66329_n6784.t6 5.18121
R315 a_66329_n6784.t1 a_66329_n6784.n1 5.18099
R316 a_66329_n6784.n8 a_66329_n6784.t4 1.9865
R317 a_66329_n6784.n6 a_66329_n6784.n3 1.65129
R318 a_66329_n6784.n1 a_66329_n6784.n0 1.59414
R319 a_66329_n6784.n4 a_66329_n6784.n5 1.15629
R320 a_66329_n6784.n2 a_66329_n6784.n4 1.15629
R321 a_66329_n6784.n3 a_66329_n6784.n2 1.15629
R322 VSS.n152 VSS.n13 1386.58
R323 VSS.n155 VSS.n152 1386.58
R324 VSS.n146 VSS.n25 1352.79
R325 VSS.n146 VSS.n26 1352.79
R326 VSS.n140 VSS.n31 1352.79
R327 VSS.n140 VSS.n32 1352.79
R328 VSS.n134 VSS.n37 1352.79
R329 VSS.n134 VSS.n133 1352.79
R330 VSS.n165 VSS.n164 1230.38
R331 VSS.n164 VSS.n163 1230.38
R332 VSS.n176 VSS.n175 823.048
R333 VSS.n118 VSS.t7 650.366
R334 VSS.t23 VSS.n32 608.688
R335 VSS.n124 VSS.n112 570.674
R336 VSS.n57 VSS.n46 570.674
R337 VSS.n183 VSS.n1 570.674
R338 VSS.n95 VSS.n86 558.308
R339 VSS.n97 VSS.n66 525.789
R340 VSS.n131 VSS.n126 496.264
R341 VSS.n126 VSS.n39 496.264
R342 VSS.n41 VSS.n39 496.264
R343 VSS.n131 VSS.n41 496.264
R344 VSS.n125 VSS.n124 466.25
R345 VSS.n156 VSS.n12 466.25
R346 VSS.n163 VSS.n162 461.212
R347 VSS.n118 VSS.n26 416.327
R348 VSS.n156 VSS.n155 397.091
R349 VSS.t5 VSS.n48 379.687
R350 VSS.t3 VSS.n8 368.695
R351 VSS.n89 VSS.n37 349.252
R352 VSS.n37 VSS.n36 349.252
R353 VSS.n36 VSS.n31 349.252
R354 VSS.n31 VSS.n30 349.252
R355 VSS.n30 VSS.n25 349.252
R356 VSS.n25 VSS.n24 349.252
R357 VSS.n24 VSS.n13 345.899
R358 VSS.n147 VSS.n21 336.462
R359 VSS.n151 VSS.n21 336.462
R360 VSS.n147 VSS.n22 336.462
R361 VSS.n151 VSS.n22 336.462
R362 VSS.n141 VSS.n27 336.462
R363 VSS.n145 VSS.n27 336.462
R364 VSS.n141 VSS.n28 336.462
R365 VSS.n145 VSS.n28 336.462
R366 VSS.n135 VSS.n33 336.462
R367 VSS.n139 VSS.n33 336.462
R368 VSS.n135 VSS.n34 336.462
R369 VSS.n139 VSS.n34 336.462
R370 VSS.n90 VSS.n87 336.462
R371 VSS.n90 VSS.n38 336.462
R372 VSS.n94 VSS.n38 336.462
R373 VSS.n94 VSS.n87 336.462
R374 VSS.n103 VSS.n98 316.474
R375 VSS.n98 VSS.n64 316.474
R376 VSS.n64 VSS.n63 316.474
R377 VSS.n103 VSS.n63 316.474
R378 VSS.n161 VSS.n9 282.764
R379 VSS.n161 VSS.n10 282.764
R380 VSS.n157 VSS.n10 282.764
R381 VSS.n157 VSS.n9 282.764
R382 VSS.n55 VSS.n50 282.764
R383 VSS.n50 VSS.n47 282.764
R384 VSS.n49 VSS.n47 282.764
R385 VSS.n55 VSS.n49 282.764
R386 VSS.n119 VSS.n113 282.764
R387 VSS.n119 VSS.n114 282.764
R388 VSS.n123 VSS.n114 282.764
R389 VSS.n123 VSS.n113 282.764
R390 VSS.n169 VSS.n166 282.764
R391 VSS.n173 VSS.n166 282.764
R392 VSS.n169 VSS.n167 282.764
R393 VSS.n173 VSS.n167 282.764
R394 VSS.n162 VSS.n8 281.673
R395 VSS.n48 VSS.n12 270.682
R396 VSS.n175 VSS.n174 264.901
R397 VSS.n20 VSS.n14 246.566
R398 VSS.n14 VSS.n7 246.566
R399 VSS.n15 VSS.n7 246.566
R400 VSS.n20 VSS.n15 246.566
R401 VSS.n177 VSS.n3 235.329
R402 VSS.n177 VSS.n4 235.329
R403 VSS.n181 VSS.n3 235.329
R404 VSS.n181 VSS.n4 235.329
R405 VSS.n165 VSS.n6 226.595
R406 VSS.n89 VSS.n66 211.648
R407 VSS.n13 VSS.n6 209.552
R408 VSS.n176 VSS.n165 209.552
R409 VSS.n155 VSS.n154 173.584
R410 VSS.n174 VSS.t9 160.933
R411 VSS.n97 VSS.n96 155.722
R412 VSS.n86 VSS.t21 144.73
R413 VSS.n105 VSS.n63 126.71
R414 VSS.n57 VSS.n56 112.212
R415 VSS.n154 VSS.n153 112.212
R416 VSS.t21 VSS.t45 111.754
R417 VSS.t45 VSS.t41 111.754
R418 VSS.t41 VSS.t17 111.754
R419 VSS.t31 VSS.t19 111.754
R420 VSS.t19 VSS.t43 111.754
R421 VSS.t43 VSS.t37 111.754
R422 VSS.t37 VSS.t35 111.754
R423 VSS.t35 VSS.t25 111.754
R424 VSS.t13 VSS.t39 111.754
R425 VSS.t39 VSS.t49 111.754
R426 VSS.t49 VSS.t33 111.754
R427 VSS.t33 VSS.t27 111.754
R428 VSS.t11 VSS.t15 111.754
R429 VSS.t15 VSS.t47 111.754
R430 VSS.t47 VSS.t29 111.754
R431 VSS.t29 VSS.t23 111.754
R432 VSS.n183 VSS.n182 111.296
R433 VSS.n133 VSS.t17 106.716
R434 VSS.n40 VSS.t11 89.3114
R435 VSS.n132 VSS.t13 88.3954
R436 VSS.n116 VSS.n112 66.4112
R437 VSS.n46 VSS.n26 49.923
R438 VSS.n117 VSS.n116 45.8009
R439 VSS.n125 VSS.n32 41.6789
R440 VSS.t7 VSS.n117 32.5188
R441 VSS.n56 VSS.t5 32.5188
R442 VSS.n153 VSS.t3 32.5188
R443 VSS.t9 VSS.n2 32.5188
R444 VSS.n105 VSS.t4 32.0943
R445 VSS.n66 VSS.t2 27.6255
R446 VSS.t4 VSS.t1 24.7817
R447 VSS.t2 VSS.t0 24.7817
R448 VSS.t25 VSS.n132 23.3587
R449 VSS.t27 VSS.n40 22.4427
R450 VSS.t0 VSS.n65 16.4536
R451 VSS.n185 VSS.n184 14.7588
R452 VSS.n110 VSS.n109 13.5005
R453 VSS.n110 VSS.n42 13.5005
R454 VSS.n60 VSS.n42 13.5005
R455 VSS.n106 VSS.n105 13.0989
R456 VSS.n96 VSS.n95 12.3666
R457 VSS.n154 VSS.n0 12.111
R458 VSS.n62 VSS.t24 11.2257
R459 VSS.n85 VSS.t22 11.2245
R460 VSS.n86 VSS.n85 11.0164
R461 VSS.n68 VSS.n67 10.2897
R462 VSS.n70 VSS.n69 10.2897
R463 VSS.n72 VSS.n71 10.2897
R464 VSS.n74 VSS.n73 10.2897
R465 VSS.n76 VSS.n75 10.2897
R466 VSS.n78 VSS.n77 10.2897
R467 VSS.n80 VSS.n79 10.2897
R468 VSS.n82 VSS.n81 10.2897
R469 VSS.n84 VSS.n83 10.2897
R470 VSS VSS.n185 10.2753
R471 VSS.n106 VSS 8.95964
R472 VSS.n59 VSS.n58 6.98379
R473 VSS.n111 VSS.n110 6.96369
R474 VSS.n59 VSS.n45 6.74471
R475 VSS.n109 VSS.n61 6.74333
R476 VSS.n44 VSS.n43 6.74333
R477 VSS.n130 VSS.n129 6.38103
R478 VSS.n129 VSS.n128 6.38103
R479 VSS.n128 VSS.n127 6.38103
R480 VSS.n130 VSS.n127 6.38103
R481 VSS.n107 VSS.n62 5.45103
R482 VSS.t1 VSS.n104 5.18019
R483 VSS.n133 VSS.t31 5.03855
R484 VSS.n163 VSS.n1 5.03855
R485 VSS.n148 VSS.n23 4.32642
R486 VSS.n150 VSS.n23 4.32642
R487 VSS.n150 VSS.n149 4.32642
R488 VSS.n149 VSS.n148 4.32642
R489 VSS.n142 VSS.n29 4.32642
R490 VSS.n144 VSS.n29 4.32642
R491 VSS.n144 VSS.n143 4.32642
R492 VSS.n143 VSS.n142 4.32642
R493 VSS.n136 VSS.n35 4.32642
R494 VSS.n138 VSS.n35 4.32642
R495 VSS.n138 VSS.n137 4.32642
R496 VSS.n137 VSS.n136 4.32642
R497 VSS.n91 VSS.n88 4.32642
R498 VSS.n92 VSS.n91 4.32642
R499 VSS.n93 VSS.n88 4.32642
R500 VSS.n93 VSS.n92 4.32642
R501 VSS.n102 VSS.n101 4.06945
R502 VSS.n101 VSS.n100 4.06945
R503 VSS.n100 VSS.n99 4.06945
R504 VSS.n102 VSS.n99 4.06945
R505 VSS.n160 VSS.n11 3.63603
R506 VSS.n160 VSS.n159 3.63603
R507 VSS.n159 VSS.n158 3.63603
R508 VSS.n158 VSS.n11 3.63603
R509 VSS.n54 VSS.n53 3.63603
R510 VSS.n53 VSS.n52 3.63603
R511 VSS.n52 VSS.n51 3.63603
R512 VSS.n54 VSS.n51 3.63603
R513 VSS.n120 VSS.n115 3.63603
R514 VSS.n121 VSS.n120 3.63603
R515 VSS.n122 VSS.n121 3.63603
R516 VSS.n122 VSS.n115 3.63603
R517 VSS.n170 VSS.n168 3.63603
R518 VSS.n172 VSS.n168 3.63603
R519 VSS.n171 VSS.n170 3.63603
R520 VSS.n172 VSS.n171 3.63603
R521 VSS.n112 VSS.n111 3.21476
R522 VSS.n19 VSS.n16 3.17063
R523 VSS.n17 VSS.n16 3.17063
R524 VSS.n18 VSS.n17 3.17063
R525 VSS.n19 VSS.n18 3.17063
R526 VSS.n104 VSS.n65 3.14894
R527 VSS.n178 VSS.n5 3.02616
R528 VSS.n179 VSS.n178 3.02616
R529 VSS.n180 VSS.n5 3.02616
R530 VSS.n180 VSS.n179 3.02616
R531 VSS.n58 VSS.t6 2.00831
R532 VSS.n111 VSS.t8 2.00069
R533 VSS.n184 VSS.t10 1.9865
R534 VSS.n58 VSS.n57 1.73383
R535 VSS.n184 VSS.n183 1.73383
R536 VSS.n107 VSS.n106 1.36388
R537 VSS.n182 VSS.n2 0.916509
R538 VSS.n108 VSS.n0 0.700336
R539 VSS.n185 VSS.n0 0.510623
R540 VSS.n108 VSS.n107 0.493902
R541 VSS.n67 VSS.t48 0.4685
R542 VSS.n67 VSS.t30 0.4685
R543 VSS.n69 VSS.t12 0.4685
R544 VSS.n69 VSS.t16 0.4685
R545 VSS.n71 VSS.t34 0.4685
R546 VSS.n71 VSS.t28 0.4685
R547 VSS.n73 VSS.t40 0.4685
R548 VSS.n73 VSS.t50 0.4685
R549 VSS.n75 VSS.t26 0.4685
R550 VSS.n75 VSS.t14 0.4685
R551 VSS.n77 VSS.t38 0.4685
R552 VSS.n77 VSS.t36 0.4685
R553 VSS.n79 VSS.t20 0.4685
R554 VSS.n79 VSS.t44 0.4685
R555 VSS.n81 VSS.t18 0.4685
R556 VSS.n81 VSS.t32 0.4685
R557 VSS.n83 VSS.t46 0.4685
R558 VSS.n83 VSS.t42 0.4685
R559 VSS.n109 VSS.n108 0.333185
R560 VSS.n178 VSS.n177 0.2605
R561 VSS.n177 VSS.n176 0.2605
R562 VSS.n181 VSS.n180 0.2605
R563 VSS.n182 VSS.n181 0.2605
R564 VSS.n16 VSS.n14 0.226587
R565 VSS.n14 VSS.n6 0.226587
R566 VSS.n18 VSS.n15 0.226587
R567 VSS.n15 VSS.n8 0.226587
R568 VSS.n179 VSS.n4 0.17981
R569 VSS.n175 VSS.n4 0.17981
R570 VSS.n20 VSS.n19 0.17981
R571 VSS.n152 VSS.n20 0.17981
R572 VSS.n151 VSS.n150 0.17981
R573 VSS.n152 VSS.n151 0.17981
R574 VSS.n148 VSS.n147 0.17981
R575 VSS.n147 VSS.n146 0.17981
R576 VSS.n145 VSS.n144 0.17981
R577 VSS.n146 VSS.n145 0.17981
R578 VSS.n142 VSS.n141 0.17981
R579 VSS.n141 VSS.n140 0.17981
R580 VSS.n139 VSS.n138 0.17981
R581 VSS.n140 VSS.n139 0.17981
R582 VSS.n88 VSS.n87 0.17981
R583 VSS.n87 VSS.n65 0.17981
R584 VSS.n92 VSS.n38 0.17981
R585 VSS.n134 VSS.n38 0.17981
R586 VSS.n136 VSS.n135 0.17981
R587 VSS.n135 VSS.n134 0.17981
R588 VSS.n17 VSS.n7 0.17981
R589 VSS.n164 VSS.n7 0.17981
R590 VSS.n5 VSS.n3 0.17981
R591 VSS.n164 VSS.n3 0.17981
R592 VSS.n115 VSS.n113 0.17981
R593 VSS.n117 VSS.n113 0.17981
R594 VSS.n121 VSS.n114 0.17981
R595 VSS.n117 VSS.n114 0.17981
R596 VSS.n55 VSS.n54 0.17981
R597 VSS.n56 VSS.n55 0.17981
R598 VSS.n52 VSS.n47 0.17981
R599 VSS.n56 VSS.n47 0.17981
R600 VSS.n11 VSS.n9 0.17981
R601 VSS.n153 VSS.n9 0.17981
R602 VSS.n159 VSS.n10 0.17981
R603 VSS.n153 VSS.n10 0.17981
R604 VSS.n168 VSS.n166 0.17981
R605 VSS.n166 VSS.n2 0.17981
R606 VSS.n171 VSS.n167 0.17981
R607 VSS.n167 VSS.n2 0.17981
R608 VSS.n85 VSS.n84 0.16925
R609 VSS.n68 VSS.n62 0.16925
R610 VSS.n173 VSS.n172 0.163
R611 VSS.n174 VSS.n173 0.163
R612 VSS.n99 VSS.n63 0.163
R613 VSS.n101 VSS.n98 0.163
R614 VSS.n98 VSS.n97 0.163
R615 VSS.n127 VSS.n41 0.163
R616 VSS.n96 VSS.n41 0.163
R617 VSS.n129 VSS.n126 0.163
R618 VSS.n126 VSS.n125 0.163
R619 VSS.n123 VSS.n122 0.163
R620 VSS.n124 VSS.n123 0.163
R621 VSS.n120 VSS.n119 0.163
R622 VSS.n119 VSS.n118 0.163
R623 VSS.n51 VSS.n49 0.163
R624 VSS.n49 VSS.n46 0.163
R625 VSS.n53 VSS.n50 0.163
R626 VSS.n50 VSS.n12 0.163
R627 VSS.n158 VSS.n157 0.163
R628 VSS.n157 VSS.n156 0.163
R629 VSS.n161 VSS.n160 0.163
R630 VSS.n162 VSS.n161 0.163
R631 VSS.n170 VSS.n169 0.163
R632 VSS.n169 VSS.n1 0.163
R633 VSS.n84 VSS.n82 0.153
R634 VSS.n82 VSS.n80 0.153
R635 VSS.n80 VSS.n78 0.153
R636 VSS.n78 VSS.n76 0.153
R637 VSS.n76 VSS.n74 0.153
R638 VSS.n74 VSS.n72 0.153
R639 VSS.n72 VSS.n70 0.153
R640 VSS.n70 VSS.n68 0.153
R641 VSS.n103 VSS.n102 0.144944
R642 VSS.n104 VSS.n103 0.144944
R643 VSS.n100 VSS.n64 0.144944
R644 VSS.n104 VSS.n64 0.144944
R645 VSS.n91 VSS.n90 0.118682
R646 VSS.n90 VSS.n89 0.118682
R647 VSS.n35 VSS.n33 0.118682
R648 VSS.n36 VSS.n33 0.118682
R649 VSS.n29 VSS.n27 0.118682
R650 VSS.n30 VSS.n27 0.118682
R651 VSS.n23 VSS.n21 0.118682
R652 VSS.n24 VSS.n21 0.118682
R653 VSS.n94 VSS.n93 0.118682
R654 VSS.n95 VSS.n94 0.118682
R655 VSS.n137 VSS.n34 0.118682
R656 VSS.n40 VSS.n34 0.118682
R657 VSS.n143 VSS.n28 0.118682
R658 VSS.n116 VSS.n28 0.118682
R659 VSS.n149 VSS.n22 0.118682
R660 VSS.n48 VSS.n22 0.118682
R661 VSS.n131 VSS.n130 0.0663228
R662 VSS.n132 VSS.n131 0.0663228
R663 VSS.n128 VSS.n39 0.0663228
R664 VSS.n132 VSS.n39 0.0663228
R665 VSS.n109 VSS.n44 0.0256748
R666 VSS.n60 VSS.n43 0.0163409
R667 VSS.n61 VSS.n60 0.0163409
R668 VSS.n61 VSS.n59 0.0163409
R669 VSS.n110 VSS.n43 0.0163409
R670 VSS.n45 VSS.n44 0.0135757
R671 VSS.n45 VSS.n42 0.0135757
R672 a_55035_n6784.n0 a_55035_n6784.t5 31.5452
R673 a_55035_n6784.n0 a_55035_n6784.t4 31.5433
R674 a_55035_n6784.n1 a_55035_n6784.t0 31.4426
R675 a_55035_n6784.n0 a_55035_n6784.t3 31.2562
R676 a_55035_n6784.n0 a_55035_n6784.t6 31.2562
R677 a_55035_n6784.n2 a_55035_n6784.n0 18.5063
R678 a_55035_n6784.t2 a_55035_n6784.n2 14.5399
R679 a_55035_n6784.n2 a_55035_n6784.n1 10.5733
R680 a_55035_n6784.n1 a_55035_n6784.t1 2.46966
R681 a_79287_n10784.t2 a_79287_n10784.t0 14.6706
R682 a_79287_n10784.t1 a_79287_n10784.t2 14.6695
R683 VINP.n0 VINP.t5 49.8994
R684 VINP.n8 VINP.t4 49.6105
R685 VINP.n0 VINP.t3 49.6105
R686 VINP.n1 VINP.t9 49.6105
R687 VINP.n2 VINP.t7 49.6105
R688 VINP.n3 VINP.t1 49.6105
R689 VINP.n4 VINP.t0 49.6105
R690 VINP.n5 VINP.t6 49.6105
R691 VINP.n6 VINP.t2 49.6105
R692 VINP.n7 VINP.t8 49.6105
R693 VINP VINP.n8 21.7674
R694 VINP.n7 VINP.n6 0.289447
R695 VINP.n6 VINP.n5 0.289447
R696 VINP.n5 VINP.n4 0.289447
R697 VINP.n4 VINP.n3 0.289447
R698 VINP.n3 VINP.n2 0.289447
R699 VINP.n2 VINP.n1 0.289447
R700 VINP.n1 VINP.n0 0.289447
R701 VINP.n8 VINP.n7 0.226684
C0 VINN VDD 0.696662f
C1 IB w_54815_n7004 0.044345f
C2 w_70815_n7004 IB 0.387961f
C3 IB w_75815_n7004 0.387961f
C4 w_57815_n7004 IB 0.082524f
C5 VINN w_60815_n7004 0.387961f
C6 OUT IB 3.7759f
C7 IB VDD 11.506201f
C8 VINP w_65815_n7004 0.387961f
C9 OUT VDD 11.5628f
C10 VINP IB 0.822556f
C11 VSS OUT 8.207049f
C12 VINN IB 0.53823f
C13 VINP VDD 3.40615f
C14 VSS a_55043_n10784 0.443171f
C15 OUT a_53801_n12052 97.8273f
C16 VINP a_53801_n12052 62.24887f
C17 VINN a_53801_n12052 56.24142f
C18 IB a_53801_n12052 0.109142p
C19 VSS a_53801_n12052 0.269017p
C20 VDD a_53801_n12052 0.142194p
C21 a_55043_n10784 a_53801_n12052 1.97668f
C22 VINP.n8 a_53801_n12052 0.040687f
C23 a_79287_n10784.t0 a_53801_n12052 0.077925f
C24 a_79287_n10784.t1 a_53801_n12052 0.077819f
C25 a_79287_n10784.t2 a_53801_n12052 3.04426f
C26 a_55035_n6784.n0 a_53801_n12052 0.626928f
C27 a_55035_n6784.t1 a_53801_n12052 0.039343f
C28 a_55035_n6784.t0 a_53801_n12052 0.037798f
C29 a_55035_n6784.n1 a_53801_n12052 0.071066f
C30 a_55035_n6784.t5 a_53801_n12052 0.037861f
C31 a_55035_n6784.t6 a_53801_n12052 0.037695f
C32 a_55035_n6784.t4 a_53801_n12052 0.03786f
C33 a_55035_n6784.t3 a_53801_n12052 0.037695f
C34 a_55035_n6784.n2 a_53801_n12052 1.88231f
C35 a_55035_n6784.t2 a_53801_n12052 0.191442f
C36 VSS.n0 a_53801_n12052 0.012175f
C37 VSS.n1 a_53801_n12052 0.013626f
C38 VSS.n6 a_53801_n12052 0.110951f
C39 VSS.n8 a_53801_n12052 0.015393f
C40 VSS.n12 a_53801_n12052 0.017441f
C41 VSS.n13 a_53801_n12052 0.143708f
C42 VSS.n24 a_53801_n12052 0.176839f
C43 VSS.n25 a_53801_n12052 0.18016f
C44 VSS.n26 a_53801_n12052 0.013503f
C45 VSS.n30 a_53801_n12052 0.177692f
C46 VSS.n31 a_53801_n12052 0.18016f
C47 VSS.n32 a_53801_n12052 0.01786f
C48 VSS.n36 a_53801_n12052 0.177692f
C49 VSS.n37 a_53801_n12052 0.18016f
C50 VSS.t23 a_53801_n12052 0.017051f
C51 VSS.n46 a_53801_n12052 0.014688f
C52 VSS.n48 a_53801_n12052 0.015393f
C53 VSS.n57 a_53801_n12052 0.01601f
C54 VSS.n63 a_53801_n12052 5.57733f
C55 VSS.t0 a_53801_n12052 0.019847f
C56 VSS.t2 a_53801_n12052 0.025224f
C57 VSS.n66 a_53801_n12052 0.079581f
C58 VSS.n86 a_53801_n12052 0.016466f
C59 VSS.n89 a_53801_n12052 0.142687f
C60 VSS.n95 a_53801_n12052 0.013507f
C61 VSS.n97 a_53801_n12052 0.01613f
C62 VSS.t1 a_53801_n12052 0.014421f
C63 VSS.t4 a_53801_n12052 0.027375f
C64 VSS.n105 a_53801_n12052 0.083907f
C65 VSS.n106 a_53801_n12052 0.104518f
C66 VSS.n107 a_53801_n12052 0.021379f
C67 VSS.n108 a_53801_n12052 0.013739f
C68 VSS.n112 a_53801_n12052 0.014957f
C69 VSS.t7 a_53801_n12052 0.016162f
C70 VSS.n118 a_53801_n12052 0.025246f
C71 VSS.n124 a_53801_n12052 0.024542f
C72 VSS.n125 a_53801_n12052 0.012021f
C73 VSS.n155 a_53801_n12052 0.015914f
C74 VSS.n156 a_53801_n12052 0.020433f
C75 VSS.n162 a_53801_n12052 0.017582f
C76 VSS.n163 a_53801_n12052 0.013748f
C77 VSS.n165 a_53801_n12052 0.113664f
C78 VSS.t9 a_53801_n12052 0.01671f
C79 VSS.n174 a_53801_n12052 0.922641f
C80 VSS.n175 a_53801_n12052 1.56057f
C81 VSS.n176 a_53801_n12052 2.76461f
C82 VSS.n183 a_53801_n12052 0.015989f
C83 VSS.n185 a_53801_n12052 0.105635f
C84 a_66329_n6784.n0 a_53801_n12052 1.15805f
C85 a_66329_n6784.n1 a_53801_n12052 7.42529f
C86 a_66329_n6784.n2 a_53801_n12052 0.292895f
C87 a_66329_n6784.n3 a_53801_n12052 0.292895f
C88 a_66329_n6784.n4 a_53801_n12052 0.292895f
C89 a_66329_n6784.n5 a_53801_n12052 0.282049f
C90 a_66329_n6784.n6 a_53801_n12052 0.420764f
C91 a_66329_n6784.t0 a_53801_n12052 0.175353f
C92 a_66329_n6784.t5 a_53801_n12052 0.403984f
C93 a_66329_n6784.t6 a_53801_n12052 0.395506f
C94 a_66329_n6784.t3 a_53801_n12052 0.395506f
C95 a_66329_n6784.t2 a_53801_n12052 0.404038f
C96 a_66329_n6784.t1 a_53801_n12052 0.395497f
C97 a_66329_n6784.t23 a_53801_n12052 0.131027f
C98 a_66329_n6784.t11 a_53801_n12052 0.13045f
C99 a_66329_n6784.t13 a_53801_n12052 0.13045f
C100 a_66329_n6784.t25 a_53801_n12052 0.13045f
C101 a_66329_n6784.t18 a_53801_n12052 0.13045f
C102 a_66329_n6784.t24 a_53801_n12052 0.13045f
C103 a_66329_n6784.t12 a_53801_n12052 0.13045f
C104 a_66329_n6784.t15 a_53801_n12052 0.13045f
C105 a_66329_n6784.t16 a_53801_n12052 0.13045f
C106 a_66329_n6784.t21 a_53801_n12052 0.13045f
C107 a_66329_n6784.t27 a_53801_n12052 0.13045f
C108 a_66329_n6784.t14 a_53801_n12052 0.13045f
C109 a_66329_n6784.t9 a_53801_n12052 0.13045f
C110 a_66329_n6784.t17 a_53801_n12052 0.13045f
C111 a_66329_n6784.t20 a_53801_n12052 0.13045f
C112 a_66329_n6784.t28 a_53801_n12052 0.13045f
C113 a_66329_n6784.t26 a_53801_n12052 0.13045f
C114 a_66329_n6784.t10 a_53801_n12052 0.13045f
C115 a_66329_n6784.t19 a_53801_n12052 0.13045f
C116 a_66329_n6784.t22 a_53801_n12052 0.13045f
C117 a_66329_n6784.t8 a_53801_n12052 0.235332f
C118 a_66329_n6784.t7 a_53801_n12052 0.211657f
C119 a_66329_n6784.n7 a_53801_n12052 0.584493f
C120 a_66329_n6784.t4 a_53801_n12052 0.114506f
C121 a_66329_n6784.n8 a_53801_n12052 1.70971f
C122 OUT.t40 a_53801_n12052 5.03676f
C123 OUT.n2 a_53801_n12052 0.026335f
C124 OUT.n4 a_53801_n12052 0.012185f
C125 OUT.n6 a_53801_n12052 0.012185f
C126 OUT.n8 a_53801_n12052 0.012185f
C127 OUT.n10 a_53801_n12052 0.012185f
C128 OUT.n12 a_53801_n12052 0.012185f
C129 OUT.n14 a_53801_n12052 0.012185f
C130 OUT.n16 a_53801_n12052 0.012185f
C131 OUT.n18 a_53801_n12052 0.01449f
C132 OUT.n19 a_53801_n12052 0.015084f
C133 OUT.n20 a_53801_n12052 0.014538f
C134 OUT.n21 a_53801_n12052 0.066254f
C135 OUT.n22 a_53801_n12052 0.014538f
C136 OUT.n23 a_53801_n12052 0.027312f
C137 OUT.n24 a_53801_n12052 0.014538f
C138 OUT.n25 a_53801_n12052 0.021783f
C139 OUT.n26 a_53801_n12052 0.014982f
C140 OUT.n27 a_53801_n12052 0.014538f
C141 OUT.n28 a_53801_n12052 0.05895f
C142 OUT.n29 a_53801_n12052 0.014538f
C143 OUT.n30 a_53801_n12052 0.027312f
C144 OUT.n31 a_53801_n12052 0.014538f
C145 OUT.n32 a_53801_n12052 0.027312f
C146 OUT.n33 a_53801_n12052 0.014538f
C147 OUT.n34 a_53801_n12052 0.092248f
C148 OUT.n35 a_53801_n12052 0.014538f
C149 OUT.n36 a_53801_n12052 0.0854f
C150 OUT.n37 a_53801_n12052 0.054683f
C151 OUT.n38 a_53801_n12052 0.163471f
C152 OUT.n39 a_53801_n12052 0.902001f
C153 VDD.n0 a_53801_n12052 0.010417f
C154 VDD.t36 a_53801_n12052 0.061714f
C155 VDD.t0 a_53801_n12052 0.038615f
C156 VDD.t1 a_53801_n12052 0.023667f
C157 VDD.n2 a_53801_n12052 0.063941f
C158 VDD.t37 a_53801_n12052 0.023677f
C159 VDD.n3 a_53801_n12052 0.04464f
C160 VDD.n8 a_53801_n12052 0.03146f
C161 VDD.n9 a_53801_n12052 0.074757f
C162 VDD.t34 a_53801_n12052 0.067171f
C163 VDD.t35 a_53801_n12052 0.010712f
C164 VDD.n10 a_53801_n12052 0.079996f
C165 VDD.n11 a_53801_n12052 0.757225f
C166 VDD.t18 a_53801_n12052 0.061714f
C167 VDD.t24 a_53801_n12052 0.032314f
C168 VDD.t42 a_53801_n12052 0.032314f
C169 VDD.t12 a_53801_n12052 0.032314f
C170 VDD.t32 a_53801_n12052 0.032314f
C171 VDD.t30 a_53801_n12052 0.032314f
C172 VDD.t16 a_53801_n12052 0.032314f
C173 VDD.t28 a_53801_n12052 0.032314f
C174 VDD.t44 a_53801_n12052 0.032314f
C175 VDD.t4 a_53801_n12052 0.038306f
C176 VDD.t5 a_53801_n12052 0.021236f
C177 VDD.n12 a_53801_n12052 0.063112f
C178 VDD.n13 a_53801_n12052 0.012f
C179 VDD.n14 a_53801_n12052 0.030188f
C180 VDD.n15 a_53801_n12052 0.012f
C181 VDD.n16 a_53801_n12052 0.028665f
C182 VDD.n17 a_53801_n12052 0.012f
C183 VDD.n18 a_53801_n12052 0.028665f
C184 VDD.n19 a_53801_n12052 0.012f
C185 VDD.n20 a_53801_n12052 0.030243f
C186 VDD.t19 a_53801_n12052 0.021236f
C187 VDD.n21 a_53801_n12052 0.050937f
C188 VDD.t15 a_53801_n12052 0.021596f
C189 VDD.n22 a_53801_n12052 0.012f
C190 VDD.n23 a_53801_n12052 0.050843f
C191 VDD.n24 a_53801_n12052 0.012f
C192 VDD.n25 a_53801_n12052 0.028665f
C193 VDD.n26 a_53801_n12052 0.012f
C194 VDD.n27 a_53801_n12052 0.028665f
C195 VDD.n28 a_53801_n12052 0.012f
C196 VDD.n29 a_53801_n12052 0.030216f
C197 VDD.t9 a_53801_n12052 0.021236f
C198 VDD.n30 a_53801_n12052 0.023038f
C199 VDD.t14 a_53801_n12052 0.061714f
C200 VDD.t20 a_53801_n12052 0.032314f
C201 VDD.t38 a_53801_n12052 0.032314f
C202 VDD.t6 a_53801_n12052 0.032314f
C203 VDD.t2 a_53801_n12052 0.032314f
C204 VDD.t26 a_53801_n12052 0.032314f
C205 VDD.t10 a_53801_n12052 0.032314f
C206 VDD.t22 a_53801_n12052 0.032314f
C207 VDD.t40 a_53801_n12052 0.032314f
C208 VDD.t8 a_53801_n12052 0.038302f
C209 VDD.n31 a_53801_n12052 0.070559f
C210 VDD.n32 a_53801_n12052 0.309878f
C211 VDD.n33 a_53801_n12052 2.77737f
C212 IB.n19 a_53801_n12052 0.023906f
C213 IB.n20 a_53801_n12052 0.387549f
C214 IB.n21 a_53801_n12052 0.456531f
C215 a_61329_n6784.n0 a_53801_n12052 1.0042f
C216 a_61329_n6784.n1 a_53801_n12052 1.15261f
C217 a_61329_n6784.t3 a_53801_n12052 0.029681f
C218 a_61329_n6784.t12 a_53801_n12052 0.10051f
C219 a_61329_n6784.t0 a_53801_n12052 0.089675f
C220 a_61329_n6784.n2 a_53801_n12052 1.12675f
C221 a_61329_n6784.t1 a_53801_n12052 0.204966f
C222 a_61329_n6784.n3 a_53801_n12052 0.613163f
C223 a_61329_n6784.t6 a_53801_n12052 0.029681f
C224 a_61329_n6784.t2 a_53801_n12052 0.029681f
C225 a_61329_n6784.n4 a_53801_n12052 0.14255f
C226 a_61329_n6784.t8 a_53801_n12052 0.029681f
C227 a_61329_n6784.t4 a_53801_n12052 0.029681f
C228 a_61329_n6784.n5 a_53801_n12052 0.141137f
C229 a_61329_n6784.t9 a_53801_n12052 0.029681f
C230 a_61329_n6784.t10 a_53801_n12052 0.029681f
C231 a_61329_n6784.n6 a_53801_n12052 0.141137f
C232 a_61329_n6784.t7 a_53801_n12052 0.029681f
C233 a_61329_n6784.t5 a_53801_n12052 0.029681f
C234 a_61329_n6784.n7 a_53801_n12052 0.145365f
C235 a_61329_n6784.n8 a_53801_n12052 0.141133f
C236 a_61329_n6784.t11 a_53801_n12052 0.029681f
C237 dw_60815_n7004.n0 a_53801_n12052 5.88733f
C238 dw_60815_n7004.t21 a_53801_n12052 0.186518f
C239 dw_60815_n7004.t15 a_53801_n12052 0.186518f
C240 dw_60815_n7004.t13 a_53801_n12052 0.186518f
C241 dw_60815_n7004.t11 a_53801_n12052 0.186518f
C242 dw_60815_n7004.t6 a_53801_n12052 0.186621f
C243 dw_60815_n7004.t4 a_53801_n12052 0.186621f
C244 dw_60815_n7004.t9 a_53801_n12052 0.186621f
C245 dw_60815_n7004.t28 a_53801_n12052 0.276498f
C246 dw_60815_n7004.t1 a_53801_n12052 0.186618f
C247 dw_60815_n7004.n1 a_53801_n12052 1.2724f
C248 dw_60815_n7004.t30 a_53801_n12052 0.644166f
C249 dw_60815_n7004.t5 a_53801_n12052 0.337288f
C250 dw_60815_n7004.t29 a_53801_n12052 0.337288f
C251 dw_60815_n7004.t7 a_53801_n12052 0.337288f
C252 dw_60815_n7004.t3 a_53801_n12052 0.337288f
C253 dw_60815_n7004.t8 a_53801_n12052 0.337288f
C254 dw_60815_n7004.t32 a_53801_n12052 0.337288f
C255 dw_60815_n7004.t0 a_53801_n12052 0.337288f
C256 dw_60815_n7004.t2 a_53801_n12052 0.337288f
C257 dw_60815_n7004.t26 a_53801_n12052 0.399833f
C258 dw_60815_n7004.t27 a_53801_n12052 0.221663f
C259 dw_60815_n7004.t17 a_53801_n12052 0.221663f
C260 dw_60815_n7004.t19 a_53801_n12052 0.221663f
C261 dw_60815_n7004.t16 a_53801_n12052 0.644166f
C262 dw_60815_n7004.t20 a_53801_n12052 0.337288f
C263 dw_60815_n7004.t25 a_53801_n12052 0.337288f
C264 dw_60815_n7004.t14 a_53801_n12052 0.337288f
C265 dw_60815_n7004.t24 a_53801_n12052 0.337288f
C266 dw_60815_n7004.t23 a_53801_n12052 0.337288f
C267 dw_60815_n7004.t12 a_53801_n12052 0.337288f
C268 dw_60815_n7004.t22 a_53801_n12052 0.337288f
C269 dw_60815_n7004.t10 a_53801_n12052 0.337288f
C270 dw_60815_n7004.t18 a_53801_n12052 0.399794f
C271 dw_60815_n7004.t31 a_53801_n12052 0.221663f
C272 VINN.n8 a_53801_n12052 0.011626f
C273 OUT.t40 a_79287_n10784.t2 1.5p
.ends

