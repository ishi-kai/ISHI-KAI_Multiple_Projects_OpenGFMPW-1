* Extracted by KLayout with GF180MCU LVS runset on : 06/12/2023 23:06

.SUBCKT TOP VSS OUT VDD VINN VINP IB
M$1 OUT IB VDD VDD pfet_06v0_dn L=0.7U W=140U AS=43.54P AD=43.54P PS=166.44U
+ PD=166.44U
M$11 \$565 VINP \$1321 \$1321 pfet_06v0_dn L=0.7U W=70U AS=21.77P AD=21.77P
+ PS=83.22U PD=83.22U
M$21 \$633 VINN \$1321 \$1321 pfet_06v0_dn L=0.7U W=70U AS=21.77P AD=21.77P
+ PS=83.22U PD=83.22U
M$41 \$1321 IB VDD VDD pfet_06v0_dn L=0.7U W=14U AS=7.21P AD=7.21P PS=23.06U
+ PD=23.06U
M$43 VDD IB \$566 VDD pfet_06v0_dn L=0.7U W=7U AS=5.39P AD=5.39P PS=15.54U
+ PD=15.54U
M$44 \$335 \$566 \$565 VSS nfet_06v0_dn L=0.7U W=14U AS=5.285P AD=5.285P
+ PS=20.52U PD=20.52U
M$48 \$566 \$566 \$329 VSS nfet_06v0_dn L=0.7U W=3.5U AS=2.555P AD=2.555P
+ PS=8.46U PD=8.46U
M$49 \$565 \$633 VSS VSS nfet_06v0_dn L=0.7U W=3.5U AS=2.555P AD=2.555P
+ PS=8.46U PD=8.46U
M$50 OUT \$565 VSS VSS nfet_06v0_dn L=0.7U W=70U AS=19.845P AD=19.845P
+ PS=84.84U PD=84.84U
M$70 VSS \$329 \$329 VSS nfet_06v0_dn L=0.7U W=3.5U AS=2.555P AD=2.555P
+ PS=8.46U PD=8.46U
M$71 VSS \$633 \$633 VSS nfet_06v0_dn L=0.7U W=3.5U AS=2.555P AD=2.555P
+ PS=8.46U PD=8.46U
C$72 \$335 OUT 1.49994e-12 cap_mim_2f0ff A=749.97P P=116.46U
.ENDS TOP
