* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VSS OUT VINP VDD VINN IB
X0 a_61329_n6784 VINN dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X1 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X2 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X3 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X4 a_66329_n6784 a_55035_n6784 a_79287_n10784 VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X5 VDD IB IB VDD pfet_06v0 ad=5.39p pd=15.539999u as=5.39p ps=15.539999u w=7u l=0.7u
X6 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X7 a_79287_n10784 a_55035_n6784 a_66329_n6784 VSS nfet_06v0 ad=0.91p pd=4.02u as=2.555p ps=8.46u w=3.5u l=0.7u
X8 dw_60815_n7004 VINP a_66329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X9 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X10 a_66329_n6784 VINP dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X11 VSS a_55043_n10784 a_55043_n10784 VSS nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X12 dw_60815_n7004 VINP a_66329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X13 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X14 a_66329_n6784 a_55035_n6784 a_79287_n10784 VSS nfet_06v0 ad=2.555p pd=8.46u as=0.91p ps=4.02u w=3.5u l=0.7u
X15 dw_60815_n7004 VINP a_66329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X16 a_66329_n6784 a_61329_n6784 VSS VSS nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X17 dw_60815_n7004 IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X18 a_61329_n6784 VINN dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X19 dw_60815_n7004 VINN a_61329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X20 dw_60815_n7004 VINN a_61329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X21 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X22 VDD IB a_55035_n6784 VDD pfet_06v0 ad=5.39p pd=15.539999u as=5.39p ps=15.539999u w=7u l=0.7u
X23 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X24 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X25 dw_60815_n7004 VINN a_61329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X26 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X27 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X28 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X29 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X30 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X31 w_62417_n11436 a_61329_n6784 a_61329_n6784 w_62417_n11436 nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X32 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X33 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X34 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X35 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X36 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X37 dw_60815_n7004 VINP a_66329_n6784 dw_60815_n7004 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X38 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X39 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X40 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X41 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X42 a_66329_n6784 VINP dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X43 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X44 a_66329_n6784 VINP dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X45 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X46 OUT a_79287_n10784 cap_mim_2f0_m4m5_noshield c_width=39u c_length=19.23u
X47 dw_60815_n7004 VINN a_61329_n6784 dw_60815_n7004 pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X48 a_79287_n10784 a_55035_n6784 a_66329_n6784 VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X49 a_61329_n6784 VINN dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X50 dw_60815_n7004 VINP a_66329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X51 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=2.555p ps=8.46u w=3.5u l=0.7u
X52 a_61329_n6784 VINN dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X53 VDD IB OUT VDD pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X54 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X55 dw_60815_n7004 VINN a_61329_n6784 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X56 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X57 VDD IB OUT VDD pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X58 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=2.555p pd=8.46u as=0.91p ps=4.02u w=3.5u l=0.7u
X59 a_66329_n6784 VINP dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X60 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=5.39p ps=15.539999u w=7u l=0.7u
X61 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X62 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X63 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X64 OUT IB VDD VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X65 a_66329_n6784 VINP dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X66 a_61329_n6784 VINN dw_60815_n7004 dw_60815_n7004 pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X67 VDD IB OUT VDD pfet_06v0 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.7u
X68 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X69 VSS a_66329_n6784 OUT VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X70 VDD IB dw_60815_n7004 VDD pfet_06v0 ad=5.39p pd=15.539999u as=1.82p ps=7.52u w=7u l=0.7u
X71 a_55035_n6784 a_55035_n6784 a_55043_n10784 VSS nfet_06v0 ad=2.555p pd=8.46u as=2.555p ps=8.46u w=3.5u l=0.7u
X72 OUT a_66329_n6784 VSS VSS nfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
.ends

