magic
tech gf180mcuD
magscale 1 10
timestamp 1699608903
<< metal1 >>
rect 1344 36874 78624 36908
rect 1344 36822 10874 36874
rect 10926 36822 10978 36874
rect 11030 36822 11082 36874
rect 11134 36822 30194 36874
rect 30246 36822 30298 36874
rect 30350 36822 30402 36874
rect 30454 36822 49514 36874
rect 49566 36822 49618 36874
rect 49670 36822 49722 36874
rect 49774 36822 68834 36874
rect 68886 36822 68938 36874
rect 68990 36822 69042 36874
rect 69094 36822 78624 36874
rect 1344 36788 78624 36822
rect 1344 36090 78784 36124
rect 1344 36038 20534 36090
rect 20586 36038 20638 36090
rect 20690 36038 20742 36090
rect 20794 36038 39854 36090
rect 39906 36038 39958 36090
rect 40010 36038 40062 36090
rect 40114 36038 59174 36090
rect 59226 36038 59278 36090
rect 59330 36038 59382 36090
rect 59434 36038 78494 36090
rect 78546 36038 78598 36090
rect 78650 36038 78702 36090
rect 78754 36038 78784 36090
rect 1344 36004 78784 36038
rect 1344 35306 78624 35340
rect 1344 35254 10874 35306
rect 10926 35254 10978 35306
rect 11030 35254 11082 35306
rect 11134 35254 30194 35306
rect 30246 35254 30298 35306
rect 30350 35254 30402 35306
rect 30454 35254 49514 35306
rect 49566 35254 49618 35306
rect 49670 35254 49722 35306
rect 49774 35254 68834 35306
rect 68886 35254 68938 35306
rect 68990 35254 69042 35306
rect 69094 35254 78624 35306
rect 1344 35220 78624 35254
rect 1344 34522 78784 34556
rect 1344 34470 20534 34522
rect 20586 34470 20638 34522
rect 20690 34470 20742 34522
rect 20794 34470 39854 34522
rect 39906 34470 39958 34522
rect 40010 34470 40062 34522
rect 40114 34470 59174 34522
rect 59226 34470 59278 34522
rect 59330 34470 59382 34522
rect 59434 34470 78494 34522
rect 78546 34470 78598 34522
rect 78650 34470 78702 34522
rect 78754 34470 78784 34522
rect 1344 34436 78784 34470
rect 1344 33738 78624 33772
rect 1344 33686 10874 33738
rect 10926 33686 10978 33738
rect 11030 33686 11082 33738
rect 11134 33686 30194 33738
rect 30246 33686 30298 33738
rect 30350 33686 30402 33738
rect 30454 33686 49514 33738
rect 49566 33686 49618 33738
rect 49670 33686 49722 33738
rect 49774 33686 68834 33738
rect 68886 33686 68938 33738
rect 68990 33686 69042 33738
rect 69094 33686 78624 33738
rect 1344 33652 78624 33686
rect 1344 32954 78784 32988
rect 1344 32902 20534 32954
rect 20586 32902 20638 32954
rect 20690 32902 20742 32954
rect 20794 32902 39854 32954
rect 39906 32902 39958 32954
rect 40010 32902 40062 32954
rect 40114 32902 59174 32954
rect 59226 32902 59278 32954
rect 59330 32902 59382 32954
rect 59434 32902 78494 32954
rect 78546 32902 78598 32954
rect 78650 32902 78702 32954
rect 78754 32902 78784 32954
rect 1344 32868 78784 32902
rect 1344 32170 78624 32204
rect 1344 32118 10874 32170
rect 10926 32118 10978 32170
rect 11030 32118 11082 32170
rect 11134 32118 30194 32170
rect 30246 32118 30298 32170
rect 30350 32118 30402 32170
rect 30454 32118 49514 32170
rect 49566 32118 49618 32170
rect 49670 32118 49722 32170
rect 49774 32118 68834 32170
rect 68886 32118 68938 32170
rect 68990 32118 69042 32170
rect 69094 32118 78624 32170
rect 1344 32084 78624 32118
rect 1344 31386 78784 31420
rect 1344 31334 20534 31386
rect 20586 31334 20638 31386
rect 20690 31334 20742 31386
rect 20794 31334 39854 31386
rect 39906 31334 39958 31386
rect 40010 31334 40062 31386
rect 40114 31334 59174 31386
rect 59226 31334 59278 31386
rect 59330 31334 59382 31386
rect 59434 31334 78494 31386
rect 78546 31334 78598 31386
rect 78650 31334 78702 31386
rect 78754 31334 78784 31386
rect 1344 31300 78784 31334
rect 1344 30602 78624 30636
rect 1344 30550 10874 30602
rect 10926 30550 10978 30602
rect 11030 30550 11082 30602
rect 11134 30550 30194 30602
rect 30246 30550 30298 30602
rect 30350 30550 30402 30602
rect 30454 30550 49514 30602
rect 49566 30550 49618 30602
rect 49670 30550 49722 30602
rect 49774 30550 68834 30602
rect 68886 30550 68938 30602
rect 68990 30550 69042 30602
rect 69094 30550 78624 30602
rect 1344 30516 78624 30550
rect 1344 29818 78784 29852
rect 1344 29766 20534 29818
rect 20586 29766 20638 29818
rect 20690 29766 20742 29818
rect 20794 29766 39854 29818
rect 39906 29766 39958 29818
rect 40010 29766 40062 29818
rect 40114 29766 59174 29818
rect 59226 29766 59278 29818
rect 59330 29766 59382 29818
rect 59434 29766 78494 29818
rect 78546 29766 78598 29818
rect 78650 29766 78702 29818
rect 78754 29766 78784 29818
rect 1344 29732 78784 29766
rect 1344 29034 78624 29068
rect 1344 28982 10874 29034
rect 10926 28982 10978 29034
rect 11030 28982 11082 29034
rect 11134 28982 30194 29034
rect 30246 28982 30298 29034
rect 30350 28982 30402 29034
rect 30454 28982 49514 29034
rect 49566 28982 49618 29034
rect 49670 28982 49722 29034
rect 49774 28982 68834 29034
rect 68886 28982 68938 29034
rect 68990 28982 69042 29034
rect 69094 28982 78624 29034
rect 1344 28948 78624 28982
rect 1344 28250 78784 28284
rect 1344 28198 20534 28250
rect 20586 28198 20638 28250
rect 20690 28198 20742 28250
rect 20794 28198 39854 28250
rect 39906 28198 39958 28250
rect 40010 28198 40062 28250
rect 40114 28198 59174 28250
rect 59226 28198 59278 28250
rect 59330 28198 59382 28250
rect 59434 28198 78494 28250
rect 78546 28198 78598 28250
rect 78650 28198 78702 28250
rect 78754 28198 78784 28250
rect 1344 28164 78784 28198
rect 1344 27466 78624 27500
rect 1344 27414 10874 27466
rect 10926 27414 10978 27466
rect 11030 27414 11082 27466
rect 11134 27414 30194 27466
rect 30246 27414 30298 27466
rect 30350 27414 30402 27466
rect 30454 27414 49514 27466
rect 49566 27414 49618 27466
rect 49670 27414 49722 27466
rect 49774 27414 68834 27466
rect 68886 27414 68938 27466
rect 68990 27414 69042 27466
rect 69094 27414 78624 27466
rect 1344 27380 78624 27414
rect 1344 26682 78784 26716
rect 1344 26630 20534 26682
rect 20586 26630 20638 26682
rect 20690 26630 20742 26682
rect 20794 26630 39854 26682
rect 39906 26630 39958 26682
rect 40010 26630 40062 26682
rect 40114 26630 59174 26682
rect 59226 26630 59278 26682
rect 59330 26630 59382 26682
rect 59434 26630 78494 26682
rect 78546 26630 78598 26682
rect 78650 26630 78702 26682
rect 78754 26630 78784 26682
rect 1344 26596 78784 26630
rect 1344 25898 78624 25932
rect 1344 25846 10874 25898
rect 10926 25846 10978 25898
rect 11030 25846 11082 25898
rect 11134 25846 30194 25898
rect 30246 25846 30298 25898
rect 30350 25846 30402 25898
rect 30454 25846 49514 25898
rect 49566 25846 49618 25898
rect 49670 25846 49722 25898
rect 49774 25846 68834 25898
rect 68886 25846 68938 25898
rect 68990 25846 69042 25898
rect 69094 25846 78624 25898
rect 1344 25812 78624 25846
rect 1344 25114 78784 25148
rect 1344 25062 20534 25114
rect 20586 25062 20638 25114
rect 20690 25062 20742 25114
rect 20794 25062 39854 25114
rect 39906 25062 39958 25114
rect 40010 25062 40062 25114
rect 40114 25062 59174 25114
rect 59226 25062 59278 25114
rect 59330 25062 59382 25114
rect 59434 25062 78494 25114
rect 78546 25062 78598 25114
rect 78650 25062 78702 25114
rect 78754 25062 78784 25114
rect 1344 25028 78784 25062
rect 1344 24330 78624 24364
rect 1344 24278 10874 24330
rect 10926 24278 10978 24330
rect 11030 24278 11082 24330
rect 11134 24278 30194 24330
rect 30246 24278 30298 24330
rect 30350 24278 30402 24330
rect 30454 24278 49514 24330
rect 49566 24278 49618 24330
rect 49670 24278 49722 24330
rect 49774 24278 68834 24330
rect 68886 24278 68938 24330
rect 68990 24278 69042 24330
rect 69094 24278 78624 24330
rect 1344 24244 78624 24278
rect 1344 23546 78784 23580
rect 1344 23494 20534 23546
rect 20586 23494 20638 23546
rect 20690 23494 20742 23546
rect 20794 23494 39854 23546
rect 39906 23494 39958 23546
rect 40010 23494 40062 23546
rect 40114 23494 59174 23546
rect 59226 23494 59278 23546
rect 59330 23494 59382 23546
rect 59434 23494 78494 23546
rect 78546 23494 78598 23546
rect 78650 23494 78702 23546
rect 78754 23494 78784 23546
rect 1344 23460 78784 23494
rect 1344 22762 78624 22796
rect 1344 22710 10874 22762
rect 10926 22710 10978 22762
rect 11030 22710 11082 22762
rect 11134 22710 30194 22762
rect 30246 22710 30298 22762
rect 30350 22710 30402 22762
rect 30454 22710 49514 22762
rect 49566 22710 49618 22762
rect 49670 22710 49722 22762
rect 49774 22710 68834 22762
rect 68886 22710 68938 22762
rect 68990 22710 69042 22762
rect 69094 22710 78624 22762
rect 1344 22676 78624 22710
rect 1344 21978 78784 22012
rect 1344 21926 20534 21978
rect 20586 21926 20638 21978
rect 20690 21926 20742 21978
rect 20794 21926 39854 21978
rect 39906 21926 39958 21978
rect 40010 21926 40062 21978
rect 40114 21926 59174 21978
rect 59226 21926 59278 21978
rect 59330 21926 59382 21978
rect 59434 21926 78494 21978
rect 78546 21926 78598 21978
rect 78650 21926 78702 21978
rect 78754 21926 78784 21978
rect 1344 21892 78784 21926
rect 1344 21194 78624 21228
rect 1344 21142 10874 21194
rect 10926 21142 10978 21194
rect 11030 21142 11082 21194
rect 11134 21142 30194 21194
rect 30246 21142 30298 21194
rect 30350 21142 30402 21194
rect 30454 21142 49514 21194
rect 49566 21142 49618 21194
rect 49670 21142 49722 21194
rect 49774 21142 68834 21194
rect 68886 21142 68938 21194
rect 68990 21142 69042 21194
rect 69094 21142 78624 21194
rect 1344 21108 78624 21142
rect 1344 20410 78784 20444
rect 1344 20358 20534 20410
rect 20586 20358 20638 20410
rect 20690 20358 20742 20410
rect 20794 20358 39854 20410
rect 39906 20358 39958 20410
rect 40010 20358 40062 20410
rect 40114 20358 59174 20410
rect 59226 20358 59278 20410
rect 59330 20358 59382 20410
rect 59434 20358 78494 20410
rect 78546 20358 78598 20410
rect 78650 20358 78702 20410
rect 78754 20358 78784 20410
rect 1344 20324 78784 20358
rect 1344 19626 78624 19660
rect 1344 19574 10874 19626
rect 10926 19574 10978 19626
rect 11030 19574 11082 19626
rect 11134 19574 30194 19626
rect 30246 19574 30298 19626
rect 30350 19574 30402 19626
rect 30454 19574 49514 19626
rect 49566 19574 49618 19626
rect 49670 19574 49722 19626
rect 49774 19574 68834 19626
rect 68886 19574 68938 19626
rect 68990 19574 69042 19626
rect 69094 19574 78624 19626
rect 1344 19540 78624 19574
rect 1344 18842 78784 18876
rect 1344 18790 20534 18842
rect 20586 18790 20638 18842
rect 20690 18790 20742 18842
rect 20794 18790 39854 18842
rect 39906 18790 39958 18842
rect 40010 18790 40062 18842
rect 40114 18790 59174 18842
rect 59226 18790 59278 18842
rect 59330 18790 59382 18842
rect 59434 18790 78494 18842
rect 78546 18790 78598 18842
rect 78650 18790 78702 18842
rect 78754 18790 78784 18842
rect 1344 18756 78784 18790
rect 1344 18058 78624 18092
rect 1344 18006 10874 18058
rect 10926 18006 10978 18058
rect 11030 18006 11082 18058
rect 11134 18006 30194 18058
rect 30246 18006 30298 18058
rect 30350 18006 30402 18058
rect 30454 18006 49514 18058
rect 49566 18006 49618 18058
rect 49670 18006 49722 18058
rect 49774 18006 68834 18058
rect 68886 18006 68938 18058
rect 68990 18006 69042 18058
rect 69094 18006 78624 18058
rect 1344 17972 78624 18006
rect 1344 17274 78784 17308
rect 1344 17222 20534 17274
rect 20586 17222 20638 17274
rect 20690 17222 20742 17274
rect 20794 17222 39854 17274
rect 39906 17222 39958 17274
rect 40010 17222 40062 17274
rect 40114 17222 59174 17274
rect 59226 17222 59278 17274
rect 59330 17222 59382 17274
rect 59434 17222 78494 17274
rect 78546 17222 78598 17274
rect 78650 17222 78702 17274
rect 78754 17222 78784 17274
rect 1344 17188 78784 17222
rect 1344 16490 78624 16524
rect 1344 16438 10874 16490
rect 10926 16438 10978 16490
rect 11030 16438 11082 16490
rect 11134 16438 30194 16490
rect 30246 16438 30298 16490
rect 30350 16438 30402 16490
rect 30454 16438 49514 16490
rect 49566 16438 49618 16490
rect 49670 16438 49722 16490
rect 49774 16438 68834 16490
rect 68886 16438 68938 16490
rect 68990 16438 69042 16490
rect 69094 16438 78624 16490
rect 1344 16404 78624 16438
rect 1344 15706 78784 15740
rect 1344 15654 20534 15706
rect 20586 15654 20638 15706
rect 20690 15654 20742 15706
rect 20794 15654 39854 15706
rect 39906 15654 39958 15706
rect 40010 15654 40062 15706
rect 40114 15654 59174 15706
rect 59226 15654 59278 15706
rect 59330 15654 59382 15706
rect 59434 15654 78494 15706
rect 78546 15654 78598 15706
rect 78650 15654 78702 15706
rect 78754 15654 78784 15706
rect 1344 15620 78784 15654
rect 35746 15374 35758 15426
rect 35810 15374 35822 15426
rect 34738 15150 34750 15202
rect 34802 15150 34814 15202
rect 1344 14922 78624 14956
rect 1344 14870 10874 14922
rect 10926 14870 10978 14922
rect 11030 14870 11082 14922
rect 11134 14870 30194 14922
rect 30246 14870 30298 14922
rect 30350 14870 30402 14922
rect 30454 14870 49514 14922
rect 49566 14870 49618 14922
rect 49670 14870 49722 14922
rect 49774 14870 68834 14922
rect 68886 14870 68938 14922
rect 68990 14870 69042 14922
rect 69094 14870 78624 14922
rect 1344 14836 78624 14870
rect 34850 14590 34862 14642
rect 34914 14590 34926 14642
rect 37326 14418 37378 14430
rect 33842 14366 33854 14418
rect 33906 14366 33918 14418
rect 37326 14354 37378 14366
rect 38110 14418 38162 14430
rect 38110 14354 38162 14366
rect 37102 14306 37154 14318
rect 37102 14242 37154 14254
rect 37214 14306 37266 14318
rect 37214 14242 37266 14254
rect 37998 14306 38050 14318
rect 37998 14242 38050 14254
rect 38558 14306 38610 14318
rect 38558 14242 38610 14254
rect 1344 14138 78784 14172
rect 1344 14086 20534 14138
rect 20586 14086 20638 14138
rect 20690 14086 20742 14138
rect 20794 14086 39854 14138
rect 39906 14086 39958 14138
rect 40010 14086 40062 14138
rect 40114 14086 59174 14138
rect 59226 14086 59278 14138
rect 59330 14086 59382 14138
rect 59434 14086 78494 14138
rect 78546 14086 78598 14138
rect 78650 14086 78702 14138
rect 78754 14086 78784 14138
rect 1344 14052 78784 14086
rect 34526 13858 34578 13870
rect 35298 13806 35310 13858
rect 35362 13806 35374 13858
rect 39890 13806 39902 13858
rect 39954 13806 39966 13858
rect 34526 13794 34578 13806
rect 13246 13634 13298 13646
rect 13246 13570 13298 13582
rect 32174 13634 32226 13646
rect 32174 13570 32226 13582
rect 32510 13634 32562 13646
rect 32510 13570 32562 13582
rect 33182 13634 33234 13646
rect 33182 13570 33234 13582
rect 33742 13634 33794 13646
rect 33742 13570 33794 13582
rect 34638 13634 34690 13646
rect 41134 13634 41186 13646
rect 36306 13582 36318 13634
rect 36370 13582 36382 13634
rect 38882 13582 38894 13634
rect 38946 13582 38958 13634
rect 34638 13570 34690 13582
rect 41134 13570 41186 13582
rect 34750 13522 34802 13534
rect 31938 13470 31950 13522
rect 32002 13519 32014 13522
rect 32498 13519 32510 13522
rect 32002 13473 32510 13519
rect 32002 13470 32014 13473
rect 32498 13470 32510 13473
rect 32562 13470 32574 13522
rect 34750 13458 34802 13470
rect 1344 13354 78624 13388
rect 1344 13302 10874 13354
rect 10926 13302 10978 13354
rect 11030 13302 11082 13354
rect 11134 13302 30194 13354
rect 30246 13302 30298 13354
rect 30350 13302 30402 13354
rect 30454 13302 49514 13354
rect 49566 13302 49618 13354
rect 49670 13302 49722 13354
rect 49774 13302 68834 13354
rect 68886 13302 68938 13354
rect 68990 13302 69042 13354
rect 69094 13302 78624 13354
rect 1344 13268 78624 13302
rect 39902 13074 39954 13086
rect 12898 13022 12910 13074
rect 12962 13022 12974 13074
rect 33506 13022 33518 13074
rect 33570 13022 33582 13074
rect 35634 13022 35646 13074
rect 35698 13022 35710 13074
rect 37762 13022 37774 13074
rect 37826 13022 37838 13074
rect 46162 13022 46174 13074
rect 46226 13022 46238 13074
rect 39902 13010 39954 13022
rect 31950 12962 32002 12974
rect 10098 12910 10110 12962
rect 10162 12910 10174 12962
rect 13570 12910 13582 12962
rect 13634 12910 13646 12962
rect 19394 12910 19406 12962
rect 19458 12910 19470 12962
rect 36306 12910 36318 12962
rect 36370 12910 36382 12962
rect 36978 12910 36990 12962
rect 37042 12910 37054 12962
rect 31950 12898 32002 12910
rect 41246 12850 41298 12862
rect 10770 12798 10782 12850
rect 10834 12798 10846 12850
rect 41246 12786 41298 12798
rect 41358 12850 41410 12862
rect 47506 12798 47518 12850
rect 47570 12798 47582 12850
rect 41358 12786 41410 12798
rect 13806 12738 13858 12750
rect 13806 12674 13858 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 20862 12738 20914 12750
rect 20862 12674 20914 12686
rect 21758 12738 21810 12750
rect 21758 12674 21810 12686
rect 22878 12738 22930 12750
rect 22878 12674 22930 12686
rect 23662 12738 23714 12750
rect 23662 12674 23714 12686
rect 24110 12738 24162 12750
rect 24110 12674 24162 12686
rect 24446 12738 24498 12750
rect 24446 12674 24498 12686
rect 25006 12738 25058 12750
rect 25006 12674 25058 12686
rect 25342 12738 25394 12750
rect 25342 12674 25394 12686
rect 25902 12738 25954 12750
rect 25902 12674 25954 12686
rect 26686 12738 26738 12750
rect 26686 12674 26738 12686
rect 27134 12738 27186 12750
rect 27134 12674 27186 12686
rect 27582 12738 27634 12750
rect 27582 12674 27634 12686
rect 30494 12738 30546 12750
rect 30494 12674 30546 12686
rect 31054 12738 31106 12750
rect 31054 12674 31106 12686
rect 31726 12738 31778 12750
rect 31726 12674 31778 12686
rect 32510 12738 32562 12750
rect 32510 12674 32562 12686
rect 33294 12738 33346 12750
rect 40798 12738 40850 12750
rect 40450 12686 40462 12738
rect 40514 12686 40526 12738
rect 33294 12674 33346 12686
rect 40798 12674 40850 12686
rect 41582 12738 41634 12750
rect 41582 12674 41634 12686
rect 42030 12738 42082 12750
rect 42030 12674 42082 12686
rect 42478 12738 42530 12750
rect 42478 12674 42530 12686
rect 42814 12738 42866 12750
rect 42814 12674 42866 12686
rect 45166 12738 45218 12750
rect 45166 12674 45218 12686
rect 45614 12738 45666 12750
rect 45614 12674 45666 12686
rect 48078 12738 48130 12750
rect 48078 12674 48130 12686
rect 48638 12738 48690 12750
rect 48638 12674 48690 12686
rect 1344 12570 78784 12604
rect 1344 12518 20534 12570
rect 20586 12518 20638 12570
rect 20690 12518 20742 12570
rect 20794 12518 39854 12570
rect 39906 12518 39958 12570
rect 40010 12518 40062 12570
rect 40114 12518 59174 12570
rect 59226 12518 59278 12570
rect 59330 12518 59382 12570
rect 59434 12518 78494 12570
rect 78546 12518 78598 12570
rect 78650 12518 78702 12570
rect 78754 12518 78784 12570
rect 1344 12484 78784 12518
rect 11230 12402 11282 12414
rect 11230 12338 11282 12350
rect 22542 12402 22594 12414
rect 22542 12338 22594 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 27358 12402 27410 12414
rect 27358 12338 27410 12350
rect 33406 12402 33458 12414
rect 33406 12338 33458 12350
rect 40238 12402 40290 12414
rect 40238 12338 40290 12350
rect 31838 12290 31890 12302
rect 12898 12238 12910 12290
rect 12962 12238 12974 12290
rect 14354 12238 14366 12290
rect 14418 12238 14430 12290
rect 20290 12238 20302 12290
rect 20354 12238 20366 12290
rect 23538 12238 23550 12290
rect 23602 12238 23614 12290
rect 29362 12238 29374 12290
rect 29426 12238 29438 12290
rect 31838 12226 31890 12238
rect 32286 12290 32338 12302
rect 32286 12226 32338 12238
rect 32510 12290 32562 12302
rect 48750 12290 48802 12302
rect 44034 12238 44046 12290
rect 44098 12238 44110 12290
rect 45602 12238 45614 12290
rect 45666 12238 45678 12290
rect 32510 12226 32562 12238
rect 48750 12226 48802 12238
rect 49310 12290 49362 12302
rect 49310 12226 49362 12238
rect 11566 12178 11618 12190
rect 11566 12114 11618 12126
rect 12014 12178 12066 12190
rect 17502 12178 17554 12190
rect 24222 12178 24274 12190
rect 40350 12178 40402 12190
rect 13122 12126 13134 12178
rect 13186 12126 13198 12178
rect 13682 12126 13694 12178
rect 13746 12126 13758 12178
rect 20962 12126 20974 12178
rect 21026 12126 21038 12178
rect 23650 12126 23662 12178
rect 23714 12126 23726 12178
rect 33170 12126 33182 12178
rect 33234 12126 33246 12178
rect 37650 12126 37662 12178
rect 37714 12126 37726 12178
rect 39890 12126 39902 12178
rect 39954 12126 39966 12178
rect 44706 12126 44718 12178
rect 44770 12126 44782 12178
rect 12014 12114 12066 12126
rect 17502 12114 17554 12126
rect 24222 12114 24274 12126
rect 40350 12114 40402 12126
rect 21534 12066 21586 12078
rect 16482 12014 16494 12066
rect 16546 12014 16558 12066
rect 18162 12014 18174 12066
rect 18226 12014 18238 12066
rect 21534 12002 21586 12014
rect 22206 12066 22258 12078
rect 22206 12002 22258 12014
rect 23102 12066 23154 12078
rect 23102 12002 23154 12014
rect 25790 12066 25842 12078
rect 25790 12002 25842 12014
rect 26238 12066 26290 12078
rect 26238 12002 26290 12014
rect 26686 12066 26738 12078
rect 26686 12002 26738 12014
rect 27918 12066 27970 12078
rect 27918 12002 27970 12014
rect 28366 12066 28418 12078
rect 28366 12002 28418 12014
rect 28814 12066 28866 12078
rect 31390 12066 31442 12078
rect 30594 12014 30606 12066
rect 30658 12014 30670 12066
rect 28814 12002 28866 12014
rect 31390 12002 31442 12014
rect 32398 12066 32450 12078
rect 41246 12066 41298 12078
rect 47742 12066 47794 12078
rect 35298 12014 35310 12066
rect 35362 12014 35374 12066
rect 40898 12014 40910 12066
rect 40962 12014 40974 12066
rect 41794 12014 41806 12066
rect 41858 12014 41870 12066
rect 32398 12002 32450 12014
rect 41246 12002 41298 12014
rect 47742 12002 47794 12014
rect 49870 12066 49922 12078
rect 49870 12002 49922 12014
rect 50318 12066 50370 12078
rect 50318 12002 50370 12014
rect 50878 12066 50930 12078
rect 50878 12002 50930 12014
rect 12350 11954 12402 11966
rect 12350 11890 12402 11902
rect 24558 11954 24610 11966
rect 33518 11954 33570 11966
rect 31378 11902 31390 11954
rect 31442 11951 31454 11954
rect 31826 11951 31838 11954
rect 31442 11905 31838 11951
rect 31442 11902 31454 11905
rect 31826 11902 31838 11905
rect 31890 11902 31902 11954
rect 24558 11890 24610 11902
rect 33518 11890 33570 11902
rect 39566 11954 39618 11966
rect 39566 11890 39618 11902
rect 39902 11954 39954 11966
rect 39902 11890 39954 11902
rect 1344 11786 78624 11820
rect 1344 11734 10874 11786
rect 10926 11734 10978 11786
rect 11030 11734 11082 11786
rect 11134 11734 30194 11786
rect 30246 11734 30298 11786
rect 30350 11734 30402 11786
rect 30454 11734 49514 11786
rect 49566 11734 49618 11786
rect 49670 11734 49722 11786
rect 49774 11734 68834 11786
rect 68886 11734 68938 11786
rect 68990 11734 69042 11786
rect 69094 11734 78624 11786
rect 1344 11700 78624 11734
rect 14142 11618 14194 11630
rect 14142 11554 14194 11566
rect 19518 11618 19570 11630
rect 69010 11566 69022 11618
rect 69074 11615 69086 11618
rect 70466 11615 70478 11618
rect 69074 11569 70478 11615
rect 69074 11566 69086 11569
rect 70466 11566 70478 11569
rect 70530 11566 70542 11618
rect 19518 11554 19570 11566
rect 28254 11506 28306 11518
rect 23426 11454 23438 11506
rect 23490 11454 23502 11506
rect 28254 11442 28306 11454
rect 29374 11506 29426 11518
rect 29374 11442 29426 11454
rect 33518 11506 33570 11518
rect 33518 11442 33570 11454
rect 38110 11506 38162 11518
rect 38110 11442 38162 11454
rect 43262 11506 43314 11518
rect 49646 11506 49698 11518
rect 46162 11454 46174 11506
rect 46226 11454 46238 11506
rect 43262 11442 43314 11454
rect 49646 11442 49698 11454
rect 50094 11506 50146 11518
rect 50530 11454 50542 11506
rect 50594 11454 50606 11506
rect 50094 11442 50146 11454
rect 14478 11394 14530 11406
rect 14478 11330 14530 11342
rect 19854 11394 19906 11406
rect 36990 11394 37042 11406
rect 20626 11342 20638 11394
rect 20690 11342 20702 11394
rect 26226 11342 26238 11394
rect 26290 11342 26302 11394
rect 32834 11342 32846 11394
rect 32898 11342 32910 11394
rect 36306 11342 36318 11394
rect 36370 11342 36382 11394
rect 19854 11330 19906 11342
rect 36990 11330 37042 11342
rect 37214 11394 37266 11406
rect 43150 11394 43202 11406
rect 37874 11342 37886 11394
rect 37938 11342 37950 11394
rect 41682 11342 41694 11394
rect 41746 11342 41758 11394
rect 42354 11342 42366 11394
rect 42418 11342 42430 11394
rect 37214 11330 37266 11342
rect 43150 11330 43202 11342
rect 43486 11394 43538 11406
rect 43486 11330 43538 11342
rect 44382 11394 44434 11406
rect 69022 11394 69074 11406
rect 49186 11342 49198 11394
rect 49250 11342 49262 11394
rect 44382 11330 44434 11342
rect 69022 11330 69074 11342
rect 22206 11282 22258 11294
rect 29486 11282 29538 11294
rect 38222 11282 38274 11294
rect 42814 11282 42866 11294
rect 14690 11230 14702 11282
rect 14754 11230 14766 11282
rect 15138 11230 15150 11282
rect 15202 11230 15214 11282
rect 20402 11230 20414 11282
rect 20466 11230 20478 11282
rect 25554 11230 25566 11282
rect 25618 11230 25630 11282
rect 32162 11230 32174 11282
rect 32226 11230 32238 11282
rect 35634 11230 35646 11282
rect 35698 11230 35710 11282
rect 41010 11230 41022 11282
rect 41074 11230 41086 11282
rect 22206 11218 22258 11230
rect 29486 11218 29538 11230
rect 38222 11218 38274 11230
rect 42814 11218 42866 11230
rect 43710 11282 43762 11294
rect 43710 11218 43762 11230
rect 43934 11282 43986 11294
rect 43934 11218 43986 11230
rect 44830 11282 44882 11294
rect 48402 11230 48414 11282
rect 48466 11230 48478 11282
rect 51538 11230 51550 11282
rect 51602 11230 51614 11282
rect 44830 11218 44882 11230
rect 12238 11170 12290 11182
rect 12238 11106 12290 11118
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 15822 11170 15874 11182
rect 15822 11106 15874 11118
rect 17726 11170 17778 11182
rect 17726 11106 17778 11118
rect 18286 11170 18338 11182
rect 18286 11106 18338 11118
rect 18846 11170 18898 11182
rect 18846 11106 18898 11118
rect 21422 11170 21474 11182
rect 21422 11106 21474 11118
rect 21870 11170 21922 11182
rect 21870 11106 21922 11118
rect 22766 11170 22818 11182
rect 22766 11106 22818 11118
rect 23102 11170 23154 11182
rect 23102 11106 23154 11118
rect 26798 11170 26850 11182
rect 26798 11106 26850 11118
rect 27246 11170 27298 11182
rect 27246 11106 27298 11118
rect 27806 11170 27858 11182
rect 27806 11106 27858 11118
rect 28590 11170 28642 11182
rect 28590 11106 28642 11118
rect 29262 11170 29314 11182
rect 44158 11170 44210 11182
rect 29922 11118 29934 11170
rect 29986 11118 29998 11170
rect 37538 11118 37550 11170
rect 37602 11118 37614 11170
rect 38770 11118 38782 11170
rect 38834 11118 38846 11170
rect 42130 11118 42142 11170
rect 42194 11118 42206 11170
rect 29262 11106 29314 11118
rect 44158 11106 44210 11118
rect 44942 11170 44994 11182
rect 44942 11106 44994 11118
rect 45166 11170 45218 11182
rect 45166 11106 45218 11118
rect 45390 11170 45442 11182
rect 45390 11106 45442 11118
rect 68574 11170 68626 11182
rect 68574 11106 68626 11118
rect 69470 11170 69522 11182
rect 69470 11106 69522 11118
rect 69918 11170 69970 11182
rect 69918 11106 69970 11118
rect 70366 11170 70418 11182
rect 70366 11106 70418 11118
rect 70702 11170 70754 11182
rect 70702 11106 70754 11118
rect 71262 11170 71314 11182
rect 71262 11106 71314 11118
rect 71710 11170 71762 11182
rect 71710 11106 71762 11118
rect 72158 11170 72210 11182
rect 72158 11106 72210 11118
rect 72494 11170 72546 11182
rect 72494 11106 72546 11118
rect 72942 11170 72994 11182
rect 72942 11106 72994 11118
rect 73838 11170 73890 11182
rect 73838 11106 73890 11118
rect 1344 11002 78784 11036
rect 1344 10950 20534 11002
rect 20586 10950 20638 11002
rect 20690 10950 20742 11002
rect 20794 10950 39854 11002
rect 39906 10950 39958 11002
rect 40010 10950 40062 11002
rect 40114 10950 59174 11002
rect 59226 10950 59278 11002
rect 59330 10950 59382 11002
rect 59434 10950 78494 11002
rect 78546 10950 78598 11002
rect 78650 10950 78702 11002
rect 78754 10950 78784 11002
rect 1344 10916 78784 10950
rect 16942 10834 16994 10846
rect 16942 10770 16994 10782
rect 17950 10834 18002 10846
rect 17950 10770 18002 10782
rect 25566 10834 25618 10846
rect 33854 10834 33906 10846
rect 33394 10782 33406 10834
rect 33458 10782 33470 10834
rect 25566 10770 25618 10782
rect 33854 10770 33906 10782
rect 47854 10834 47906 10846
rect 47854 10770 47906 10782
rect 76974 10834 77026 10846
rect 76974 10770 77026 10782
rect 25230 10722 25282 10734
rect 21074 10670 21086 10722
rect 21138 10670 21150 10722
rect 25230 10658 25282 10670
rect 25902 10722 25954 10734
rect 31726 10722 31778 10734
rect 39342 10722 39394 10734
rect 30146 10670 30158 10722
rect 30210 10670 30222 10722
rect 36082 10670 36094 10722
rect 36146 10670 36158 10722
rect 38658 10670 38670 10722
rect 38722 10670 38734 10722
rect 25902 10658 25954 10670
rect 31726 10658 31778 10670
rect 39342 10658 39394 10670
rect 39790 10722 39842 10734
rect 51550 10722 51602 10734
rect 48178 10670 48190 10722
rect 48242 10670 48254 10722
rect 50754 10670 50766 10722
rect 50818 10670 50830 10722
rect 39790 10658 39842 10670
rect 51550 10658 51602 10670
rect 51998 10722 52050 10734
rect 51998 10658 52050 10670
rect 70254 10722 70306 10734
rect 70254 10658 70306 10670
rect 70702 10722 70754 10734
rect 70702 10658 70754 10670
rect 71374 10722 71426 10734
rect 71374 10658 71426 10670
rect 72270 10722 72322 10734
rect 72270 10658 72322 10670
rect 77870 10722 77922 10734
rect 77870 10658 77922 10670
rect 31166 10610 31218 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 30818 10558 30830 10610
rect 30882 10558 30894 10610
rect 31166 10546 31218 10558
rect 31390 10610 31442 10622
rect 33070 10610 33122 10622
rect 31938 10558 31950 10610
rect 32002 10558 32014 10610
rect 31390 10546 31442 10558
rect 33070 10546 33122 10558
rect 40126 10610 40178 10622
rect 40126 10546 40178 10558
rect 40350 10610 40402 10622
rect 72830 10610 72882 10622
rect 40898 10558 40910 10610
rect 40962 10558 40974 10610
rect 46722 10558 46734 10610
rect 46786 10558 46798 10610
rect 46946 10558 46958 10610
rect 47010 10558 47022 10610
rect 49186 10558 49198 10610
rect 49250 10558 49262 10610
rect 70914 10558 70926 10610
rect 70978 10558 70990 10610
rect 40350 10546 40402 10558
rect 72830 10546 72882 10558
rect 78206 10610 78258 10622
rect 78206 10546 78258 10558
rect 12910 10498 12962 10510
rect 10322 10446 10334 10498
rect 10386 10446 10398 10498
rect 12450 10446 12462 10498
rect 12514 10446 12526 10498
rect 12910 10434 12962 10446
rect 13358 10498 13410 10510
rect 13358 10434 13410 10446
rect 14030 10498 14082 10510
rect 14030 10434 14082 10446
rect 15038 10498 15090 10510
rect 15038 10434 15090 10446
rect 16382 10498 16434 10510
rect 16382 10434 16434 10446
rect 17502 10498 17554 10510
rect 17502 10434 17554 10446
rect 18510 10498 18562 10510
rect 18510 10434 18562 10446
rect 26798 10498 26850 10510
rect 26798 10434 26850 10446
rect 27246 10498 27298 10510
rect 27246 10434 27298 10446
rect 27694 10498 27746 10510
rect 34414 10498 34466 10510
rect 36654 10498 36706 10510
rect 28018 10446 28030 10498
rect 28082 10446 28094 10498
rect 34738 10446 34750 10498
rect 34802 10446 34814 10498
rect 27694 10434 27746 10446
rect 34414 10434 34466 10446
rect 36654 10434 36706 10446
rect 37214 10498 37266 10510
rect 40238 10498 40290 10510
rect 46510 10498 46562 10510
rect 37538 10446 37550 10498
rect 37602 10446 37614 10498
rect 43698 10446 43710 10498
rect 43762 10446 43774 10498
rect 37214 10434 37266 10446
rect 40238 10434 40290 10446
rect 46510 10434 46562 10446
rect 48750 10498 48802 10510
rect 52558 10498 52610 10510
rect 49746 10446 49758 10498
rect 49810 10446 49822 10498
rect 48750 10434 48802 10446
rect 52558 10434 52610 10446
rect 53006 10498 53058 10510
rect 53006 10434 53058 10446
rect 53566 10498 53618 10510
rect 53566 10434 53618 10446
rect 54014 10498 54066 10510
rect 54014 10434 54066 10446
rect 63534 10498 63586 10510
rect 63534 10434 63586 10446
rect 63982 10498 64034 10510
rect 63982 10434 64034 10446
rect 64542 10498 64594 10510
rect 64542 10434 64594 10446
rect 65102 10498 65154 10510
rect 65102 10434 65154 10446
rect 65438 10498 65490 10510
rect 65438 10434 65490 10446
rect 66222 10498 66274 10510
rect 66222 10434 66274 10446
rect 67006 10498 67058 10510
rect 67006 10434 67058 10446
rect 67678 10498 67730 10510
rect 67678 10434 67730 10446
rect 68126 10498 68178 10510
rect 68126 10434 68178 10446
rect 68798 10498 68850 10510
rect 68798 10434 68850 10446
rect 69134 10498 69186 10510
rect 69134 10434 69186 10446
rect 69806 10498 69858 10510
rect 69806 10434 69858 10446
rect 73278 10498 73330 10510
rect 73278 10434 73330 10446
rect 73838 10498 73890 10510
rect 73838 10434 73890 10446
rect 74174 10498 74226 10510
rect 74174 10434 74226 10446
rect 74622 10498 74674 10510
rect 74622 10434 74674 10446
rect 75182 10498 75234 10510
rect 75182 10434 75234 10446
rect 75966 10498 76018 10510
rect 75966 10434 76018 10446
rect 76638 10498 76690 10510
rect 76638 10434 76690 10446
rect 77646 10498 77698 10510
rect 77646 10434 77698 10446
rect 39454 10386 39506 10398
rect 32274 10334 32286 10386
rect 32338 10334 32350 10386
rect 52658 10334 52670 10386
rect 52722 10383 52734 10386
rect 53554 10383 53566 10386
rect 52722 10337 53566 10383
rect 52722 10334 52734 10337
rect 53554 10334 53566 10337
rect 53618 10334 53630 10386
rect 74162 10334 74174 10386
rect 74226 10383 74238 10386
rect 74722 10383 74734 10386
rect 74226 10337 74734 10383
rect 74226 10334 74238 10337
rect 74722 10334 74734 10337
rect 74786 10334 74798 10386
rect 39454 10322 39506 10334
rect 1344 10218 78624 10252
rect 1344 10166 10874 10218
rect 10926 10166 10978 10218
rect 11030 10166 11082 10218
rect 11134 10166 30194 10218
rect 30246 10166 30298 10218
rect 30350 10166 30402 10218
rect 30454 10166 49514 10218
rect 49566 10166 49618 10218
rect 49670 10166 49722 10218
rect 49774 10166 68834 10218
rect 68886 10166 68938 10218
rect 68990 10166 69042 10218
rect 69094 10166 78624 10218
rect 1344 10132 78624 10166
rect 70142 10050 70194 10062
rect 36418 9998 36430 10050
rect 36482 9998 36494 10050
rect 70142 9986 70194 9998
rect 70478 10050 70530 10062
rect 70478 9986 70530 9998
rect 9438 9938 9490 9950
rect 18734 9938 18786 9950
rect 18274 9886 18286 9938
rect 18338 9886 18350 9938
rect 9438 9874 9490 9886
rect 18734 9874 18786 9886
rect 20302 9938 20354 9950
rect 28702 9938 28754 9950
rect 32062 9938 32114 9950
rect 35870 9938 35922 9950
rect 37998 9938 38050 9950
rect 40798 9938 40850 9950
rect 22082 9886 22094 9938
rect 22146 9886 22158 9938
rect 24210 9886 24222 9938
rect 24274 9886 24286 9938
rect 27570 9886 27582 9938
rect 27634 9886 27646 9938
rect 29922 9886 29934 9938
rect 29986 9886 29998 9938
rect 32610 9886 32622 9938
rect 32674 9886 32686 9938
rect 34738 9886 34750 9938
rect 34802 9886 34814 9938
rect 37426 9886 37438 9938
rect 37490 9886 37502 9938
rect 38882 9886 38894 9938
rect 38946 9886 38958 9938
rect 20302 9874 20354 9886
rect 28702 9874 28754 9886
rect 32062 9874 32114 9886
rect 35870 9874 35922 9886
rect 37998 9874 38050 9886
rect 40798 9874 40850 9886
rect 41470 9938 41522 9950
rect 41470 9874 41522 9886
rect 45166 9938 45218 9950
rect 54574 9938 54626 9950
rect 45826 9886 45838 9938
rect 45890 9886 45902 9938
rect 47058 9886 47070 9938
rect 47122 9886 47134 9938
rect 49298 9886 49310 9938
rect 49362 9886 49374 9938
rect 45166 9874 45218 9886
rect 54574 9874 54626 9886
rect 11566 9826 11618 9838
rect 28142 9826 28194 9838
rect 36094 9826 36146 9838
rect 12114 9774 12126 9826
rect 12178 9774 12190 9826
rect 15362 9774 15374 9826
rect 15426 9774 15438 9826
rect 21410 9774 21422 9826
rect 21474 9774 21486 9826
rect 29250 9774 29262 9826
rect 29314 9774 29326 9826
rect 35522 9774 35534 9826
rect 35586 9774 35598 9826
rect 11566 9762 11618 9774
rect 28142 9762 28194 9774
rect 36094 9762 36146 9774
rect 36990 9826 37042 9838
rect 63086 9826 63138 9838
rect 45714 9774 45726 9826
rect 45778 9774 45790 9826
rect 49970 9774 49982 9826
rect 50034 9774 50046 9826
rect 71250 9774 71262 9826
rect 71314 9774 71326 9826
rect 72594 9774 72606 9826
rect 72658 9774 72670 9826
rect 78082 9774 78094 9826
rect 78146 9774 78158 9826
rect 36990 9762 37042 9774
rect 63086 9762 63138 9774
rect 10222 9714 10274 9726
rect 10222 9650 10274 9662
rect 10558 9714 10610 9726
rect 10558 9650 10610 9662
rect 11230 9714 11282 9726
rect 14366 9714 14418 9726
rect 12338 9662 12350 9714
rect 12402 9662 12414 9714
rect 11230 9650 11282 9662
rect 14366 9650 14418 9662
rect 14702 9714 14754 9726
rect 46622 9714 46674 9726
rect 16146 9662 16158 9714
rect 16210 9662 16222 9714
rect 26450 9662 26462 9714
rect 26514 9662 26526 9714
rect 39890 9662 39902 9714
rect 39954 9662 39966 9714
rect 42018 9662 42030 9714
rect 42082 9662 42094 9714
rect 14702 9650 14754 9662
rect 46622 9650 46674 9662
rect 50766 9714 50818 9726
rect 50766 9650 50818 9662
rect 65662 9714 65714 9726
rect 65662 9650 65714 9662
rect 66782 9714 66834 9726
rect 66782 9650 66834 9662
rect 67454 9714 67506 9726
rect 67454 9650 67506 9662
rect 67790 9714 67842 9726
rect 72046 9714 72098 9726
rect 74062 9714 74114 9726
rect 71026 9662 71038 9714
rect 71090 9662 71102 9714
rect 73042 9662 73054 9714
rect 73106 9662 73118 9714
rect 67790 9650 67842 9662
rect 72046 9650 72098 9662
rect 74062 9650 74114 9662
rect 76862 9714 76914 9726
rect 76862 9650 76914 9662
rect 77198 9714 77250 9726
rect 77198 9650 77250 9662
rect 77870 9714 77922 9726
rect 77870 9650 77922 9662
rect 9998 9602 10050 9614
rect 9998 9538 10050 9550
rect 12910 9602 12962 9614
rect 12910 9538 12962 9550
rect 13582 9602 13634 9614
rect 13582 9538 13634 9550
rect 14142 9602 14194 9614
rect 14142 9538 14194 9550
rect 19182 9602 19234 9614
rect 19182 9538 19234 9550
rect 19854 9602 19906 9614
rect 19854 9538 19906 9550
rect 20862 9602 20914 9614
rect 20862 9538 20914 9550
rect 24894 9602 24946 9614
rect 24894 9538 24946 9550
rect 25342 9602 25394 9614
rect 25342 9538 25394 9550
rect 25790 9602 25842 9614
rect 25790 9538 25842 9550
rect 38670 9602 38722 9614
rect 38670 9538 38722 9550
rect 44382 9602 44434 9614
rect 44382 9538 44434 9550
rect 50542 9602 50594 9614
rect 50542 9538 50594 9550
rect 50654 9602 50706 9614
rect 50654 9538 50706 9550
rect 51102 9602 51154 9614
rect 51102 9538 51154 9550
rect 51550 9602 51602 9614
rect 51550 9538 51602 9550
rect 51998 9602 52050 9614
rect 51998 9538 52050 9550
rect 52670 9602 52722 9614
rect 52670 9538 52722 9550
rect 53118 9602 53170 9614
rect 53118 9538 53170 9550
rect 53566 9602 53618 9614
rect 53566 9538 53618 9550
rect 54014 9602 54066 9614
rect 54014 9538 54066 9550
rect 55022 9602 55074 9614
rect 55022 9538 55074 9550
rect 59950 9602 60002 9614
rect 59950 9538 60002 9550
rect 60846 9602 60898 9614
rect 60846 9538 60898 9550
rect 61294 9602 61346 9614
rect 61294 9538 61346 9550
rect 62526 9602 62578 9614
rect 62526 9538 62578 9550
rect 63422 9602 63474 9614
rect 63422 9538 63474 9550
rect 64206 9602 64258 9614
rect 64206 9538 64258 9550
rect 64766 9602 64818 9614
rect 64766 9538 64818 9550
rect 65326 9602 65378 9614
rect 65326 9538 65378 9550
rect 66222 9602 66274 9614
rect 66222 9538 66274 9550
rect 67006 9602 67058 9614
rect 67006 9538 67058 9550
rect 68574 9602 68626 9614
rect 68574 9538 68626 9550
rect 69022 9602 69074 9614
rect 69022 9538 69074 9550
rect 69470 9602 69522 9614
rect 69470 9538 69522 9550
rect 71710 9602 71762 9614
rect 71710 9538 71762 9550
rect 72382 9602 72434 9614
rect 72382 9538 72434 9550
rect 73390 9602 73442 9614
rect 73390 9538 73442 9550
rect 73726 9602 73778 9614
rect 73726 9538 73778 9550
rect 74398 9602 74450 9614
rect 74398 9538 74450 9550
rect 74958 9602 75010 9614
rect 74958 9538 75010 9550
rect 75406 9602 75458 9614
rect 75406 9538 75458 9550
rect 76190 9602 76242 9614
rect 76190 9538 76242 9550
rect 1344 9434 78784 9468
rect 1344 9382 20534 9434
rect 20586 9382 20638 9434
rect 20690 9382 20742 9434
rect 20794 9382 39854 9434
rect 39906 9382 39958 9434
rect 40010 9382 40062 9434
rect 40114 9382 59174 9434
rect 59226 9382 59278 9434
rect 59330 9382 59382 9434
rect 59434 9382 78494 9434
rect 78546 9382 78598 9434
rect 78650 9382 78702 9434
rect 78754 9382 78784 9434
rect 1344 9348 78784 9382
rect 17502 9266 17554 9278
rect 17502 9202 17554 9214
rect 18846 9266 18898 9278
rect 18846 9202 18898 9214
rect 22542 9266 22594 9278
rect 22542 9202 22594 9214
rect 26462 9266 26514 9278
rect 34190 9266 34242 9278
rect 30930 9214 30942 9266
rect 30994 9214 31006 9266
rect 26462 9202 26514 9214
rect 34190 9202 34242 9214
rect 34638 9266 34690 9278
rect 34638 9202 34690 9214
rect 41694 9266 41746 9278
rect 41694 9202 41746 9214
rect 47854 9266 47906 9278
rect 47854 9202 47906 9214
rect 58942 9266 58994 9278
rect 58942 9202 58994 9214
rect 59390 9266 59442 9278
rect 59390 9202 59442 9214
rect 60174 9266 60226 9278
rect 60174 9202 60226 9214
rect 61182 9266 61234 9278
rect 61182 9202 61234 9214
rect 63534 9266 63586 9278
rect 63534 9202 63586 9214
rect 64654 9266 64706 9278
rect 64654 9202 64706 9214
rect 65326 9266 65378 9278
rect 65326 9202 65378 9214
rect 66782 9266 66834 9278
rect 66782 9202 66834 9214
rect 69246 9266 69298 9278
rect 69246 9202 69298 9214
rect 75854 9266 75906 9278
rect 75854 9202 75906 9214
rect 9998 9154 10050 9166
rect 9998 9090 10050 9102
rect 10334 9154 10386 9166
rect 13582 9154 13634 9166
rect 12002 9102 12014 9154
rect 12066 9102 12078 9154
rect 10334 9090 10386 9102
rect 13582 9090 13634 9102
rect 17726 9154 17778 9166
rect 24110 9154 24162 9166
rect 23426 9102 23438 9154
rect 23490 9102 23502 9154
rect 17726 9090 17778 9102
rect 24110 9090 24162 9102
rect 24558 9154 24610 9166
rect 24558 9090 24610 9102
rect 25678 9154 25730 9166
rect 25678 9090 25730 9102
rect 26350 9154 26402 9166
rect 33406 9154 33458 9166
rect 41358 9154 41410 9166
rect 47742 9154 47794 9166
rect 30482 9102 30494 9154
rect 30546 9102 30558 9154
rect 31378 9102 31390 9154
rect 31442 9102 31454 9154
rect 35970 9102 35982 9154
rect 36034 9102 36046 9154
rect 37202 9102 37214 9154
rect 37266 9102 37278 9154
rect 40226 9102 40238 9154
rect 40290 9102 40302 9154
rect 47170 9102 47182 9154
rect 47234 9102 47246 9154
rect 26350 9090 26402 9102
rect 33406 9090 33458 9102
rect 41358 9090 41410 9102
rect 47742 9090 47794 9102
rect 48862 9154 48914 9166
rect 48862 9090 48914 9102
rect 49422 9154 49474 9166
rect 61966 9154 62018 9166
rect 55458 9102 55470 9154
rect 55522 9102 55534 9154
rect 49422 9090 49474 9102
rect 61966 9090 62018 9102
rect 62862 9154 62914 9166
rect 67454 9154 67506 9166
rect 65986 9102 65998 9154
rect 66050 9102 66062 9154
rect 62862 9090 62914 9102
rect 67454 9090 67506 9102
rect 67902 9154 67954 9166
rect 67902 9090 67954 9102
rect 68574 9154 68626 9166
rect 76862 9154 76914 9166
rect 69794 9102 69806 9154
rect 69858 9102 69870 9154
rect 71250 9102 71262 9154
rect 71314 9102 71326 9154
rect 73266 9102 73278 9154
rect 73330 9102 73342 9154
rect 74162 9102 74174 9154
rect 74226 9102 74238 9154
rect 68574 9090 68626 9102
rect 10670 9042 10722 9054
rect 9762 8990 9774 9042
rect 9826 8990 9838 9042
rect 10670 8978 10722 8990
rect 11118 9042 11170 9054
rect 11118 8978 11170 8990
rect 11454 9042 11506 9054
rect 17390 9042 17442 9054
rect 12114 8990 12126 9042
rect 12178 8990 12190 9042
rect 13346 8990 13358 9042
rect 13410 8990 13422 9042
rect 16818 8990 16830 9042
rect 16882 8990 16894 9042
rect 11454 8978 11506 8990
rect 17390 8978 17442 8990
rect 17838 9042 17890 9054
rect 33070 9042 33122 9054
rect 21858 8990 21870 9042
rect 21922 8990 21934 9042
rect 23650 8990 23662 9042
rect 23714 8990 23726 9042
rect 27010 8990 27022 9042
rect 27074 8990 27086 9042
rect 30706 8990 30718 9042
rect 30770 8990 30782 9042
rect 31490 8990 31502 9042
rect 31554 8990 31566 9042
rect 32498 8990 32510 9042
rect 32562 8990 32574 9042
rect 17838 8978 17890 8990
rect 33070 8978 33122 8990
rect 33518 9042 33570 9054
rect 40910 9042 40962 9054
rect 37090 8990 37102 9042
rect 37154 8990 37166 9042
rect 33518 8978 33570 8990
rect 40910 8978 40962 8990
rect 41022 9042 41074 9054
rect 41806 9042 41858 9054
rect 53902 9042 53954 9054
rect 41570 8990 41582 9042
rect 41634 8990 41646 9042
rect 45378 8990 45390 9042
rect 45442 8990 45454 9042
rect 52994 8990 53006 9042
rect 53058 8990 53070 9042
rect 41022 8978 41074 8990
rect 41806 8978 41858 8990
rect 53902 8978 53954 8990
rect 62526 9042 62578 9054
rect 62526 8978 62578 8990
rect 63198 9042 63250 9054
rect 63198 8978 63250 8990
rect 63870 9042 63922 9054
rect 65662 9042 65714 9054
rect 67118 9042 67170 9054
rect 64866 8990 64878 9042
rect 64930 8990 64942 9042
rect 66210 8990 66222 9042
rect 66274 8990 66286 9042
rect 63870 8978 63922 8990
rect 65662 8978 65714 8990
rect 67118 8978 67170 8990
rect 68238 9042 68290 9054
rect 69582 9042 69634 9054
rect 68786 8990 68798 9042
rect 68850 8990 68862 9042
rect 68238 8978 68290 8990
rect 69582 8978 69634 8990
rect 8542 8930 8594 8942
rect 8542 8866 8594 8878
rect 9102 8930 9154 8942
rect 9102 8866 9154 8878
rect 13022 8930 13074 8942
rect 33182 8930 33234 8942
rect 37998 8930 38050 8942
rect 13906 8878 13918 8930
rect 13970 8878 13982 8930
rect 16034 8878 16046 8930
rect 16098 8878 16110 8930
rect 19058 8878 19070 8930
rect 19122 8878 19134 8930
rect 21186 8878 21198 8930
rect 21250 8878 21262 8930
rect 27682 8878 27694 8930
rect 27746 8878 27758 8930
rect 29810 8878 29822 8930
rect 29874 8878 29886 8930
rect 34962 8878 34974 8930
rect 35026 8878 35038 8930
rect 37538 8878 37550 8930
rect 37602 8878 37614 8930
rect 13022 8866 13074 8878
rect 33182 8866 33234 8878
rect 37998 8866 38050 8878
rect 38558 8930 38610 8942
rect 42590 8930 42642 8942
rect 49086 8930 49138 8942
rect 39106 8878 39118 8930
rect 39170 8878 39182 8930
rect 44706 8878 44718 8930
rect 44770 8878 44782 8930
rect 45826 8878 45838 8930
rect 45890 8878 45902 8930
rect 48850 8878 48862 8930
rect 48914 8878 48926 8930
rect 38558 8866 38610 8878
rect 42590 8866 42642 8878
rect 49086 8866 49138 8878
rect 50094 8930 50146 8942
rect 53454 8930 53506 8942
rect 56814 8930 56866 8942
rect 52210 8878 52222 8930
rect 52274 8878 52286 8930
rect 54338 8878 54350 8930
rect 54402 8878 54414 8930
rect 50094 8866 50146 8878
rect 53454 8866 53506 8878
rect 56814 8866 56866 8878
rect 57150 8930 57202 8942
rect 57150 8866 57202 8878
rect 60846 8930 60898 8942
rect 60846 8866 60898 8878
rect 61742 8930 61794 8942
rect 61742 8866 61794 8878
rect 22878 8818 22930 8830
rect 22878 8754 22930 8766
rect 25566 8818 25618 8830
rect 25566 8754 25618 8766
rect 25902 8818 25954 8830
rect 25902 8754 25954 8766
rect 26574 8818 26626 8830
rect 26574 8754 26626 8766
rect 47966 8818 48018 8830
rect 69809 8818 69855 9102
rect 76862 9090 76914 9102
rect 77534 9154 77586 9166
rect 77534 9090 77586 9102
rect 70478 9042 70530 9054
rect 76190 9042 76242 9054
rect 71138 8990 71150 9042
rect 71202 8990 71214 9042
rect 77074 8990 77086 9042
rect 77138 8990 77150 9042
rect 77746 8990 77758 9042
rect 77810 8990 77822 9042
rect 70478 8978 70530 8990
rect 76190 8978 76242 8990
rect 72258 8878 72270 8930
rect 72322 8878 72334 8930
rect 75506 8878 75518 8930
rect 75570 8878 75582 8930
rect 70142 8818 70194 8830
rect 53218 8766 53230 8818
rect 53282 8815 53294 8818
rect 53442 8815 53454 8818
rect 53282 8769 53454 8815
rect 53282 8766 53294 8769
rect 53442 8766 53454 8769
rect 53506 8766 53518 8818
rect 60498 8766 60510 8818
rect 60562 8815 60574 8818
rect 61618 8815 61630 8818
rect 60562 8769 61630 8815
rect 60562 8766 60574 8769
rect 61618 8766 61630 8769
rect 61682 8766 61694 8818
rect 69794 8766 69806 8818
rect 69858 8766 69870 8818
rect 47966 8754 48018 8766
rect 70142 8754 70194 8766
rect 1344 8650 78624 8684
rect 1344 8598 10874 8650
rect 10926 8598 10978 8650
rect 11030 8598 11082 8650
rect 11134 8598 30194 8650
rect 30246 8598 30298 8650
rect 30350 8598 30402 8650
rect 30454 8598 49514 8650
rect 49566 8598 49618 8650
rect 49670 8598 49722 8650
rect 49774 8598 68834 8650
rect 68886 8598 68938 8650
rect 68990 8598 69042 8650
rect 69094 8598 78624 8650
rect 1344 8564 78624 8598
rect 17838 8482 17890 8494
rect 17838 8418 17890 8430
rect 43710 8482 43762 8494
rect 43710 8418 43762 8430
rect 14030 8370 14082 8382
rect 12002 8318 12014 8370
rect 12066 8318 12078 8370
rect 14030 8306 14082 8318
rect 19406 8370 19458 8382
rect 19406 8306 19458 8318
rect 20302 8370 20354 8382
rect 36430 8370 36482 8382
rect 23874 8318 23886 8370
rect 23938 8318 23950 8370
rect 25106 8318 25118 8370
rect 25170 8318 25182 8370
rect 27234 8318 27246 8370
rect 27298 8318 27310 8370
rect 35522 8318 35534 8370
rect 35586 8318 35598 8370
rect 20302 8306 20354 8318
rect 36430 8306 36482 8318
rect 37438 8370 37490 8382
rect 47966 8370 48018 8382
rect 42018 8318 42030 8370
rect 42082 8318 42094 8370
rect 45042 8318 45054 8370
rect 45106 8318 45118 8370
rect 48626 8318 48638 8370
rect 48690 8318 48702 8370
rect 50754 8318 50766 8370
rect 50818 8318 50830 8370
rect 51538 8318 51550 8370
rect 51602 8318 51614 8370
rect 52994 8318 53006 8370
rect 53058 8318 53070 8370
rect 53778 8318 53790 8370
rect 53842 8318 53854 8370
rect 58370 8318 58382 8370
rect 58434 8318 58446 8370
rect 62178 8318 62190 8370
rect 62242 8318 62254 8370
rect 68338 8318 68350 8370
rect 68402 8318 68414 8370
rect 70130 8318 70142 8370
rect 70194 8318 70206 8370
rect 73154 8318 73166 8370
rect 73218 8318 73230 8370
rect 73714 8318 73726 8370
rect 73778 8318 73790 8370
rect 76178 8318 76190 8370
rect 76242 8318 76254 8370
rect 37438 8306 37490 8318
rect 47966 8306 48018 8318
rect 15822 8258 15874 8270
rect 9090 8206 9102 8258
rect 9154 8206 9166 8258
rect 9874 8206 9886 8258
rect 9938 8206 9950 8258
rect 12450 8206 12462 8258
rect 12514 8206 12526 8258
rect 15138 8206 15150 8258
rect 15202 8206 15214 8258
rect 15822 8194 15874 8206
rect 16382 8258 16434 8270
rect 16382 8194 16434 8206
rect 16942 8258 16994 8270
rect 16942 8194 16994 8206
rect 17502 8258 17554 8270
rect 19854 8258 19906 8270
rect 17826 8206 17838 8258
rect 17890 8206 17902 8258
rect 19170 8206 19182 8258
rect 19234 8206 19246 8258
rect 17502 8194 17554 8206
rect 19854 8194 19906 8206
rect 20190 8258 20242 8270
rect 20190 8194 20242 8206
rect 20526 8258 20578 8270
rect 20526 8194 20578 8206
rect 21646 8258 21698 8270
rect 27918 8258 27970 8270
rect 35870 8258 35922 8270
rect 39902 8258 39954 8270
rect 44382 8258 44434 8270
rect 23538 8206 23550 8258
rect 23602 8206 23614 8258
rect 24322 8206 24334 8258
rect 24386 8206 24398 8258
rect 34402 8206 34414 8258
rect 34466 8206 34478 8258
rect 37762 8206 37774 8258
rect 37826 8206 37838 8258
rect 44034 8206 44046 8258
rect 44098 8206 44110 8258
rect 50430 8258 50482 8270
rect 62526 8258 62578 8270
rect 21646 8194 21698 8206
rect 27918 8194 27970 8206
rect 35870 8194 35922 8206
rect 39902 8194 39954 8206
rect 44382 8194 44434 8206
rect 44830 8202 44882 8214
rect 8094 8146 8146 8158
rect 8094 8082 8146 8094
rect 13806 8146 13858 8158
rect 13806 8082 13858 8094
rect 15374 8146 15426 8158
rect 15374 8082 15426 8094
rect 15934 8146 15986 8158
rect 15934 8082 15986 8094
rect 16606 8146 16658 8158
rect 16606 8082 16658 8094
rect 17166 8146 17218 8158
rect 17166 8082 17218 8094
rect 18510 8146 18562 8158
rect 18510 8082 18562 8094
rect 19518 8146 19570 8158
rect 28030 8146 28082 8158
rect 21298 8094 21310 8146
rect 21362 8094 21374 8146
rect 19518 8082 19570 8094
rect 22542 8090 22594 8102
rect 6302 8034 6354 8046
rect 6302 7970 6354 7982
rect 7422 8034 7474 8046
rect 7422 7970 7474 7982
rect 7870 8034 7922 8046
rect 7870 7970 7922 7982
rect 8430 8034 8482 8046
rect 8430 7970 8482 7982
rect 12686 8034 12738 8046
rect 12686 7970 12738 7982
rect 14590 8034 14642 8046
rect 14590 7970 14642 7982
rect 16046 8034 16098 8046
rect 16046 7970 16098 7982
rect 16718 8034 16770 8046
rect 16718 7970 16770 7982
rect 18174 8034 18226 8046
rect 18174 7970 18226 7982
rect 22094 8034 22146 8046
rect 28030 8082 28082 8094
rect 28142 8146 28194 8158
rect 34862 8146 34914 8158
rect 30258 8094 30270 8146
rect 30322 8094 30334 8146
rect 28142 8082 28194 8094
rect 34862 8082 34914 8094
rect 34974 8146 35026 8158
rect 34974 8082 35026 8094
rect 35086 8146 35138 8158
rect 35086 8082 35138 8094
rect 37214 8146 37266 8158
rect 37214 8082 37266 8094
rect 37326 8146 37378 8158
rect 37326 8082 37378 8094
rect 38894 8146 38946 8158
rect 38894 8082 38946 8094
rect 40350 8146 40402 8158
rect 51874 8206 51886 8258
rect 51938 8206 51950 8258
rect 58482 8206 58494 8258
rect 58546 8206 58558 8258
rect 61730 8206 61742 8258
rect 61794 8206 61806 8258
rect 50430 8194 50482 8206
rect 62526 8194 62578 8206
rect 63534 8258 63586 8270
rect 63534 8194 63586 8206
rect 63646 8258 63698 8270
rect 64430 8258 64482 8270
rect 63858 8206 63870 8258
rect 63922 8206 63934 8258
rect 63646 8194 63698 8206
rect 64430 8194 64482 8206
rect 64990 8258 65042 8270
rect 65538 8206 65550 8258
rect 65602 8206 65614 8258
rect 66882 8206 66894 8258
rect 66946 8206 66958 8258
rect 67554 8206 67566 8258
rect 67618 8206 67630 8258
rect 64990 8194 65042 8206
rect 43362 8094 43374 8146
rect 43426 8094 43438 8146
rect 44830 8138 44882 8150
rect 45278 8146 45330 8158
rect 52670 8146 52722 8158
rect 45826 8094 45838 8146
rect 45890 8094 45902 8146
rect 49634 8094 49646 8146
rect 49698 8094 49710 8146
rect 51986 8094 51998 8146
rect 52050 8094 52062 8146
rect 40350 8082 40402 8094
rect 45278 8082 45330 8094
rect 52670 8082 52722 8094
rect 52894 8146 52946 8158
rect 57934 8146 57986 8158
rect 55010 8094 55022 8146
rect 55074 8094 55086 8146
rect 52894 8082 52946 8094
rect 57934 8082 57986 8094
rect 61070 8146 61122 8158
rect 61070 8082 61122 8094
rect 65998 8146 66050 8158
rect 65998 8082 66050 8094
rect 66334 8146 66386 8158
rect 66334 8082 66386 8094
rect 66670 8146 66722 8158
rect 69346 8094 69358 8146
rect 69410 8094 69422 8146
rect 71250 8094 71262 8146
rect 71314 8094 71326 8146
rect 72034 8094 72046 8146
rect 72098 8094 72110 8146
rect 74722 8094 74734 8146
rect 74786 8094 74798 8146
rect 77522 8094 77534 8146
rect 77586 8094 77598 8146
rect 66670 8082 66722 8094
rect 22542 8026 22594 8038
rect 22990 8034 23042 8046
rect 41022 8034 41074 8046
rect 22094 7970 22146 7982
rect 28578 7982 28590 8034
rect 28642 7982 28654 8034
rect 22990 7970 23042 7982
rect 41022 7970 41074 7982
rect 43822 8034 43874 8046
rect 43822 7970 43874 7982
rect 45054 8034 45106 8046
rect 45054 7970 45106 7982
rect 50654 8034 50706 8046
rect 50654 7970 50706 7982
rect 55470 8034 55522 8046
rect 55470 7970 55522 7982
rect 55918 8034 55970 8046
rect 55918 7970 55970 7982
rect 56366 8034 56418 8046
rect 56366 7970 56418 7982
rect 56814 8034 56866 8046
rect 56814 7970 56866 7982
rect 57262 8034 57314 8046
rect 57262 7970 57314 7982
rect 59054 8034 59106 8046
rect 59054 7970 59106 7982
rect 59502 8034 59554 8046
rect 59502 7970 59554 7982
rect 60622 8034 60674 8046
rect 62302 8034 62354 8046
rect 61506 7982 61518 8034
rect 61570 7982 61582 8034
rect 60622 7970 60674 7982
rect 62302 7970 62354 7982
rect 63310 8034 63362 8046
rect 63310 7970 63362 7982
rect 63422 8034 63474 8046
rect 67342 8034 67394 8046
rect 65314 7982 65326 8034
rect 65378 7982 65390 8034
rect 63422 7970 63474 7982
rect 67342 7970 67394 7982
rect 75518 8034 75570 8046
rect 75518 7970 75570 7982
rect 77982 8034 78034 8046
rect 77982 7970 78034 7982
rect 1344 7866 78784 7900
rect 1344 7814 20534 7866
rect 20586 7814 20638 7866
rect 20690 7814 20742 7866
rect 20794 7814 39854 7866
rect 39906 7814 39958 7866
rect 40010 7814 40062 7866
rect 40114 7814 59174 7866
rect 59226 7814 59278 7866
rect 59330 7814 59382 7866
rect 59434 7814 78494 7866
rect 78546 7814 78598 7866
rect 78650 7814 78702 7866
rect 78754 7814 78784 7866
rect 1344 7780 78784 7814
rect 7758 7698 7810 7710
rect 7758 7634 7810 7646
rect 9998 7698 10050 7710
rect 9998 7634 10050 7646
rect 10670 7698 10722 7710
rect 10670 7634 10722 7646
rect 17726 7698 17778 7710
rect 17726 7634 17778 7646
rect 24670 7698 24722 7710
rect 24670 7634 24722 7646
rect 26798 7698 26850 7710
rect 26798 7634 26850 7646
rect 29262 7698 29314 7710
rect 29262 7634 29314 7646
rect 29822 7698 29874 7710
rect 29822 7634 29874 7646
rect 30158 7698 30210 7710
rect 30158 7634 30210 7646
rect 30606 7698 30658 7710
rect 30606 7634 30658 7646
rect 38446 7698 38498 7710
rect 38446 7634 38498 7646
rect 38558 7698 38610 7710
rect 38558 7634 38610 7646
rect 38670 7698 38722 7710
rect 38670 7634 38722 7646
rect 41134 7698 41186 7710
rect 41134 7634 41186 7646
rect 41582 7698 41634 7710
rect 41582 7634 41634 7646
rect 43822 7698 43874 7710
rect 43822 7634 43874 7646
rect 44270 7698 44322 7710
rect 44270 7634 44322 7646
rect 47854 7698 47906 7710
rect 47854 7634 47906 7646
rect 48078 7698 48130 7710
rect 48078 7634 48130 7646
rect 48974 7698 49026 7710
rect 48974 7634 49026 7646
rect 53902 7698 53954 7710
rect 53902 7634 53954 7646
rect 54350 7698 54402 7710
rect 55470 7698 55522 7710
rect 54786 7646 54798 7698
rect 54850 7646 54862 7698
rect 54350 7634 54402 7646
rect 55470 7634 55522 7646
rect 56590 7698 56642 7710
rect 56590 7634 56642 7646
rect 58606 7698 58658 7710
rect 77086 7698 77138 7710
rect 66658 7646 66670 7698
rect 66722 7646 66734 7698
rect 58606 7634 58658 7646
rect 70814 7642 70866 7654
rect 6078 7586 6130 7598
rect 6078 7522 6130 7534
rect 7310 7586 7362 7598
rect 23662 7586 23714 7598
rect 8754 7534 8766 7586
rect 8818 7534 8830 7586
rect 7310 7522 7362 7534
rect 23662 7522 23714 7534
rect 25342 7586 25394 7598
rect 25342 7522 25394 7534
rect 25902 7586 25954 7598
rect 25902 7522 25954 7534
rect 26350 7586 26402 7598
rect 33518 7586 33570 7598
rect 47182 7586 47234 7598
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 31938 7534 31950 7586
rect 32002 7534 32014 7586
rect 35746 7534 35758 7586
rect 35810 7534 35822 7586
rect 36642 7534 36654 7586
rect 36706 7534 36718 7586
rect 42914 7534 42926 7586
rect 42978 7534 42990 7586
rect 45714 7534 45726 7586
rect 45778 7534 45790 7586
rect 26350 7522 26402 7534
rect 33518 7522 33570 7534
rect 47182 7522 47234 7534
rect 48750 7586 48802 7598
rect 53454 7586 53506 7598
rect 52322 7534 52334 7586
rect 52386 7534 52398 7586
rect 48750 7522 48802 7534
rect 53454 7522 53506 7534
rect 54462 7586 54514 7598
rect 57262 7586 57314 7598
rect 55794 7534 55806 7586
rect 55858 7534 55870 7586
rect 56914 7534 56926 7586
rect 56978 7534 56990 7586
rect 54462 7522 54514 7534
rect 57262 7522 57314 7534
rect 58382 7586 58434 7598
rect 58382 7522 58434 7534
rect 59278 7586 59330 7598
rect 59278 7522 59330 7534
rect 59726 7586 59778 7598
rect 59726 7522 59778 7534
rect 60174 7586 60226 7598
rect 60174 7522 60226 7534
rect 60958 7586 61010 7598
rect 65326 7586 65378 7598
rect 77086 7634 77138 7646
rect 62850 7534 62862 7586
rect 62914 7534 62926 7586
rect 65874 7534 65886 7586
rect 65938 7534 65950 7586
rect 67330 7534 67342 7586
rect 67394 7534 67406 7586
rect 70018 7534 70030 7586
rect 70082 7534 70094 7586
rect 70814 7578 70866 7590
rect 71486 7586 71538 7598
rect 77758 7586 77810 7598
rect 72370 7534 72382 7586
rect 72434 7534 72446 7586
rect 74386 7534 74398 7586
rect 74450 7534 74462 7586
rect 60958 7522 61010 7534
rect 65326 7522 65378 7534
rect 71486 7522 71538 7534
rect 77758 7522 77810 7534
rect 6974 7474 7026 7486
rect 5842 7422 5854 7474
rect 5906 7422 5918 7474
rect 6974 7410 7026 7422
rect 8094 7474 8146 7486
rect 9662 7474 9714 7486
rect 24110 7474 24162 7486
rect 34414 7474 34466 7486
rect 39454 7474 39506 7486
rect 46622 7474 46674 7486
rect 8866 7422 8878 7474
rect 8930 7422 8942 7474
rect 10434 7422 10446 7474
rect 10498 7422 10510 7474
rect 13122 7422 13134 7474
rect 13186 7422 13198 7474
rect 16482 7422 16494 7474
rect 16546 7422 16558 7474
rect 21746 7422 21758 7474
rect 21810 7422 21822 7474
rect 25666 7422 25678 7474
rect 25730 7422 25742 7474
rect 26562 7422 26574 7474
rect 26626 7422 26638 7474
rect 34066 7422 34078 7474
rect 34130 7422 34142 7474
rect 36194 7422 36206 7474
rect 36258 7422 36270 7474
rect 36418 7422 36430 7474
rect 36482 7422 36494 7474
rect 38994 7422 39006 7474
rect 39058 7422 39070 7474
rect 39890 7422 39902 7474
rect 39954 7422 39966 7474
rect 8094 7410 8146 7422
rect 9662 7410 9714 7422
rect 24110 7410 24162 7422
rect 34414 7410 34466 7422
rect 39454 7410 39506 7422
rect 46622 7410 46674 7422
rect 46734 7474 46786 7486
rect 46734 7410 46786 7422
rect 46846 7474 46898 7486
rect 46846 7410 46898 7422
rect 47518 7474 47570 7486
rect 47518 7410 47570 7422
rect 48190 7474 48242 7486
rect 48190 7410 48242 7422
rect 49086 7474 49138 7486
rect 49086 7410 49138 7422
rect 49310 7474 49362 7486
rect 55134 7474 55186 7486
rect 52994 7422 53006 7474
rect 53058 7422 53070 7474
rect 49310 7410 49362 7422
rect 55134 7410 55186 7422
rect 57486 7474 57538 7486
rect 71150 7474 71202 7486
rect 57698 7422 57710 7474
rect 57762 7422 57774 7474
rect 64530 7422 64542 7474
rect 64594 7422 64606 7474
rect 66322 7422 66334 7474
rect 66386 7422 66398 7474
rect 66882 7422 66894 7474
rect 66946 7422 66958 7474
rect 77298 7422 77310 7474
rect 77362 7422 77374 7474
rect 77970 7422 77982 7474
rect 78034 7422 78046 7474
rect 57486 7410 57538 7422
rect 71150 7410 71202 7422
rect 5518 7362 5570 7374
rect 5518 7298 5570 7310
rect 6526 7362 6578 7374
rect 33182 7362 33234 7374
rect 40350 7362 40402 7374
rect 47854 7362 47906 7374
rect 58494 7362 58546 7374
rect 18834 7310 18846 7362
rect 18898 7310 18910 7362
rect 26786 7310 26798 7362
rect 26850 7310 26862 7362
rect 28354 7310 28366 7362
rect 28418 7310 28430 7362
rect 30930 7310 30942 7362
rect 30994 7310 31006 7362
rect 38210 7310 38222 7362
rect 38274 7310 38286 7362
rect 41906 7310 41918 7362
rect 41970 7310 41982 7362
rect 44706 7310 44718 7362
rect 44770 7310 44782 7362
rect 50082 7310 50094 7362
rect 50146 7310 50158 7362
rect 6526 7298 6578 7310
rect 33182 7298 33234 7310
rect 40350 7298 40402 7310
rect 47854 7298 47906 7310
rect 58494 7298 58546 7310
rect 59166 7362 59218 7374
rect 63534 7362 63586 7374
rect 76526 7362 76578 7374
rect 61506 7310 61518 7362
rect 61570 7310 61582 7362
rect 64866 7310 64878 7362
rect 64930 7310 64942 7362
rect 68450 7310 68462 7362
rect 68514 7310 68526 7362
rect 69010 7310 69022 7362
rect 69074 7310 69086 7362
rect 73714 7310 73726 7362
rect 73778 7310 73790 7362
rect 59166 7298 59218 7310
rect 63534 7298 63586 7310
rect 76526 7298 76578 7310
rect 11230 7250 11282 7262
rect 11230 7186 11282 7198
rect 14142 7250 14194 7262
rect 14142 7186 14194 7198
rect 26014 7250 26066 7262
rect 26014 7186 26066 7198
rect 59054 7250 59106 7262
rect 59054 7186 59106 7198
rect 63422 7250 63474 7262
rect 63422 7186 63474 7198
rect 63758 7250 63810 7262
rect 63758 7186 63810 7198
rect 63870 7250 63922 7262
rect 63870 7186 63922 7198
rect 1344 7082 78624 7116
rect 1344 7030 10874 7082
rect 10926 7030 10978 7082
rect 11030 7030 11082 7082
rect 11134 7030 30194 7082
rect 30246 7030 30298 7082
rect 30350 7030 30402 7082
rect 30454 7030 49514 7082
rect 49566 7030 49618 7082
rect 49670 7030 49722 7082
rect 49774 7030 68834 7082
rect 68886 7030 68938 7082
rect 68990 7030 69042 7082
rect 69094 7030 78624 7082
rect 1344 6996 78624 7030
rect 14366 6914 14418 6926
rect 14366 6850 14418 6862
rect 20078 6914 20130 6926
rect 42030 6914 42082 6926
rect 55694 6914 55746 6926
rect 26450 6862 26462 6914
rect 26514 6911 26526 6914
rect 26514 6865 26623 6911
rect 26514 6862 26526 6865
rect 20078 6850 20130 6862
rect 9874 6750 9886 6802
rect 9938 6750 9950 6802
rect 16034 6750 16046 6802
rect 16098 6750 16110 6802
rect 20402 6750 20414 6802
rect 20466 6750 20478 6802
rect 6302 6690 6354 6702
rect 14702 6690 14754 6702
rect 15710 6690 15762 6702
rect 21198 6690 21250 6702
rect 5730 6638 5742 6690
rect 5794 6638 5806 6690
rect 7074 6638 7086 6690
rect 7138 6638 7150 6690
rect 7746 6638 7758 6690
rect 7810 6638 7822 6690
rect 12450 6638 12462 6690
rect 12514 6638 12526 6690
rect 13906 6638 13918 6690
rect 13970 6638 13982 6690
rect 15250 6638 15262 6690
rect 15314 6638 15326 6690
rect 18834 6638 18846 6690
rect 18898 6638 18910 6690
rect 19506 6638 19518 6690
rect 19570 6638 19582 6690
rect 6302 6626 6354 6638
rect 14702 6626 14754 6638
rect 15710 6626 15762 6638
rect 21198 6626 21250 6638
rect 21646 6690 21698 6702
rect 21646 6626 21698 6638
rect 21758 6690 21810 6702
rect 25118 6690 25170 6702
rect 23538 6638 23550 6690
rect 23602 6638 23614 6690
rect 24546 6638 24558 6690
rect 24610 6638 24622 6690
rect 25666 6638 25678 6690
rect 25730 6638 25742 6690
rect 21758 6626 21810 6638
rect 25118 6626 25170 6638
rect 4734 6578 4786 6590
rect 4734 6514 4786 6526
rect 5070 6578 5122 6590
rect 5070 6514 5122 6526
rect 6638 6578 6690 6590
rect 22990 6578 23042 6590
rect 11330 6526 11342 6578
rect 11394 6526 11406 6578
rect 13682 6526 13694 6578
rect 13746 6526 13758 6578
rect 18162 6526 18174 6578
rect 18226 6526 18238 6578
rect 19282 6526 19294 6578
rect 19346 6526 19358 6578
rect 24770 6526 24782 6578
rect 24834 6526 24846 6578
rect 25554 6526 25566 6578
rect 25618 6526 25630 6578
rect 6638 6514 6690 6526
rect 22990 6514 23042 6526
rect 4510 6466 4562 6478
rect 4510 6402 4562 6414
rect 5966 6466 6018 6478
rect 5966 6402 6018 6414
rect 20302 6466 20354 6478
rect 20302 6402 20354 6414
rect 21534 6466 21586 6478
rect 21534 6402 21586 6414
rect 22654 6466 22706 6478
rect 22654 6402 22706 6414
rect 23102 6466 23154 6478
rect 23102 6402 23154 6414
rect 23326 6466 23378 6478
rect 23326 6402 23378 6414
rect 26462 6466 26514 6478
rect 26577 6466 26623 6865
rect 40674 6862 40686 6914
rect 40738 6911 40750 6914
rect 41346 6911 41358 6914
rect 40738 6865 41358 6911
rect 40738 6862 40750 6865
rect 41346 6862 41358 6865
rect 41410 6862 41422 6914
rect 43138 6862 43150 6914
rect 43202 6862 43214 6914
rect 45154 6862 45166 6914
rect 45218 6911 45230 6914
rect 45490 6911 45502 6914
rect 45218 6865 45502 6911
rect 45218 6862 45230 6865
rect 45490 6862 45502 6865
rect 45554 6862 45566 6914
rect 50306 6911 50318 6914
rect 50097 6865 50318 6911
rect 42030 6850 42082 6862
rect 26910 6802 26962 6814
rect 34078 6802 34130 6814
rect 27122 6750 27134 6802
rect 27186 6750 27198 6802
rect 29362 6750 29374 6802
rect 29426 6750 29438 6802
rect 26910 6738 26962 6750
rect 34078 6738 34130 6750
rect 40014 6802 40066 6814
rect 40014 6738 40066 6750
rect 40910 6802 40962 6814
rect 45938 6750 45950 6802
rect 46002 6750 46014 6802
rect 49186 6750 49198 6802
rect 49250 6750 49262 6802
rect 40910 6738 40962 6750
rect 40238 6690 40290 6702
rect 29586 6638 29598 6690
rect 29650 6638 29662 6690
rect 31154 6638 31166 6690
rect 31218 6638 31230 6690
rect 36082 6638 36094 6690
rect 36146 6638 36158 6690
rect 36978 6638 36990 6690
rect 37042 6638 37054 6690
rect 37986 6638 37998 6690
rect 38050 6638 38062 6690
rect 39106 6638 39118 6690
rect 39170 6638 39182 6690
rect 39778 6638 39790 6690
rect 39842 6638 39854 6690
rect 40238 6626 40290 6638
rect 40350 6690 40402 6702
rect 40350 6626 40402 6638
rect 40462 6690 40514 6702
rect 42254 6690 42306 6702
rect 45614 6690 45666 6702
rect 50097 6690 50143 6865
rect 50306 6862 50318 6865
rect 50370 6862 50382 6914
rect 52546 6862 52558 6914
rect 52610 6911 52622 6914
rect 52770 6911 52782 6914
rect 52610 6865 52782 6911
rect 52610 6862 52622 6865
rect 52770 6862 52782 6865
rect 52834 6862 52846 6914
rect 55694 6850 55746 6862
rect 59614 6914 59666 6926
rect 59614 6850 59666 6862
rect 75630 6914 75682 6926
rect 75630 6850 75682 6862
rect 51774 6802 51826 6814
rect 50194 6750 50206 6802
rect 50258 6750 50270 6802
rect 41794 6638 41806 6690
rect 41858 6638 41870 6690
rect 42802 6638 42814 6690
rect 42866 6638 42878 6690
rect 43698 6638 43710 6690
rect 43762 6638 43774 6690
rect 44034 6638 44046 6690
rect 44098 6638 44110 6690
rect 50082 6638 50094 6690
rect 50146 6638 50158 6690
rect 40462 6626 40514 6638
rect 42254 6626 42306 6638
rect 45614 6626 45666 6638
rect 29150 6578 29202 6590
rect 39566 6578 39618 6590
rect 28130 6526 28142 6578
rect 28194 6526 28206 6578
rect 38210 6526 38222 6578
rect 38274 6526 38286 6578
rect 38882 6526 38894 6578
rect 38946 6526 38958 6578
rect 29150 6514 29202 6526
rect 39566 6514 39618 6526
rect 41582 6578 41634 6590
rect 41582 6514 41634 6526
rect 42478 6578 42530 6590
rect 42478 6514 42530 6526
rect 43038 6578 43090 6590
rect 50209 6578 50255 6750
rect 51774 6738 51826 6750
rect 52110 6802 52162 6814
rect 52110 6738 52162 6750
rect 52894 6802 52946 6814
rect 52894 6738 52946 6750
rect 58718 6802 58770 6814
rect 58718 6738 58770 6750
rect 60734 6802 60786 6814
rect 72830 6802 72882 6814
rect 61506 6750 61518 6802
rect 61570 6750 61582 6802
rect 63410 6750 63422 6802
rect 63474 6750 63486 6802
rect 65650 6750 65662 6802
rect 65714 6750 65726 6802
rect 69794 6750 69806 6802
rect 69858 6750 69870 6802
rect 77634 6750 77646 6802
rect 77698 6750 77710 6802
rect 60734 6738 60786 6750
rect 72830 6738 72882 6750
rect 51102 6690 51154 6702
rect 50754 6638 50766 6690
rect 50818 6638 50830 6690
rect 51102 6626 51154 6638
rect 51438 6690 51490 6702
rect 58930 6638 58942 6690
rect 58994 6638 59006 6690
rect 63298 6638 63310 6690
rect 63362 6638 63374 6690
rect 66546 6638 66558 6690
rect 66610 6638 66622 6690
rect 67666 6638 67678 6690
rect 67730 6638 67742 6690
rect 51438 6626 51490 6638
rect 58606 6578 58658 6590
rect 47058 6526 47070 6578
rect 47122 6526 47134 6578
rect 48066 6526 48078 6578
rect 48130 6526 48142 6578
rect 50194 6526 50206 6578
rect 50258 6526 50270 6578
rect 55346 6526 55358 6578
rect 55410 6526 55422 6578
rect 58146 6526 58158 6578
rect 58210 6526 58222 6578
rect 43038 6514 43090 6526
rect 58606 6514 58658 6526
rect 59502 6578 59554 6590
rect 63982 6578 64034 6590
rect 62850 6526 62862 6578
rect 62914 6526 62926 6578
rect 64530 6526 64542 6578
rect 64594 6526 64606 6578
rect 66658 6526 66670 6578
rect 66722 6526 66734 6578
rect 68562 6526 68574 6578
rect 68626 6526 68638 6578
rect 70354 6526 70366 6578
rect 70418 6526 70430 6578
rect 73490 6526 73502 6578
rect 73554 6526 73566 6578
rect 76290 6526 76302 6578
rect 76354 6526 76366 6578
rect 59502 6514 59554 6526
rect 63982 6514 64034 6526
rect 31950 6466 32002 6478
rect 42030 6466 42082 6478
rect 26562 6414 26574 6466
rect 26626 6414 26638 6466
rect 38098 6414 38110 6466
rect 38162 6414 38174 6466
rect 26462 6402 26514 6414
rect 31950 6402 32002 6414
rect 42030 6402 42082 6414
rect 44942 6466 44994 6478
rect 44942 6402 44994 6414
rect 49870 6466 49922 6478
rect 49870 6402 49922 6414
rect 50318 6466 50370 6478
rect 50318 6402 50370 6414
rect 50990 6466 51042 6478
rect 50990 6402 51042 6414
rect 51550 6466 51602 6478
rect 51550 6402 51602 6414
rect 59726 6466 59778 6478
rect 59726 6402 59778 6414
rect 59950 6466 60002 6478
rect 59950 6402 60002 6414
rect 61070 6466 61122 6478
rect 61070 6402 61122 6414
rect 63534 6466 63586 6478
rect 63534 6402 63586 6414
rect 63758 6466 63810 6478
rect 77982 6466 78034 6478
rect 67442 6414 67454 6466
rect 67506 6414 67518 6466
rect 63758 6402 63810 6414
rect 77982 6402 78034 6414
rect 1344 6298 78784 6332
rect 1344 6246 20534 6298
rect 20586 6246 20638 6298
rect 20690 6246 20742 6298
rect 20794 6246 39854 6298
rect 39906 6246 39958 6298
rect 40010 6246 40062 6298
rect 40114 6246 59174 6298
rect 59226 6246 59278 6298
rect 59330 6246 59382 6298
rect 59434 6246 78494 6298
rect 78546 6246 78598 6298
rect 78650 6246 78702 6298
rect 78754 6246 78784 6298
rect 1344 6212 78784 6246
rect 9662 6130 9714 6142
rect 9662 6066 9714 6078
rect 17614 6130 17666 6142
rect 17614 6066 17666 6078
rect 18510 6130 18562 6142
rect 18510 6066 18562 6078
rect 19518 6130 19570 6142
rect 40238 6130 40290 6142
rect 41694 6130 41746 6142
rect 24322 6078 24334 6130
rect 24386 6078 24398 6130
rect 33842 6078 33854 6130
rect 33906 6078 33918 6130
rect 40898 6078 40910 6130
rect 40962 6078 40974 6130
rect 19518 6066 19570 6078
rect 40238 6066 40290 6078
rect 41694 6066 41746 6078
rect 42926 6130 42978 6142
rect 42926 6066 42978 6078
rect 43934 6130 43986 6142
rect 43934 6066 43986 6078
rect 52334 6130 52386 6142
rect 52334 6066 52386 6078
rect 53902 6130 53954 6142
rect 53902 6066 53954 6078
rect 56702 6130 56754 6142
rect 56702 6066 56754 6078
rect 77646 6130 77698 6142
rect 77646 6066 77698 6078
rect 17726 6018 17778 6030
rect 10322 5966 10334 6018
rect 10386 5966 10398 6018
rect 10546 5966 10558 6018
rect 10610 5966 10622 6018
rect 17726 5954 17778 5966
rect 18174 6018 18226 6030
rect 23214 6018 23266 6030
rect 18834 5966 18846 6018
rect 18898 5966 18910 6018
rect 21970 5966 21982 6018
rect 22034 5966 22046 6018
rect 18174 5954 18226 5966
rect 23214 5954 23266 5966
rect 25342 6018 25394 6030
rect 25342 5954 25394 5966
rect 27470 6018 27522 6030
rect 27470 5954 27522 5966
rect 27806 6018 27858 6030
rect 33182 6018 33234 6030
rect 29362 5966 29374 6018
rect 29426 5966 29438 6018
rect 27806 5954 27858 5966
rect 33182 5954 33234 5966
rect 33294 6018 33346 6030
rect 33294 5954 33346 5966
rect 33406 6018 33458 6030
rect 33406 5954 33458 5966
rect 40014 6018 40066 6030
rect 40014 5954 40066 5966
rect 40350 6018 40402 6030
rect 40350 5954 40402 5966
rect 42254 6018 42306 6030
rect 44382 6018 44434 6030
rect 54238 6018 54290 6030
rect 55470 6018 55522 6030
rect 43138 5966 43150 6018
rect 43202 5966 43214 6018
rect 46498 5966 46510 6018
rect 46562 5966 46574 6018
rect 51314 5966 51326 6018
rect 51378 5966 51390 6018
rect 54562 5966 54574 6018
rect 54626 5966 54638 6018
rect 42254 5954 42306 5966
rect 44382 5954 44434 5966
rect 54238 5954 54290 5966
rect 55470 5954 55522 5966
rect 57262 6018 57314 6030
rect 57262 5954 57314 5966
rect 58046 6018 58098 6030
rect 64542 6018 64594 6030
rect 67790 6018 67842 6030
rect 71038 6018 71090 6030
rect 77870 6018 77922 6030
rect 58706 5966 58718 6018
rect 58770 5966 58782 6018
rect 61730 5966 61742 6018
rect 61794 5966 61806 6018
rect 62738 5966 62750 6018
rect 62802 5966 62814 6018
rect 65090 5966 65102 6018
rect 65154 5966 65166 6018
rect 68338 5966 68350 6018
rect 68402 5966 68414 6018
rect 72370 5966 72382 6018
rect 72434 5966 72446 6018
rect 75170 5966 75182 6018
rect 75234 5966 75246 6018
rect 58046 5954 58098 5966
rect 64542 5954 64594 5966
rect 67790 5954 67842 5966
rect 71038 5954 71090 5966
rect 77870 5954 77922 5966
rect 9998 5906 10050 5918
rect 23326 5906 23378 5918
rect 5954 5854 5966 5906
rect 6018 5854 6030 5906
rect 8978 5854 8990 5906
rect 9042 5854 9054 5906
rect 11778 5854 11790 5906
rect 11842 5854 11854 5906
rect 16370 5854 16382 5906
rect 16434 5854 16446 5906
rect 17378 5854 17390 5906
rect 17442 5854 17454 5906
rect 19282 5854 19294 5906
rect 19346 5854 19358 5906
rect 22754 5854 22766 5906
rect 22818 5854 22830 5906
rect 9998 5842 10050 5854
rect 23326 5842 23378 5854
rect 23438 5906 23490 5918
rect 23438 5842 23490 5854
rect 24670 5906 24722 5918
rect 24670 5842 24722 5854
rect 25678 5906 25730 5918
rect 25678 5842 25730 5854
rect 25902 5906 25954 5918
rect 41806 5906 41858 5918
rect 26562 5854 26574 5906
rect 26626 5854 26638 5906
rect 27682 5854 27694 5906
rect 27746 5854 27758 5906
rect 29922 5854 29934 5906
rect 29986 5854 29998 5906
rect 36866 5854 36878 5906
rect 36930 5854 36942 5906
rect 39330 5854 39342 5906
rect 39394 5854 39406 5906
rect 41122 5854 41134 5906
rect 41186 5854 41198 5906
rect 25902 5842 25954 5854
rect 15138 5742 15150 5794
rect 15202 5742 15214 5794
rect 19842 5742 19854 5794
rect 19906 5742 19918 5794
rect 5070 5682 5122 5694
rect 5070 5618 5122 5630
rect 7982 5682 8034 5694
rect 12786 5630 12798 5682
rect 12850 5630 12862 5682
rect 23874 5630 23886 5682
rect 23938 5630 23950 5682
rect 27346 5630 27358 5682
rect 27410 5679 27422 5682
rect 27697 5679 27743 5854
rect 41806 5842 41858 5854
rect 42142 5906 42194 5918
rect 42142 5842 42194 5854
rect 42590 5906 42642 5918
rect 42590 5842 42642 5854
rect 42814 5906 42866 5918
rect 47294 5906 47346 5918
rect 48862 5906 48914 5918
rect 43362 5854 43374 5906
rect 43426 5854 43438 5906
rect 47618 5854 47630 5906
rect 47682 5854 47694 5906
rect 42814 5842 42866 5854
rect 47294 5842 47346 5854
rect 48862 5842 48914 5854
rect 53230 5906 53282 5918
rect 55806 5906 55858 5918
rect 54786 5854 54798 5906
rect 54850 5854 54862 5906
rect 53230 5842 53282 5854
rect 55806 5842 55858 5854
rect 56030 5906 56082 5918
rect 59502 5906 59554 5918
rect 58930 5854 58942 5906
rect 58994 5854 59006 5906
rect 63074 5854 63086 5906
rect 63138 5854 63150 5906
rect 63746 5854 63758 5906
rect 63810 5854 63822 5906
rect 71250 5854 71262 5906
rect 71314 5854 71326 5906
rect 78082 5854 78094 5906
rect 78146 5854 78158 5906
rect 56030 5842 56082 5854
rect 59502 5842 59554 5854
rect 44830 5794 44882 5806
rect 48190 5794 48242 5806
rect 28130 5742 28142 5794
rect 28194 5742 28206 5794
rect 45378 5742 45390 5794
rect 45442 5742 45454 5794
rect 44830 5730 44882 5742
rect 48190 5730 48242 5742
rect 49310 5794 49362 5806
rect 51886 5794 51938 5806
rect 50194 5742 50206 5794
rect 50258 5742 50270 5794
rect 49310 5730 49362 5742
rect 51886 5730 51938 5742
rect 52782 5794 52834 5806
rect 52782 5730 52834 5742
rect 55918 5794 55970 5806
rect 55918 5730 55970 5742
rect 57598 5794 57650 5806
rect 57598 5730 57650 5742
rect 59950 5794 60002 5806
rect 62414 5794 62466 5806
rect 74510 5794 74562 5806
rect 60162 5742 60174 5794
rect 60226 5742 60238 5794
rect 60386 5742 60398 5794
rect 60450 5742 60462 5794
rect 62850 5742 62862 5794
rect 62914 5742 62926 5794
rect 67330 5742 67342 5794
rect 67394 5742 67406 5794
rect 70578 5742 70590 5794
rect 70642 5742 70654 5794
rect 59950 5730 60002 5742
rect 27410 5633 27743 5679
rect 30942 5682 30994 5694
rect 27410 5630 27422 5633
rect 7982 5618 8034 5630
rect 30942 5618 30994 5630
rect 34526 5682 34578 5694
rect 34526 5618 34578 5630
rect 37438 5682 37490 5694
rect 43810 5630 43822 5682
rect 43874 5679 43886 5682
rect 44258 5679 44270 5682
rect 43874 5633 44270 5679
rect 43874 5630 43886 5633
rect 44258 5630 44270 5633
rect 44322 5630 44334 5682
rect 52098 5630 52110 5682
rect 52162 5679 52174 5682
rect 52658 5679 52670 5682
rect 52162 5633 52670 5679
rect 52162 5630 52174 5633
rect 52658 5630 52670 5633
rect 52722 5630 52734 5682
rect 59378 5630 59390 5682
rect 59442 5679 59454 5682
rect 60177 5679 60223 5742
rect 62414 5730 62466 5742
rect 74510 5730 74562 5742
rect 59442 5633 60223 5679
rect 59442 5630 59454 5633
rect 37438 5618 37490 5630
rect 1344 5514 78624 5548
rect 1344 5462 10874 5514
rect 10926 5462 10978 5514
rect 11030 5462 11082 5514
rect 11134 5462 30194 5514
rect 30246 5462 30298 5514
rect 30350 5462 30402 5514
rect 30454 5462 49514 5514
rect 49566 5462 49618 5514
rect 49670 5462 49722 5514
rect 49774 5462 68834 5514
rect 68886 5462 68938 5514
rect 68990 5462 69042 5514
rect 69094 5462 78624 5514
rect 1344 5428 78624 5462
rect 17278 5346 17330 5358
rect 6738 5294 6750 5346
rect 6802 5294 6814 5346
rect 17278 5282 17330 5294
rect 21310 5346 21362 5358
rect 56254 5346 56306 5358
rect 22754 5294 22766 5346
rect 22818 5294 22830 5346
rect 25778 5294 25790 5346
rect 25842 5294 25854 5346
rect 37762 5294 37774 5346
rect 37826 5294 37838 5346
rect 45378 5294 45390 5346
rect 45442 5294 45454 5346
rect 47170 5294 47182 5346
rect 47234 5343 47246 5346
rect 47618 5343 47630 5346
rect 47234 5297 47630 5343
rect 47234 5294 47246 5297
rect 47618 5294 47630 5297
rect 47682 5294 47694 5346
rect 52658 5294 52670 5346
rect 52722 5294 52734 5346
rect 60386 5294 60398 5346
rect 60450 5343 60462 5346
rect 61058 5343 61070 5346
rect 60450 5297 61070 5343
rect 60450 5294 60462 5297
rect 61058 5294 61070 5297
rect 61122 5294 61134 5346
rect 21310 5282 21362 5294
rect 56254 5282 56306 5294
rect 2494 5234 2546 5246
rect 2494 5170 2546 5182
rect 3838 5234 3890 5246
rect 3838 5170 3890 5182
rect 5966 5234 6018 5246
rect 5966 5170 6018 5182
rect 6190 5234 6242 5246
rect 26910 5234 26962 5246
rect 30494 5234 30546 5246
rect 39454 5234 39506 5246
rect 46510 5234 46562 5246
rect 7074 5182 7086 5234
rect 7138 5182 7150 5234
rect 9202 5182 9214 5234
rect 9266 5182 9278 5234
rect 14466 5182 14478 5234
rect 14530 5182 14542 5234
rect 16594 5182 16606 5234
rect 16658 5182 16670 5234
rect 27346 5182 27358 5234
rect 27410 5182 27422 5234
rect 32946 5182 32958 5234
rect 33010 5182 33022 5234
rect 35186 5182 35198 5234
rect 35250 5182 35262 5234
rect 37874 5182 37886 5234
rect 37938 5182 37950 5234
rect 42690 5182 42702 5234
rect 42754 5182 42766 5234
rect 44034 5182 44046 5234
rect 44098 5182 44110 5234
rect 6190 5170 6242 5182
rect 26910 5170 26962 5182
rect 30494 5170 30546 5182
rect 39454 5170 39506 5182
rect 46510 5170 46562 5182
rect 46846 5234 46898 5246
rect 53230 5234 53282 5246
rect 52098 5182 52110 5234
rect 52162 5182 52174 5234
rect 46846 5170 46898 5182
rect 53230 5170 53282 5182
rect 53454 5234 53506 5246
rect 60622 5234 60674 5246
rect 70590 5234 70642 5246
rect 59714 5182 59726 5234
rect 59778 5182 59790 5234
rect 61506 5182 61518 5234
rect 61570 5182 61582 5234
rect 66098 5182 66110 5234
rect 66162 5182 66174 5234
rect 71250 5182 71262 5234
rect 71314 5182 71326 5234
rect 74050 5182 74062 5234
rect 74114 5182 74126 5234
rect 76178 5182 76190 5234
rect 76242 5182 76254 5234
rect 53454 5170 53506 5182
rect 60622 5170 60674 5182
rect 70590 5170 70642 5182
rect 2942 5122 2994 5134
rect 2942 5058 2994 5070
rect 3390 5122 3442 5134
rect 5070 5122 5122 5134
rect 4610 5070 4622 5122
rect 4674 5070 4686 5122
rect 3390 5058 3442 5070
rect 5070 5058 5122 5070
rect 6414 5122 6466 5134
rect 21422 5122 21474 5134
rect 22318 5122 22370 5134
rect 23438 5122 23490 5134
rect 9874 5070 9886 5122
rect 9938 5070 9950 5122
rect 12562 5070 12574 5122
rect 12626 5070 12638 5122
rect 13682 5070 13694 5122
rect 13746 5070 13758 5122
rect 16930 5070 16942 5122
rect 16994 5070 17006 5122
rect 19954 5070 19966 5122
rect 20018 5070 20030 5122
rect 20738 5070 20750 5122
rect 20802 5070 20814 5122
rect 21634 5070 21646 5122
rect 21698 5070 21710 5122
rect 21970 5070 21982 5122
rect 22034 5070 22046 5122
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 6414 5058 6466 5070
rect 21422 5058 21474 5070
rect 22318 5058 22370 5070
rect 23438 5058 23490 5070
rect 24670 5122 24722 5134
rect 25230 5122 25282 5134
rect 24994 5070 25006 5122
rect 25058 5070 25070 5122
rect 24670 5058 24722 5070
rect 25230 5058 25282 5070
rect 25342 5122 25394 5134
rect 25342 5058 25394 5070
rect 29262 5122 29314 5134
rect 30606 5122 30658 5134
rect 38446 5122 38498 5134
rect 44830 5122 44882 5134
rect 29810 5070 29822 5122
rect 29874 5070 29886 5122
rect 31378 5070 31390 5122
rect 31442 5070 31454 5122
rect 35970 5070 35982 5122
rect 36034 5070 36046 5122
rect 37202 5070 37214 5122
rect 37266 5070 37278 5122
rect 41346 5070 41358 5122
rect 41410 5070 41422 5122
rect 42242 5070 42254 5122
rect 42306 5070 42318 5122
rect 42914 5070 42926 5122
rect 42978 5070 42990 5122
rect 29262 5058 29314 5070
rect 30606 5058 30658 5070
rect 38446 5058 38498 5070
rect 44830 5058 44882 5070
rect 45054 5122 45106 5134
rect 45054 5058 45106 5070
rect 45950 5122 46002 5134
rect 45950 5058 46002 5070
rect 48302 5122 48354 5134
rect 48302 5058 48354 5070
rect 48638 5122 48690 5134
rect 48638 5058 48690 5070
rect 50318 5122 50370 5134
rect 50318 5058 50370 5070
rect 53006 5122 53058 5134
rect 53006 5058 53058 5070
rect 59390 5122 59442 5134
rect 59390 5058 59442 5070
rect 59502 5122 59554 5134
rect 61070 5122 61122 5134
rect 59938 5070 59950 5122
rect 60002 5070 60014 5122
rect 59502 5058 59554 5070
rect 61070 5058 61122 5070
rect 22206 5010 22258 5022
rect 22206 4946 22258 4958
rect 23326 5010 23378 5022
rect 23326 4946 23378 4958
rect 24334 5010 24386 5022
rect 29150 5010 29202 5022
rect 28242 4958 28254 5010
rect 28306 4958 28318 5010
rect 24334 4946 24386 4958
rect 29150 4946 29202 4958
rect 43486 5010 43538 5022
rect 43486 4946 43538 4958
rect 45614 5010 45666 5022
rect 47954 4958 47966 5010
rect 48018 4958 48030 5010
rect 48962 4958 48974 5010
rect 49026 4958 49038 5010
rect 51090 4958 51102 5010
rect 51154 4958 51166 5010
rect 55906 4958 55918 5010
rect 55970 4958 55982 5010
rect 58370 4958 58382 5010
rect 58434 4958 58446 5010
rect 62626 4958 62638 5010
rect 62690 4958 62702 5010
rect 65650 4958 65662 5010
rect 65714 4958 65726 5010
rect 67218 4958 67230 5010
rect 67282 4958 67294 5010
rect 68450 4958 68462 5010
rect 68514 4958 68526 5010
rect 73154 4958 73166 5010
rect 73218 4958 73230 5010
rect 74946 4958 74958 5010
rect 75010 4958 75022 5010
rect 77522 4958 77534 5010
rect 77586 4958 77598 5010
rect 45614 4946 45666 4958
rect 2046 4898 2098 4910
rect 2046 4834 2098 4846
rect 4286 4898 4338 4910
rect 4286 4834 4338 4846
rect 11902 4898 11954 4910
rect 11902 4834 11954 4846
rect 17166 4898 17218 4910
rect 26350 4898 26402 4910
rect 42478 4898 42530 4910
rect 17714 4846 17726 4898
rect 17778 4846 17790 4898
rect 23874 4846 23886 4898
rect 23938 4846 23950 4898
rect 38770 4846 38782 4898
rect 38834 4846 38846 4898
rect 17166 4834 17218 4846
rect 26350 4834 26402 4846
rect 42478 4834 42530 4846
rect 42702 4898 42754 4910
rect 42702 4834 42754 4846
rect 43710 4898 43762 4910
rect 43710 4834 43762 4846
rect 43934 4898 43986 4910
rect 43934 4834 43986 4846
rect 44046 4898 44098 4910
rect 44046 4834 44098 4846
rect 45838 4898 45890 4910
rect 45838 4834 45890 4846
rect 47294 4898 47346 4910
rect 47294 4834 47346 4846
rect 49422 4898 49474 4910
rect 49422 4834 49474 4846
rect 49870 4898 49922 4910
rect 49870 4834 49922 4846
rect 59726 4898 59778 4910
rect 59726 4834 59778 4846
rect 63198 4898 63250 4910
rect 63198 4834 63250 4846
rect 77982 4898 78034 4910
rect 77982 4834 78034 4846
rect 1344 4730 78784 4764
rect 1344 4678 20534 4730
rect 20586 4678 20638 4730
rect 20690 4678 20742 4730
rect 20794 4678 39854 4730
rect 39906 4678 39958 4730
rect 40010 4678 40062 4730
rect 40114 4678 59174 4730
rect 59226 4678 59278 4730
rect 59330 4678 59382 4730
rect 59434 4678 78494 4730
rect 78546 4678 78598 4730
rect 78650 4678 78702 4730
rect 78754 4678 78784 4730
rect 1344 4644 78784 4678
rect 2494 4562 2546 4574
rect 2494 4498 2546 4510
rect 10670 4562 10722 4574
rect 10670 4498 10722 4510
rect 17838 4562 17890 4574
rect 17838 4498 17890 4510
rect 24222 4562 24274 4574
rect 24222 4498 24274 4510
rect 27694 4562 27746 4574
rect 27694 4498 27746 4510
rect 44158 4562 44210 4574
rect 44158 4498 44210 4510
rect 44830 4562 44882 4574
rect 44830 4498 44882 4510
rect 48638 4562 48690 4574
rect 48638 4498 48690 4510
rect 51662 4562 51714 4574
rect 51662 4498 51714 4510
rect 51774 4562 51826 4574
rect 51774 4498 51826 4510
rect 52334 4562 52386 4574
rect 52334 4498 52386 4510
rect 54350 4562 54402 4574
rect 54350 4498 54402 4510
rect 72158 4562 72210 4574
rect 72158 4498 72210 4510
rect 17390 4450 17442 4462
rect 13010 4398 13022 4450
rect 13074 4398 13086 4450
rect 17390 4386 17442 4398
rect 17614 4450 17666 4462
rect 22206 4450 22258 4462
rect 18946 4398 18958 4450
rect 19010 4398 19022 4450
rect 17614 4386 17666 4398
rect 22206 4386 22258 4398
rect 22542 4450 22594 4462
rect 22542 4386 22594 4398
rect 23326 4450 23378 4462
rect 23326 4386 23378 4398
rect 23438 4450 23490 4462
rect 23438 4386 23490 4398
rect 25902 4450 25954 4462
rect 25902 4386 25954 4398
rect 26798 4450 26850 4462
rect 33182 4450 33234 4462
rect 29138 4398 29150 4450
rect 29202 4398 29214 4450
rect 26798 4386 26850 4398
rect 33182 4386 33234 4398
rect 34526 4450 34578 4462
rect 52222 4450 52274 4462
rect 47954 4398 47966 4450
rect 48018 4398 48030 4450
rect 50978 4398 50990 4450
rect 51042 4398 51054 4450
rect 34526 4386 34578 4398
rect 52222 4386 52274 4398
rect 55470 4450 55522 4462
rect 55470 4386 55522 4398
rect 55806 4450 55858 4462
rect 55806 4386 55858 4398
rect 56814 4450 56866 4462
rect 56814 4386 56866 4398
rect 57038 4450 57090 4462
rect 77870 4450 77922 4462
rect 58594 4398 58606 4450
rect 58658 4398 58670 4450
rect 61730 4398 61742 4450
rect 61794 4398 61806 4450
rect 62514 4398 62526 4450
rect 62578 4398 62590 4450
rect 64530 4398 64542 4450
rect 64594 4398 64606 4450
rect 67666 4398 67678 4450
rect 67730 4398 67742 4450
rect 71026 4398 71038 4450
rect 71090 4398 71102 4450
rect 74274 4398 74286 4450
rect 74338 4398 74350 4450
rect 75170 4398 75182 4450
rect 75234 4398 75246 4450
rect 57038 4386 57090 4398
rect 77870 4386 77922 4398
rect 78206 4450 78258 4462
rect 78206 4386 78258 4398
rect 9550 4338 9602 4350
rect 18062 4338 18114 4350
rect 24558 4338 24610 4350
rect 26350 4338 26402 4350
rect 2258 4286 2270 4338
rect 2322 4286 2334 4338
rect 5618 4286 5630 4338
rect 5682 4286 5694 4338
rect 8978 4286 8990 4338
rect 9042 4286 9054 4338
rect 13682 4286 13694 4338
rect 13746 4286 13758 4338
rect 16706 4286 16718 4338
rect 16770 4286 16782 4338
rect 18722 4286 18734 4338
rect 18786 4286 18798 4338
rect 21522 4286 21534 4338
rect 21586 4286 21598 4338
rect 23090 4286 23102 4338
rect 23154 4286 23166 4338
rect 26114 4286 26126 4338
rect 26178 4286 26190 4338
rect 9550 4274 9602 4286
rect 18062 4274 18114 4286
rect 24558 4274 24610 4286
rect 26350 4274 26402 4286
rect 26574 4338 26626 4350
rect 44046 4338 44098 4350
rect 29922 4286 29934 4338
rect 29986 4286 29998 4338
rect 33954 4286 33966 4338
rect 34018 4286 34030 4338
rect 34850 4286 34862 4338
rect 34914 4286 34926 4338
rect 40338 4286 40350 4338
rect 40402 4286 40414 4338
rect 43026 4286 43038 4338
rect 43090 4286 43102 4338
rect 43810 4286 43822 4338
rect 43874 4286 43886 4338
rect 26574 4274 26626 4286
rect 44046 4274 44098 4286
rect 44270 4338 44322 4350
rect 44270 4274 44322 4286
rect 44382 4338 44434 4350
rect 44382 4274 44434 4286
rect 45054 4338 45106 4350
rect 52110 4338 52162 4350
rect 45378 4286 45390 4338
rect 45442 4286 45454 4338
rect 45054 4274 45106 4286
rect 52110 4274 52162 4286
rect 52782 4338 52834 4350
rect 52782 4274 52834 4286
rect 53342 4338 53394 4350
rect 54798 4338 54850 4350
rect 53890 4286 53902 4338
rect 53954 4286 53966 4338
rect 53342 4274 53394 4286
rect 54798 4274 54850 4286
rect 55246 4338 55298 4350
rect 55246 4274 55298 4286
rect 1934 4226 1986 4238
rect 1934 4162 1986 4174
rect 3278 4226 3330 4238
rect 25678 4226 25730 4238
rect 4834 4174 4846 4226
rect 4898 4174 4910 4226
rect 7858 4174 7870 4226
rect 7922 4174 7934 4226
rect 10882 4174 10894 4226
rect 10946 4174 10958 4226
rect 15698 4174 15710 4226
rect 15762 4174 15774 4226
rect 3278 4162 3330 4174
rect 25678 4162 25730 4174
rect 26686 4226 26738 4238
rect 44942 4226 44994 4238
rect 27234 4174 27246 4226
rect 27298 4174 27310 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 32162 4174 32174 4226
rect 32226 4174 32238 4226
rect 33618 4174 33630 4226
rect 33682 4174 33694 4226
rect 36194 4174 36206 4226
rect 36258 4174 36270 4226
rect 38322 4174 38334 4226
rect 38386 4174 38398 4226
rect 26686 4162 26738 4174
rect 44942 4162 44994 4174
rect 52558 4226 52610 4238
rect 66670 4226 66722 4238
rect 56690 4174 56702 4226
rect 56754 4174 56766 4226
rect 57586 4174 57598 4226
rect 57650 4174 57662 4226
rect 63858 4174 63870 4226
rect 63922 4174 63934 4226
rect 52558 4162 52610 4174
rect 66670 4162 66722 4174
rect 69470 4226 69522 4238
rect 77310 4226 77362 4238
rect 70242 4174 70254 4226
rect 70306 4174 70318 4226
rect 69470 4162 69522 4174
rect 77310 4162 77362 4174
rect 9774 4114 9826 4126
rect 19518 4114 19570 4126
rect 41134 4114 41186 4126
rect 10098 4062 10110 4114
rect 10162 4062 10174 4114
rect 23874 4062 23886 4114
rect 23938 4062 23950 4114
rect 9774 4050 9826 4062
rect 19518 4050 19570 4062
rect 41134 4050 41186 4062
rect 45614 4114 45666 4126
rect 45614 4050 45666 4062
rect 53566 4114 53618 4126
rect 53566 4050 53618 4062
rect 55022 4114 55074 4126
rect 55022 4050 55074 4062
rect 59278 4114 59330 4126
rect 59278 4050 59330 4062
rect 1344 3946 78624 3980
rect 1344 3894 10874 3946
rect 10926 3894 10978 3946
rect 11030 3894 11082 3946
rect 11134 3894 30194 3946
rect 30246 3894 30298 3946
rect 30350 3894 30402 3946
rect 30454 3894 49514 3946
rect 49566 3894 49618 3946
rect 49670 3894 49722 3946
rect 49774 3894 68834 3946
rect 68886 3894 68938 3946
rect 68990 3894 69042 3946
rect 69094 3894 78624 3946
rect 1344 3860 78624 3894
rect 26126 3778 26178 3790
rect 26126 3714 26178 3726
rect 27358 3778 27410 3790
rect 27358 3714 27410 3726
rect 32510 3778 32562 3790
rect 44606 3778 44658 3790
rect 43698 3726 43710 3778
rect 43762 3726 43774 3778
rect 32510 3714 32562 3726
rect 44606 3714 44658 3726
rect 59166 3778 59218 3790
rect 59166 3714 59218 3726
rect 59390 3778 59442 3790
rect 59390 3714 59442 3726
rect 65326 3778 65378 3790
rect 65326 3714 65378 3726
rect 66334 3778 66386 3790
rect 66334 3714 66386 3726
rect 4958 3666 5010 3678
rect 4958 3602 5010 3614
rect 7758 3666 7810 3678
rect 7758 3602 7810 3614
rect 11566 3666 11618 3678
rect 11566 3602 11618 3614
rect 17614 3666 17666 3678
rect 27582 3666 27634 3678
rect 21858 3614 21870 3666
rect 21922 3614 21934 3666
rect 17614 3602 17666 3614
rect 27582 3602 27634 3614
rect 31390 3666 31442 3678
rect 31390 3602 31442 3614
rect 32398 3666 32450 3678
rect 32398 3602 32450 3614
rect 34414 3666 34466 3678
rect 34414 3602 34466 3614
rect 40686 3666 40738 3678
rect 46510 3666 46562 3678
rect 52222 3666 52274 3678
rect 44146 3614 44158 3666
rect 44210 3614 44222 3666
rect 48402 3614 48414 3666
rect 48466 3614 48478 3666
rect 51874 3614 51886 3666
rect 51938 3614 51950 3666
rect 40686 3602 40738 3614
rect 46510 3602 46562 3614
rect 52222 3602 52274 3614
rect 52558 3666 52610 3678
rect 52558 3602 52610 3614
rect 52670 3666 52722 3678
rect 52670 3602 52722 3614
rect 53230 3666 53282 3678
rect 55470 3666 55522 3678
rect 53666 3614 53678 3666
rect 53730 3614 53742 3666
rect 53230 3602 53282 3614
rect 55470 3602 55522 3614
rect 55918 3666 55970 3678
rect 55918 3602 55970 3614
rect 56926 3666 56978 3678
rect 56926 3602 56978 3614
rect 57598 3666 57650 3678
rect 57598 3602 57650 3614
rect 61070 3666 61122 3678
rect 72594 3614 72606 3666
rect 72658 3614 72670 3666
rect 61070 3602 61122 3614
rect 4062 3554 4114 3566
rect 9326 3554 9378 3566
rect 13134 3554 13186 3566
rect 23662 3554 23714 3566
rect 2258 3502 2270 3554
rect 2322 3502 2334 3554
rect 3602 3502 3614 3554
rect 3666 3502 3678 3554
rect 4498 3502 4510 3554
rect 4562 3502 4574 3554
rect 5618 3502 5630 3554
rect 5682 3502 5694 3554
rect 8754 3502 8766 3554
rect 8818 3502 8830 3554
rect 12562 3502 12574 3554
rect 12626 3502 12638 3554
rect 16258 3502 16270 3554
rect 16322 3502 16334 3554
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 4062 3490 4114 3502
rect 9326 3490 9378 3502
rect 13134 3490 13186 3502
rect 23662 3490 23714 3502
rect 25006 3554 25058 3566
rect 25006 3490 25058 3502
rect 25566 3554 25618 3566
rect 26350 3554 26402 3566
rect 25890 3502 25902 3554
rect 25954 3502 25966 3554
rect 25566 3490 25618 3502
rect 26350 3490 26402 3502
rect 26574 3554 26626 3566
rect 27806 3554 27858 3566
rect 43934 3554 43986 3566
rect 46174 3554 46226 3566
rect 26898 3502 26910 3554
rect 26962 3502 26974 3554
rect 27122 3502 27134 3554
rect 27186 3502 27198 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 29026 3502 29038 3554
rect 29090 3502 29102 3554
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 38770 3502 38782 3554
rect 38834 3502 38846 3554
rect 42578 3502 42590 3554
rect 42642 3502 42654 3554
rect 45154 3502 45166 3554
rect 45218 3502 45230 3554
rect 26574 3490 26626 3502
rect 27806 3490 27858 3502
rect 43934 3490 43986 3502
rect 46174 3490 46226 3502
rect 46846 3554 46898 3566
rect 46846 3490 46898 3502
rect 47406 3554 47458 3566
rect 53566 3554 53618 3566
rect 50418 3502 50430 3554
rect 50482 3502 50494 3554
rect 52882 3502 52894 3554
rect 52946 3502 52958 3554
rect 47406 3490 47458 3502
rect 53566 3490 53618 3502
rect 55358 3554 55410 3566
rect 55358 3490 55410 3502
rect 55694 3554 55746 3566
rect 60174 3554 60226 3566
rect 56242 3502 56254 3554
rect 56306 3502 56318 3554
rect 57922 3502 57934 3554
rect 57986 3502 57998 3554
rect 59602 3502 59614 3554
rect 59666 3502 59678 3554
rect 59938 3502 59950 3554
rect 60002 3502 60014 3554
rect 55694 3490 55746 3502
rect 60174 3490 60226 3502
rect 60398 3554 60450 3566
rect 60958 3554 61010 3566
rect 60610 3502 60622 3554
rect 60674 3502 60686 3554
rect 60398 3490 60450 3502
rect 60958 3490 61010 3502
rect 61182 3554 61234 3566
rect 61182 3490 61234 3502
rect 61406 3554 61458 3566
rect 65762 3502 65774 3554
rect 65826 3502 65838 3554
rect 69458 3502 69470 3554
rect 69522 3502 69534 3554
rect 77074 3502 77086 3554
rect 77138 3502 77150 3554
rect 78082 3502 78094 3554
rect 78146 3502 78158 3554
rect 61406 3490 61458 3502
rect 1934 3442 1986 3454
rect 1934 3378 1986 3390
rect 2494 3442 2546 3454
rect 2494 3378 2546 3390
rect 2830 3442 2882 3454
rect 25342 3442 25394 3454
rect 14802 3390 14814 3442
rect 14866 3390 14878 3442
rect 23986 3390 23998 3442
rect 24050 3390 24062 3442
rect 2830 3378 2882 3390
rect 25342 3378 25394 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 32286 3442 32338 3454
rect 36318 3442 36370 3454
rect 46286 3442 46338 3454
rect 51998 3442 52050 3454
rect 35970 3390 35982 3442
rect 36034 3390 36046 3442
rect 37650 3390 37662 3442
rect 37714 3390 37726 3442
rect 47730 3390 47742 3442
rect 47794 3390 47806 3442
rect 49634 3390 49646 3442
rect 49698 3390 49710 3442
rect 51202 3390 51214 3442
rect 51266 3390 51278 3442
rect 32286 3378 32338 3390
rect 36318 3378 36370 3390
rect 46286 3378 46338 3390
rect 51998 3378 52050 3390
rect 55022 3442 55074 3454
rect 55022 3378 55074 3390
rect 56702 3442 56754 3454
rect 56702 3378 56754 3390
rect 57374 3442 57426 3454
rect 57374 3378 57426 3390
rect 60286 3442 60338 3454
rect 65550 3442 65602 3454
rect 73502 3442 73554 3454
rect 62850 3390 62862 3442
rect 62914 3390 62926 3442
rect 68450 3390 68462 3442
rect 68514 3390 68526 3442
rect 70354 3390 70366 3442
rect 70418 3390 70430 3442
rect 60286 3378 60338 3390
rect 65550 3378 65602 3390
rect 73502 3378 73554 3390
rect 73950 3442 74002 3454
rect 76862 3442 76914 3454
rect 76066 3390 76078 3442
rect 76130 3390 76142 3442
rect 73950 3378 74002 3390
rect 76862 3378 76914 3390
rect 77870 3442 77922 3454
rect 77870 3378 77922 3390
rect 3166 3330 3218 3342
rect 13470 3330 13522 3342
rect 5842 3278 5854 3330
rect 5906 3278 5918 3330
rect 9650 3278 9662 3330
rect 9714 3278 9726 3330
rect 3166 3266 3218 3278
rect 13470 3266 13522 3278
rect 17054 3330 17106 3342
rect 17054 3266 17106 3278
rect 24670 3330 24722 3342
rect 24670 3266 24722 3278
rect 26686 3330 26738 3342
rect 26686 3266 26738 3278
rect 27918 3330 27970 3342
rect 27918 3266 27970 3278
rect 40014 3330 40066 3342
rect 40014 3266 40066 3278
rect 44718 3330 44770 3342
rect 44718 3266 44770 3278
rect 44942 3330 44994 3342
rect 44942 3266 44994 3278
rect 45726 3330 45778 3342
rect 45726 3266 45778 3278
rect 45838 3330 45890 3342
rect 45838 3266 45890 3278
rect 46958 3330 47010 3342
rect 51550 3330 51602 3342
rect 50194 3278 50206 3330
rect 50258 3278 50270 3330
rect 46958 3266 47010 3278
rect 51550 3266 51602 3278
rect 54574 3330 54626 3342
rect 54574 3266 54626 3278
rect 56030 3330 56082 3342
rect 56030 3266 56082 3278
rect 56814 3330 56866 3342
rect 56814 3266 56866 3278
rect 59502 3330 59554 3342
rect 59502 3266 59554 3278
rect 61966 3330 62018 3342
rect 61966 3266 62018 3278
rect 69246 3330 69298 3342
rect 73154 3278 73166 3330
rect 73218 3278 73230 3330
rect 69246 3266 69298 3278
rect 1344 3162 78784 3196
rect 1344 3110 20534 3162
rect 20586 3110 20638 3162
rect 20690 3110 20742 3162
rect 20794 3110 39854 3162
rect 39906 3110 39958 3162
rect 40010 3110 40062 3162
rect 40114 3110 59174 3162
rect 59226 3110 59278 3162
rect 59330 3110 59382 3162
rect 59434 3110 78494 3162
rect 78546 3110 78598 3162
rect 78650 3110 78702 3162
rect 78754 3110 78784 3162
rect 1344 3076 78784 3110
rect 25442 2942 25454 2994
rect 25506 2991 25518 2994
rect 29138 2991 29150 2994
rect 25506 2945 29150 2991
rect 25506 2942 25518 2945
rect 29138 2942 29150 2945
rect 29202 2942 29214 2994
rect 43362 2942 43374 2994
rect 43426 2991 43438 2994
rect 47170 2991 47182 2994
rect 43426 2945 47182 2991
rect 43426 2942 43438 2945
rect 47170 2942 47182 2945
rect 47234 2942 47246 2994
rect 67442 2942 67454 2994
rect 67506 2991 67518 2994
rect 68002 2991 68014 2994
rect 67506 2945 68014 2991
rect 67506 2942 67518 2945
rect 68002 2942 68014 2945
rect 68066 2942 68078 2994
rect 38882 2830 38894 2882
rect 38946 2879 38958 2882
rect 40226 2879 40238 2882
rect 38946 2833 40238 2879
rect 38946 2830 38958 2833
rect 40226 2830 40238 2833
rect 40290 2879 40302 2882
rect 40290 2833 46335 2879
rect 40290 2830 40302 2833
rect 46289 2770 46335 2833
rect 61394 2830 61406 2882
rect 61458 2879 61470 2882
rect 67330 2879 67342 2882
rect 61458 2833 67342 2879
rect 61458 2830 61470 2833
rect 67330 2830 67342 2833
rect 67394 2830 67406 2882
rect 42914 2718 42926 2770
rect 42978 2767 42990 2770
rect 45490 2767 45502 2770
rect 42978 2721 45502 2767
rect 42978 2718 42990 2721
rect 45490 2718 45502 2721
rect 45554 2718 45566 2770
rect 46274 2718 46286 2770
rect 46338 2718 46350 2770
rect 62738 2718 62750 2770
rect 62802 2767 62814 2770
rect 65986 2767 65998 2770
rect 62802 2721 65998 2767
rect 62802 2718 62814 2721
rect 65986 2718 65998 2721
rect 66050 2767 66062 2770
rect 68450 2767 68462 2770
rect 66050 2721 68462 2767
rect 66050 2718 66062 2721
rect 68450 2718 68462 2721
rect 68514 2718 68526 2770
rect 42802 2606 42814 2658
rect 42866 2655 42878 2658
rect 43698 2655 43710 2658
rect 42866 2609 43710 2655
rect 42866 2606 42878 2609
rect 43698 2606 43710 2609
rect 43762 2606 43774 2658
rect 66098 2606 66110 2658
rect 66162 2655 66174 2658
rect 70242 2655 70254 2658
rect 66162 2609 70254 2655
rect 66162 2606 66174 2609
rect 70242 2606 70254 2609
rect 70306 2606 70318 2658
rect 43250 2494 43262 2546
rect 43314 2543 43326 2546
rect 44370 2543 44382 2546
rect 43314 2497 44382 2543
rect 43314 2494 43326 2497
rect 44370 2494 44382 2497
rect 44434 2494 44446 2546
rect 45378 2494 45390 2546
rect 45442 2543 45454 2546
rect 54338 2543 54350 2546
rect 45442 2497 54350 2543
rect 45442 2494 45454 2497
rect 54338 2494 54350 2497
rect 54402 2494 54414 2546
rect 46050 2382 46062 2434
rect 46114 2431 46126 2434
rect 54562 2431 54574 2434
rect 46114 2385 54574 2431
rect 46114 2382 46126 2385
rect 54562 2382 54574 2385
rect 54626 2382 54638 2434
rect 45714 2270 45726 2322
rect 45778 2319 45790 2322
rect 50866 2319 50878 2322
rect 45778 2273 50878 2319
rect 45778 2270 45790 2273
rect 50866 2270 50878 2273
rect 50930 2270 50942 2322
rect 61618 1822 61630 1874
rect 61682 1871 61694 1874
rect 64418 1871 64430 1874
rect 61682 1825 64430 1871
rect 61682 1822 61694 1825
rect 64418 1822 64430 1825
rect 64482 1822 64494 1874
rect 42354 926 42366 978
rect 42418 975 42430 978
rect 45826 975 45838 978
rect 42418 929 45838 975
rect 42418 926 42430 929
rect 45826 926 45838 929
rect 45890 926 45902 978
<< via1 >>
rect 10874 36822 10926 36874
rect 10978 36822 11030 36874
rect 11082 36822 11134 36874
rect 30194 36822 30246 36874
rect 30298 36822 30350 36874
rect 30402 36822 30454 36874
rect 49514 36822 49566 36874
rect 49618 36822 49670 36874
rect 49722 36822 49774 36874
rect 68834 36822 68886 36874
rect 68938 36822 68990 36874
rect 69042 36822 69094 36874
rect 20534 36038 20586 36090
rect 20638 36038 20690 36090
rect 20742 36038 20794 36090
rect 39854 36038 39906 36090
rect 39958 36038 40010 36090
rect 40062 36038 40114 36090
rect 59174 36038 59226 36090
rect 59278 36038 59330 36090
rect 59382 36038 59434 36090
rect 78494 36038 78546 36090
rect 78598 36038 78650 36090
rect 78702 36038 78754 36090
rect 10874 35254 10926 35306
rect 10978 35254 11030 35306
rect 11082 35254 11134 35306
rect 30194 35254 30246 35306
rect 30298 35254 30350 35306
rect 30402 35254 30454 35306
rect 49514 35254 49566 35306
rect 49618 35254 49670 35306
rect 49722 35254 49774 35306
rect 68834 35254 68886 35306
rect 68938 35254 68990 35306
rect 69042 35254 69094 35306
rect 20534 34470 20586 34522
rect 20638 34470 20690 34522
rect 20742 34470 20794 34522
rect 39854 34470 39906 34522
rect 39958 34470 40010 34522
rect 40062 34470 40114 34522
rect 59174 34470 59226 34522
rect 59278 34470 59330 34522
rect 59382 34470 59434 34522
rect 78494 34470 78546 34522
rect 78598 34470 78650 34522
rect 78702 34470 78754 34522
rect 10874 33686 10926 33738
rect 10978 33686 11030 33738
rect 11082 33686 11134 33738
rect 30194 33686 30246 33738
rect 30298 33686 30350 33738
rect 30402 33686 30454 33738
rect 49514 33686 49566 33738
rect 49618 33686 49670 33738
rect 49722 33686 49774 33738
rect 68834 33686 68886 33738
rect 68938 33686 68990 33738
rect 69042 33686 69094 33738
rect 20534 32902 20586 32954
rect 20638 32902 20690 32954
rect 20742 32902 20794 32954
rect 39854 32902 39906 32954
rect 39958 32902 40010 32954
rect 40062 32902 40114 32954
rect 59174 32902 59226 32954
rect 59278 32902 59330 32954
rect 59382 32902 59434 32954
rect 78494 32902 78546 32954
rect 78598 32902 78650 32954
rect 78702 32902 78754 32954
rect 10874 32118 10926 32170
rect 10978 32118 11030 32170
rect 11082 32118 11134 32170
rect 30194 32118 30246 32170
rect 30298 32118 30350 32170
rect 30402 32118 30454 32170
rect 49514 32118 49566 32170
rect 49618 32118 49670 32170
rect 49722 32118 49774 32170
rect 68834 32118 68886 32170
rect 68938 32118 68990 32170
rect 69042 32118 69094 32170
rect 20534 31334 20586 31386
rect 20638 31334 20690 31386
rect 20742 31334 20794 31386
rect 39854 31334 39906 31386
rect 39958 31334 40010 31386
rect 40062 31334 40114 31386
rect 59174 31334 59226 31386
rect 59278 31334 59330 31386
rect 59382 31334 59434 31386
rect 78494 31334 78546 31386
rect 78598 31334 78650 31386
rect 78702 31334 78754 31386
rect 10874 30550 10926 30602
rect 10978 30550 11030 30602
rect 11082 30550 11134 30602
rect 30194 30550 30246 30602
rect 30298 30550 30350 30602
rect 30402 30550 30454 30602
rect 49514 30550 49566 30602
rect 49618 30550 49670 30602
rect 49722 30550 49774 30602
rect 68834 30550 68886 30602
rect 68938 30550 68990 30602
rect 69042 30550 69094 30602
rect 20534 29766 20586 29818
rect 20638 29766 20690 29818
rect 20742 29766 20794 29818
rect 39854 29766 39906 29818
rect 39958 29766 40010 29818
rect 40062 29766 40114 29818
rect 59174 29766 59226 29818
rect 59278 29766 59330 29818
rect 59382 29766 59434 29818
rect 78494 29766 78546 29818
rect 78598 29766 78650 29818
rect 78702 29766 78754 29818
rect 10874 28982 10926 29034
rect 10978 28982 11030 29034
rect 11082 28982 11134 29034
rect 30194 28982 30246 29034
rect 30298 28982 30350 29034
rect 30402 28982 30454 29034
rect 49514 28982 49566 29034
rect 49618 28982 49670 29034
rect 49722 28982 49774 29034
rect 68834 28982 68886 29034
rect 68938 28982 68990 29034
rect 69042 28982 69094 29034
rect 20534 28198 20586 28250
rect 20638 28198 20690 28250
rect 20742 28198 20794 28250
rect 39854 28198 39906 28250
rect 39958 28198 40010 28250
rect 40062 28198 40114 28250
rect 59174 28198 59226 28250
rect 59278 28198 59330 28250
rect 59382 28198 59434 28250
rect 78494 28198 78546 28250
rect 78598 28198 78650 28250
rect 78702 28198 78754 28250
rect 10874 27414 10926 27466
rect 10978 27414 11030 27466
rect 11082 27414 11134 27466
rect 30194 27414 30246 27466
rect 30298 27414 30350 27466
rect 30402 27414 30454 27466
rect 49514 27414 49566 27466
rect 49618 27414 49670 27466
rect 49722 27414 49774 27466
rect 68834 27414 68886 27466
rect 68938 27414 68990 27466
rect 69042 27414 69094 27466
rect 20534 26630 20586 26682
rect 20638 26630 20690 26682
rect 20742 26630 20794 26682
rect 39854 26630 39906 26682
rect 39958 26630 40010 26682
rect 40062 26630 40114 26682
rect 59174 26630 59226 26682
rect 59278 26630 59330 26682
rect 59382 26630 59434 26682
rect 78494 26630 78546 26682
rect 78598 26630 78650 26682
rect 78702 26630 78754 26682
rect 10874 25846 10926 25898
rect 10978 25846 11030 25898
rect 11082 25846 11134 25898
rect 30194 25846 30246 25898
rect 30298 25846 30350 25898
rect 30402 25846 30454 25898
rect 49514 25846 49566 25898
rect 49618 25846 49670 25898
rect 49722 25846 49774 25898
rect 68834 25846 68886 25898
rect 68938 25846 68990 25898
rect 69042 25846 69094 25898
rect 20534 25062 20586 25114
rect 20638 25062 20690 25114
rect 20742 25062 20794 25114
rect 39854 25062 39906 25114
rect 39958 25062 40010 25114
rect 40062 25062 40114 25114
rect 59174 25062 59226 25114
rect 59278 25062 59330 25114
rect 59382 25062 59434 25114
rect 78494 25062 78546 25114
rect 78598 25062 78650 25114
rect 78702 25062 78754 25114
rect 10874 24278 10926 24330
rect 10978 24278 11030 24330
rect 11082 24278 11134 24330
rect 30194 24278 30246 24330
rect 30298 24278 30350 24330
rect 30402 24278 30454 24330
rect 49514 24278 49566 24330
rect 49618 24278 49670 24330
rect 49722 24278 49774 24330
rect 68834 24278 68886 24330
rect 68938 24278 68990 24330
rect 69042 24278 69094 24330
rect 20534 23494 20586 23546
rect 20638 23494 20690 23546
rect 20742 23494 20794 23546
rect 39854 23494 39906 23546
rect 39958 23494 40010 23546
rect 40062 23494 40114 23546
rect 59174 23494 59226 23546
rect 59278 23494 59330 23546
rect 59382 23494 59434 23546
rect 78494 23494 78546 23546
rect 78598 23494 78650 23546
rect 78702 23494 78754 23546
rect 10874 22710 10926 22762
rect 10978 22710 11030 22762
rect 11082 22710 11134 22762
rect 30194 22710 30246 22762
rect 30298 22710 30350 22762
rect 30402 22710 30454 22762
rect 49514 22710 49566 22762
rect 49618 22710 49670 22762
rect 49722 22710 49774 22762
rect 68834 22710 68886 22762
rect 68938 22710 68990 22762
rect 69042 22710 69094 22762
rect 20534 21926 20586 21978
rect 20638 21926 20690 21978
rect 20742 21926 20794 21978
rect 39854 21926 39906 21978
rect 39958 21926 40010 21978
rect 40062 21926 40114 21978
rect 59174 21926 59226 21978
rect 59278 21926 59330 21978
rect 59382 21926 59434 21978
rect 78494 21926 78546 21978
rect 78598 21926 78650 21978
rect 78702 21926 78754 21978
rect 10874 21142 10926 21194
rect 10978 21142 11030 21194
rect 11082 21142 11134 21194
rect 30194 21142 30246 21194
rect 30298 21142 30350 21194
rect 30402 21142 30454 21194
rect 49514 21142 49566 21194
rect 49618 21142 49670 21194
rect 49722 21142 49774 21194
rect 68834 21142 68886 21194
rect 68938 21142 68990 21194
rect 69042 21142 69094 21194
rect 20534 20358 20586 20410
rect 20638 20358 20690 20410
rect 20742 20358 20794 20410
rect 39854 20358 39906 20410
rect 39958 20358 40010 20410
rect 40062 20358 40114 20410
rect 59174 20358 59226 20410
rect 59278 20358 59330 20410
rect 59382 20358 59434 20410
rect 78494 20358 78546 20410
rect 78598 20358 78650 20410
rect 78702 20358 78754 20410
rect 10874 19574 10926 19626
rect 10978 19574 11030 19626
rect 11082 19574 11134 19626
rect 30194 19574 30246 19626
rect 30298 19574 30350 19626
rect 30402 19574 30454 19626
rect 49514 19574 49566 19626
rect 49618 19574 49670 19626
rect 49722 19574 49774 19626
rect 68834 19574 68886 19626
rect 68938 19574 68990 19626
rect 69042 19574 69094 19626
rect 20534 18790 20586 18842
rect 20638 18790 20690 18842
rect 20742 18790 20794 18842
rect 39854 18790 39906 18842
rect 39958 18790 40010 18842
rect 40062 18790 40114 18842
rect 59174 18790 59226 18842
rect 59278 18790 59330 18842
rect 59382 18790 59434 18842
rect 78494 18790 78546 18842
rect 78598 18790 78650 18842
rect 78702 18790 78754 18842
rect 10874 18006 10926 18058
rect 10978 18006 11030 18058
rect 11082 18006 11134 18058
rect 30194 18006 30246 18058
rect 30298 18006 30350 18058
rect 30402 18006 30454 18058
rect 49514 18006 49566 18058
rect 49618 18006 49670 18058
rect 49722 18006 49774 18058
rect 68834 18006 68886 18058
rect 68938 18006 68990 18058
rect 69042 18006 69094 18058
rect 20534 17222 20586 17274
rect 20638 17222 20690 17274
rect 20742 17222 20794 17274
rect 39854 17222 39906 17274
rect 39958 17222 40010 17274
rect 40062 17222 40114 17274
rect 59174 17222 59226 17274
rect 59278 17222 59330 17274
rect 59382 17222 59434 17274
rect 78494 17222 78546 17274
rect 78598 17222 78650 17274
rect 78702 17222 78754 17274
rect 10874 16438 10926 16490
rect 10978 16438 11030 16490
rect 11082 16438 11134 16490
rect 30194 16438 30246 16490
rect 30298 16438 30350 16490
rect 30402 16438 30454 16490
rect 49514 16438 49566 16490
rect 49618 16438 49670 16490
rect 49722 16438 49774 16490
rect 68834 16438 68886 16490
rect 68938 16438 68990 16490
rect 69042 16438 69094 16490
rect 20534 15654 20586 15706
rect 20638 15654 20690 15706
rect 20742 15654 20794 15706
rect 39854 15654 39906 15706
rect 39958 15654 40010 15706
rect 40062 15654 40114 15706
rect 59174 15654 59226 15706
rect 59278 15654 59330 15706
rect 59382 15654 59434 15706
rect 78494 15654 78546 15706
rect 78598 15654 78650 15706
rect 78702 15654 78754 15706
rect 35758 15374 35810 15426
rect 34750 15150 34802 15202
rect 10874 14870 10926 14922
rect 10978 14870 11030 14922
rect 11082 14870 11134 14922
rect 30194 14870 30246 14922
rect 30298 14870 30350 14922
rect 30402 14870 30454 14922
rect 49514 14870 49566 14922
rect 49618 14870 49670 14922
rect 49722 14870 49774 14922
rect 68834 14870 68886 14922
rect 68938 14870 68990 14922
rect 69042 14870 69094 14922
rect 34862 14590 34914 14642
rect 33854 14366 33906 14418
rect 37326 14366 37378 14418
rect 38110 14366 38162 14418
rect 37102 14254 37154 14306
rect 37214 14254 37266 14306
rect 37998 14254 38050 14306
rect 38558 14254 38610 14306
rect 20534 14086 20586 14138
rect 20638 14086 20690 14138
rect 20742 14086 20794 14138
rect 39854 14086 39906 14138
rect 39958 14086 40010 14138
rect 40062 14086 40114 14138
rect 59174 14086 59226 14138
rect 59278 14086 59330 14138
rect 59382 14086 59434 14138
rect 78494 14086 78546 14138
rect 78598 14086 78650 14138
rect 78702 14086 78754 14138
rect 34526 13806 34578 13858
rect 35310 13806 35362 13858
rect 39902 13806 39954 13858
rect 13246 13582 13298 13634
rect 32174 13582 32226 13634
rect 32510 13582 32562 13634
rect 33182 13582 33234 13634
rect 33742 13582 33794 13634
rect 34638 13582 34690 13634
rect 36318 13582 36370 13634
rect 38894 13582 38946 13634
rect 41134 13582 41186 13634
rect 31950 13470 32002 13522
rect 32510 13470 32562 13522
rect 34750 13470 34802 13522
rect 10874 13302 10926 13354
rect 10978 13302 11030 13354
rect 11082 13302 11134 13354
rect 30194 13302 30246 13354
rect 30298 13302 30350 13354
rect 30402 13302 30454 13354
rect 49514 13302 49566 13354
rect 49618 13302 49670 13354
rect 49722 13302 49774 13354
rect 68834 13302 68886 13354
rect 68938 13302 68990 13354
rect 69042 13302 69094 13354
rect 12910 13022 12962 13074
rect 33518 13022 33570 13074
rect 35646 13022 35698 13074
rect 37774 13022 37826 13074
rect 39902 13022 39954 13074
rect 46174 13022 46226 13074
rect 10110 12910 10162 12962
rect 13582 12910 13634 12962
rect 19406 12910 19458 12962
rect 31950 12910 32002 12962
rect 36318 12910 36370 12962
rect 36990 12910 37042 12962
rect 10782 12798 10834 12850
rect 41246 12798 41298 12850
rect 41358 12798 41410 12850
rect 47518 12798 47570 12850
rect 13806 12686 13858 12738
rect 19630 12686 19682 12738
rect 20862 12686 20914 12738
rect 21758 12686 21810 12738
rect 22878 12686 22930 12738
rect 23662 12686 23714 12738
rect 24110 12686 24162 12738
rect 24446 12686 24498 12738
rect 25006 12686 25058 12738
rect 25342 12686 25394 12738
rect 25902 12686 25954 12738
rect 26686 12686 26738 12738
rect 27134 12686 27186 12738
rect 27582 12686 27634 12738
rect 30494 12686 30546 12738
rect 31054 12686 31106 12738
rect 31726 12686 31778 12738
rect 32510 12686 32562 12738
rect 33294 12686 33346 12738
rect 40462 12686 40514 12738
rect 40798 12686 40850 12738
rect 41582 12686 41634 12738
rect 42030 12686 42082 12738
rect 42478 12686 42530 12738
rect 42814 12686 42866 12738
rect 45166 12686 45218 12738
rect 45614 12686 45666 12738
rect 48078 12686 48130 12738
rect 48638 12686 48690 12738
rect 20534 12518 20586 12570
rect 20638 12518 20690 12570
rect 20742 12518 20794 12570
rect 39854 12518 39906 12570
rect 39958 12518 40010 12570
rect 40062 12518 40114 12570
rect 59174 12518 59226 12570
rect 59278 12518 59330 12570
rect 59382 12518 59434 12570
rect 78494 12518 78546 12570
rect 78598 12518 78650 12570
rect 78702 12518 78754 12570
rect 11230 12350 11282 12402
rect 22542 12350 22594 12402
rect 25454 12350 25506 12402
rect 27358 12350 27410 12402
rect 33406 12350 33458 12402
rect 40238 12350 40290 12402
rect 12910 12238 12962 12290
rect 14366 12238 14418 12290
rect 20302 12238 20354 12290
rect 23550 12238 23602 12290
rect 29374 12238 29426 12290
rect 31838 12238 31890 12290
rect 32286 12238 32338 12290
rect 32510 12238 32562 12290
rect 44046 12238 44098 12290
rect 45614 12238 45666 12290
rect 48750 12238 48802 12290
rect 49310 12238 49362 12290
rect 11566 12126 11618 12178
rect 12014 12126 12066 12178
rect 13134 12126 13186 12178
rect 13694 12126 13746 12178
rect 17502 12126 17554 12178
rect 20974 12126 21026 12178
rect 23662 12126 23714 12178
rect 24222 12126 24274 12178
rect 33182 12126 33234 12178
rect 37662 12126 37714 12178
rect 39902 12126 39954 12178
rect 40350 12126 40402 12178
rect 44718 12126 44770 12178
rect 16494 12014 16546 12066
rect 18174 12014 18226 12066
rect 21534 12014 21586 12066
rect 22206 12014 22258 12066
rect 23102 12014 23154 12066
rect 25790 12014 25842 12066
rect 26238 12014 26290 12066
rect 26686 12014 26738 12066
rect 27918 12014 27970 12066
rect 28366 12014 28418 12066
rect 28814 12014 28866 12066
rect 30606 12014 30658 12066
rect 31390 12014 31442 12066
rect 32398 12014 32450 12066
rect 35310 12014 35362 12066
rect 40910 12014 40962 12066
rect 41246 12014 41298 12066
rect 41806 12014 41858 12066
rect 47742 12014 47794 12066
rect 49870 12014 49922 12066
rect 50318 12014 50370 12066
rect 50878 12014 50930 12066
rect 12350 11902 12402 11954
rect 24558 11902 24610 11954
rect 31390 11902 31442 11954
rect 31838 11902 31890 11954
rect 33518 11902 33570 11954
rect 39566 11902 39618 11954
rect 39902 11902 39954 11954
rect 10874 11734 10926 11786
rect 10978 11734 11030 11786
rect 11082 11734 11134 11786
rect 30194 11734 30246 11786
rect 30298 11734 30350 11786
rect 30402 11734 30454 11786
rect 49514 11734 49566 11786
rect 49618 11734 49670 11786
rect 49722 11734 49774 11786
rect 68834 11734 68886 11786
rect 68938 11734 68990 11786
rect 69042 11734 69094 11786
rect 14142 11566 14194 11618
rect 19518 11566 19570 11618
rect 69022 11566 69074 11618
rect 70478 11566 70530 11618
rect 23438 11454 23490 11506
rect 28254 11454 28306 11506
rect 29374 11454 29426 11506
rect 33518 11454 33570 11506
rect 38110 11454 38162 11506
rect 43262 11454 43314 11506
rect 46174 11454 46226 11506
rect 49646 11454 49698 11506
rect 50094 11454 50146 11506
rect 50542 11454 50594 11506
rect 14478 11342 14530 11394
rect 19854 11342 19906 11394
rect 20638 11342 20690 11394
rect 26238 11342 26290 11394
rect 32846 11342 32898 11394
rect 36318 11342 36370 11394
rect 36990 11342 37042 11394
rect 37214 11342 37266 11394
rect 37886 11342 37938 11394
rect 41694 11342 41746 11394
rect 42366 11342 42418 11394
rect 43150 11342 43202 11394
rect 43486 11342 43538 11394
rect 44382 11342 44434 11394
rect 49198 11342 49250 11394
rect 69022 11342 69074 11394
rect 14702 11230 14754 11282
rect 15150 11230 15202 11282
rect 20414 11230 20466 11282
rect 22206 11230 22258 11282
rect 25566 11230 25618 11282
rect 29486 11230 29538 11282
rect 32174 11230 32226 11282
rect 35646 11230 35698 11282
rect 38222 11230 38274 11282
rect 41022 11230 41074 11282
rect 42814 11230 42866 11282
rect 43710 11230 43762 11282
rect 43934 11230 43986 11282
rect 44830 11230 44882 11282
rect 48414 11230 48466 11282
rect 51550 11230 51602 11282
rect 12238 11118 12290 11170
rect 13582 11118 13634 11170
rect 15822 11118 15874 11170
rect 17726 11118 17778 11170
rect 18286 11118 18338 11170
rect 18846 11118 18898 11170
rect 21422 11118 21474 11170
rect 21870 11118 21922 11170
rect 22766 11118 22818 11170
rect 23102 11118 23154 11170
rect 26798 11118 26850 11170
rect 27246 11118 27298 11170
rect 27806 11118 27858 11170
rect 28590 11118 28642 11170
rect 29262 11118 29314 11170
rect 29934 11118 29986 11170
rect 37550 11118 37602 11170
rect 38782 11118 38834 11170
rect 42142 11118 42194 11170
rect 44158 11118 44210 11170
rect 44942 11118 44994 11170
rect 45166 11118 45218 11170
rect 45390 11118 45442 11170
rect 68574 11118 68626 11170
rect 69470 11118 69522 11170
rect 69918 11118 69970 11170
rect 70366 11118 70418 11170
rect 70702 11118 70754 11170
rect 71262 11118 71314 11170
rect 71710 11118 71762 11170
rect 72158 11118 72210 11170
rect 72494 11118 72546 11170
rect 72942 11118 72994 11170
rect 73838 11118 73890 11170
rect 20534 10950 20586 11002
rect 20638 10950 20690 11002
rect 20742 10950 20794 11002
rect 39854 10950 39906 11002
rect 39958 10950 40010 11002
rect 40062 10950 40114 11002
rect 59174 10950 59226 11002
rect 59278 10950 59330 11002
rect 59382 10950 59434 11002
rect 78494 10950 78546 11002
rect 78598 10950 78650 11002
rect 78702 10950 78754 11002
rect 16942 10782 16994 10834
rect 17950 10782 18002 10834
rect 25566 10782 25618 10834
rect 33406 10782 33458 10834
rect 33854 10782 33906 10834
rect 47854 10782 47906 10834
rect 76974 10782 77026 10834
rect 21086 10670 21138 10722
rect 25230 10670 25282 10722
rect 25902 10670 25954 10722
rect 30158 10670 30210 10722
rect 31726 10670 31778 10722
rect 36094 10670 36146 10722
rect 38670 10670 38722 10722
rect 39342 10670 39394 10722
rect 39790 10670 39842 10722
rect 48190 10670 48242 10722
rect 50766 10670 50818 10722
rect 51550 10670 51602 10722
rect 51998 10670 52050 10722
rect 70254 10670 70306 10722
rect 70702 10670 70754 10722
rect 71374 10670 71426 10722
rect 72270 10670 72322 10722
rect 77870 10670 77922 10722
rect 9550 10558 9602 10610
rect 19966 10558 20018 10610
rect 30830 10558 30882 10610
rect 31166 10558 31218 10610
rect 31390 10558 31442 10610
rect 31950 10558 32002 10610
rect 33070 10558 33122 10610
rect 40126 10558 40178 10610
rect 40350 10558 40402 10610
rect 40910 10558 40962 10610
rect 46734 10558 46786 10610
rect 46958 10558 47010 10610
rect 49198 10558 49250 10610
rect 70926 10558 70978 10610
rect 72830 10558 72882 10610
rect 78206 10558 78258 10610
rect 10334 10446 10386 10498
rect 12462 10446 12514 10498
rect 12910 10446 12962 10498
rect 13358 10446 13410 10498
rect 14030 10446 14082 10498
rect 15038 10446 15090 10498
rect 16382 10446 16434 10498
rect 17502 10446 17554 10498
rect 18510 10446 18562 10498
rect 26798 10446 26850 10498
rect 27246 10446 27298 10498
rect 27694 10446 27746 10498
rect 28030 10446 28082 10498
rect 34414 10446 34466 10498
rect 34750 10446 34802 10498
rect 36654 10446 36706 10498
rect 37214 10446 37266 10498
rect 37550 10446 37602 10498
rect 40238 10446 40290 10498
rect 43710 10446 43762 10498
rect 46510 10446 46562 10498
rect 48750 10446 48802 10498
rect 49758 10446 49810 10498
rect 52558 10446 52610 10498
rect 53006 10446 53058 10498
rect 53566 10446 53618 10498
rect 54014 10446 54066 10498
rect 63534 10446 63586 10498
rect 63982 10446 64034 10498
rect 64542 10446 64594 10498
rect 65102 10446 65154 10498
rect 65438 10446 65490 10498
rect 66222 10446 66274 10498
rect 67006 10446 67058 10498
rect 67678 10446 67730 10498
rect 68126 10446 68178 10498
rect 68798 10446 68850 10498
rect 69134 10446 69186 10498
rect 69806 10446 69858 10498
rect 73278 10446 73330 10498
rect 73838 10446 73890 10498
rect 74174 10446 74226 10498
rect 74622 10446 74674 10498
rect 75182 10446 75234 10498
rect 75966 10446 76018 10498
rect 76638 10446 76690 10498
rect 77646 10446 77698 10498
rect 32286 10334 32338 10386
rect 39454 10334 39506 10386
rect 52670 10334 52722 10386
rect 53566 10334 53618 10386
rect 74174 10334 74226 10386
rect 74734 10334 74786 10386
rect 10874 10166 10926 10218
rect 10978 10166 11030 10218
rect 11082 10166 11134 10218
rect 30194 10166 30246 10218
rect 30298 10166 30350 10218
rect 30402 10166 30454 10218
rect 49514 10166 49566 10218
rect 49618 10166 49670 10218
rect 49722 10166 49774 10218
rect 68834 10166 68886 10218
rect 68938 10166 68990 10218
rect 69042 10166 69094 10218
rect 36430 9998 36482 10050
rect 70142 9998 70194 10050
rect 70478 9998 70530 10050
rect 9438 9886 9490 9938
rect 18286 9886 18338 9938
rect 18734 9886 18786 9938
rect 20302 9886 20354 9938
rect 22094 9886 22146 9938
rect 24222 9886 24274 9938
rect 27582 9886 27634 9938
rect 28702 9886 28754 9938
rect 29934 9886 29986 9938
rect 32062 9886 32114 9938
rect 32622 9886 32674 9938
rect 34750 9886 34802 9938
rect 35870 9886 35922 9938
rect 37438 9886 37490 9938
rect 37998 9886 38050 9938
rect 38894 9886 38946 9938
rect 40798 9886 40850 9938
rect 41470 9886 41522 9938
rect 45166 9886 45218 9938
rect 45838 9886 45890 9938
rect 47070 9886 47122 9938
rect 49310 9886 49362 9938
rect 54574 9886 54626 9938
rect 11566 9774 11618 9826
rect 12126 9774 12178 9826
rect 15374 9774 15426 9826
rect 21422 9774 21474 9826
rect 28142 9774 28194 9826
rect 29262 9774 29314 9826
rect 35534 9774 35586 9826
rect 36094 9774 36146 9826
rect 36990 9774 37042 9826
rect 45726 9774 45778 9826
rect 49982 9774 50034 9826
rect 63086 9774 63138 9826
rect 71262 9774 71314 9826
rect 72606 9774 72658 9826
rect 78094 9774 78146 9826
rect 10222 9662 10274 9714
rect 10558 9662 10610 9714
rect 11230 9662 11282 9714
rect 12350 9662 12402 9714
rect 14366 9662 14418 9714
rect 14702 9662 14754 9714
rect 16158 9662 16210 9714
rect 26462 9662 26514 9714
rect 39902 9662 39954 9714
rect 42030 9662 42082 9714
rect 46622 9662 46674 9714
rect 50766 9662 50818 9714
rect 65662 9662 65714 9714
rect 66782 9662 66834 9714
rect 67454 9662 67506 9714
rect 67790 9662 67842 9714
rect 71038 9662 71090 9714
rect 72046 9662 72098 9714
rect 73054 9662 73106 9714
rect 74062 9662 74114 9714
rect 76862 9662 76914 9714
rect 77198 9662 77250 9714
rect 77870 9662 77922 9714
rect 9998 9550 10050 9602
rect 12910 9550 12962 9602
rect 13582 9550 13634 9602
rect 14142 9550 14194 9602
rect 19182 9550 19234 9602
rect 19854 9550 19906 9602
rect 20862 9550 20914 9602
rect 24894 9550 24946 9602
rect 25342 9550 25394 9602
rect 25790 9550 25842 9602
rect 38670 9550 38722 9602
rect 44382 9550 44434 9602
rect 50542 9550 50594 9602
rect 50654 9550 50706 9602
rect 51102 9550 51154 9602
rect 51550 9550 51602 9602
rect 51998 9550 52050 9602
rect 52670 9550 52722 9602
rect 53118 9550 53170 9602
rect 53566 9550 53618 9602
rect 54014 9550 54066 9602
rect 55022 9550 55074 9602
rect 59950 9550 60002 9602
rect 60846 9550 60898 9602
rect 61294 9550 61346 9602
rect 62526 9550 62578 9602
rect 63422 9550 63474 9602
rect 64206 9550 64258 9602
rect 64766 9550 64818 9602
rect 65326 9550 65378 9602
rect 66222 9550 66274 9602
rect 67006 9550 67058 9602
rect 68574 9550 68626 9602
rect 69022 9550 69074 9602
rect 69470 9550 69522 9602
rect 71710 9550 71762 9602
rect 72382 9550 72434 9602
rect 73390 9550 73442 9602
rect 73726 9550 73778 9602
rect 74398 9550 74450 9602
rect 74958 9550 75010 9602
rect 75406 9550 75458 9602
rect 76190 9550 76242 9602
rect 20534 9382 20586 9434
rect 20638 9382 20690 9434
rect 20742 9382 20794 9434
rect 39854 9382 39906 9434
rect 39958 9382 40010 9434
rect 40062 9382 40114 9434
rect 59174 9382 59226 9434
rect 59278 9382 59330 9434
rect 59382 9382 59434 9434
rect 78494 9382 78546 9434
rect 78598 9382 78650 9434
rect 78702 9382 78754 9434
rect 17502 9214 17554 9266
rect 18846 9214 18898 9266
rect 22542 9214 22594 9266
rect 26462 9214 26514 9266
rect 30942 9214 30994 9266
rect 34190 9214 34242 9266
rect 34638 9214 34690 9266
rect 41694 9214 41746 9266
rect 47854 9214 47906 9266
rect 58942 9214 58994 9266
rect 59390 9214 59442 9266
rect 60174 9214 60226 9266
rect 61182 9214 61234 9266
rect 63534 9214 63586 9266
rect 64654 9214 64706 9266
rect 65326 9214 65378 9266
rect 66782 9214 66834 9266
rect 69246 9214 69298 9266
rect 75854 9214 75906 9266
rect 9998 9102 10050 9154
rect 10334 9102 10386 9154
rect 12014 9102 12066 9154
rect 13582 9102 13634 9154
rect 17726 9102 17778 9154
rect 23438 9102 23490 9154
rect 24110 9102 24162 9154
rect 24558 9102 24610 9154
rect 25678 9102 25730 9154
rect 26350 9102 26402 9154
rect 30494 9102 30546 9154
rect 31390 9102 31442 9154
rect 33406 9102 33458 9154
rect 35982 9102 36034 9154
rect 37214 9102 37266 9154
rect 40238 9102 40290 9154
rect 41358 9102 41410 9154
rect 47182 9102 47234 9154
rect 47742 9102 47794 9154
rect 48862 9102 48914 9154
rect 49422 9102 49474 9154
rect 55470 9102 55522 9154
rect 61966 9102 62018 9154
rect 62862 9102 62914 9154
rect 65998 9102 66050 9154
rect 67454 9102 67506 9154
rect 67902 9102 67954 9154
rect 68574 9102 68626 9154
rect 69806 9102 69858 9154
rect 71262 9102 71314 9154
rect 73278 9102 73330 9154
rect 74174 9102 74226 9154
rect 76862 9102 76914 9154
rect 9774 8990 9826 9042
rect 10670 8990 10722 9042
rect 11118 8990 11170 9042
rect 11454 8990 11506 9042
rect 12126 8990 12178 9042
rect 13358 8990 13410 9042
rect 16830 8990 16882 9042
rect 17390 8990 17442 9042
rect 17838 8990 17890 9042
rect 21870 8990 21922 9042
rect 23662 8990 23714 9042
rect 27022 8990 27074 9042
rect 30718 8990 30770 9042
rect 31502 8990 31554 9042
rect 32510 8990 32562 9042
rect 33070 8990 33122 9042
rect 33518 8990 33570 9042
rect 37102 8990 37154 9042
rect 40910 8990 40962 9042
rect 41022 8990 41074 9042
rect 41582 8990 41634 9042
rect 41806 8990 41858 9042
rect 45390 8990 45442 9042
rect 53006 8990 53058 9042
rect 53902 8990 53954 9042
rect 62526 8990 62578 9042
rect 63198 8990 63250 9042
rect 63870 8990 63922 9042
rect 64878 8990 64930 9042
rect 65662 8990 65714 9042
rect 66222 8990 66274 9042
rect 67118 8990 67170 9042
rect 68238 8990 68290 9042
rect 68798 8990 68850 9042
rect 69582 8990 69634 9042
rect 8542 8878 8594 8930
rect 9102 8878 9154 8930
rect 13022 8878 13074 8930
rect 13918 8878 13970 8930
rect 16046 8878 16098 8930
rect 19070 8878 19122 8930
rect 21198 8878 21250 8930
rect 27694 8878 27746 8930
rect 29822 8878 29874 8930
rect 33182 8878 33234 8930
rect 34974 8878 35026 8930
rect 37550 8878 37602 8930
rect 37998 8878 38050 8930
rect 38558 8878 38610 8930
rect 39118 8878 39170 8930
rect 42590 8878 42642 8930
rect 44718 8878 44770 8930
rect 45838 8878 45890 8930
rect 48862 8878 48914 8930
rect 49086 8878 49138 8930
rect 50094 8878 50146 8930
rect 52222 8878 52274 8930
rect 53454 8878 53506 8930
rect 54350 8878 54402 8930
rect 56814 8878 56866 8930
rect 57150 8878 57202 8930
rect 60846 8878 60898 8930
rect 61742 8878 61794 8930
rect 22878 8766 22930 8818
rect 25566 8766 25618 8818
rect 25902 8766 25954 8818
rect 26574 8766 26626 8818
rect 77534 9102 77586 9154
rect 70478 8990 70530 9042
rect 71150 8990 71202 9042
rect 76190 8990 76242 9042
rect 77086 8990 77138 9042
rect 77758 8990 77810 9042
rect 72270 8878 72322 8930
rect 75518 8878 75570 8930
rect 47966 8766 48018 8818
rect 53230 8766 53282 8818
rect 53454 8766 53506 8818
rect 60510 8766 60562 8818
rect 61630 8766 61682 8818
rect 69806 8766 69858 8818
rect 70142 8766 70194 8818
rect 10874 8598 10926 8650
rect 10978 8598 11030 8650
rect 11082 8598 11134 8650
rect 30194 8598 30246 8650
rect 30298 8598 30350 8650
rect 30402 8598 30454 8650
rect 49514 8598 49566 8650
rect 49618 8598 49670 8650
rect 49722 8598 49774 8650
rect 68834 8598 68886 8650
rect 68938 8598 68990 8650
rect 69042 8598 69094 8650
rect 17838 8430 17890 8482
rect 43710 8430 43762 8482
rect 12014 8318 12066 8370
rect 14030 8318 14082 8370
rect 19406 8318 19458 8370
rect 20302 8318 20354 8370
rect 23886 8318 23938 8370
rect 25118 8318 25170 8370
rect 27246 8318 27298 8370
rect 35534 8318 35586 8370
rect 36430 8318 36482 8370
rect 37438 8318 37490 8370
rect 42030 8318 42082 8370
rect 45054 8318 45106 8370
rect 47966 8318 48018 8370
rect 48638 8318 48690 8370
rect 50766 8318 50818 8370
rect 51550 8318 51602 8370
rect 53006 8318 53058 8370
rect 53790 8318 53842 8370
rect 58382 8318 58434 8370
rect 62190 8318 62242 8370
rect 68350 8318 68402 8370
rect 70142 8318 70194 8370
rect 73166 8318 73218 8370
rect 73726 8318 73778 8370
rect 76190 8318 76242 8370
rect 9102 8206 9154 8258
rect 9886 8206 9938 8258
rect 12462 8206 12514 8258
rect 15150 8206 15202 8258
rect 15822 8206 15874 8258
rect 16382 8206 16434 8258
rect 16942 8206 16994 8258
rect 17502 8206 17554 8258
rect 17838 8206 17890 8258
rect 19182 8206 19234 8258
rect 19854 8206 19906 8258
rect 20190 8206 20242 8258
rect 20526 8206 20578 8258
rect 21646 8206 21698 8258
rect 23550 8206 23602 8258
rect 24334 8206 24386 8258
rect 27918 8206 27970 8258
rect 34414 8206 34466 8258
rect 35870 8206 35922 8258
rect 37774 8206 37826 8258
rect 39902 8206 39954 8258
rect 44046 8206 44098 8258
rect 44382 8206 44434 8258
rect 8094 8094 8146 8146
rect 13806 8094 13858 8146
rect 15374 8094 15426 8146
rect 15934 8094 15986 8146
rect 16606 8094 16658 8146
rect 17166 8094 17218 8146
rect 18510 8094 18562 8146
rect 19518 8094 19570 8146
rect 21310 8094 21362 8146
rect 6302 7982 6354 8034
rect 7422 7982 7474 8034
rect 7870 7982 7922 8034
rect 8430 7982 8482 8034
rect 12686 7982 12738 8034
rect 14590 7982 14642 8034
rect 16046 7982 16098 8034
rect 16718 7982 16770 8034
rect 18174 7982 18226 8034
rect 22094 7982 22146 8034
rect 22542 8038 22594 8090
rect 28030 8094 28082 8146
rect 28142 8094 28194 8146
rect 30270 8094 30322 8146
rect 34862 8094 34914 8146
rect 34974 8094 35026 8146
rect 35086 8094 35138 8146
rect 37214 8094 37266 8146
rect 37326 8094 37378 8146
rect 38894 8094 38946 8146
rect 44830 8150 44882 8202
rect 50430 8206 50482 8258
rect 51886 8206 51938 8258
rect 58494 8206 58546 8258
rect 61742 8206 61794 8258
rect 62526 8206 62578 8258
rect 63534 8206 63586 8258
rect 63646 8206 63698 8258
rect 63870 8206 63922 8258
rect 64430 8206 64482 8258
rect 64990 8206 65042 8258
rect 65550 8206 65602 8258
rect 66894 8206 66946 8258
rect 67566 8206 67618 8258
rect 40350 8094 40402 8146
rect 43374 8094 43426 8146
rect 45278 8094 45330 8146
rect 45838 8094 45890 8146
rect 49646 8094 49698 8146
rect 51998 8094 52050 8146
rect 52670 8094 52722 8146
rect 52894 8094 52946 8146
rect 55022 8094 55074 8146
rect 57934 8094 57986 8146
rect 61070 8094 61122 8146
rect 65998 8094 66050 8146
rect 66334 8094 66386 8146
rect 66670 8094 66722 8146
rect 69358 8094 69410 8146
rect 71262 8094 71314 8146
rect 72046 8094 72098 8146
rect 74734 8094 74786 8146
rect 77534 8094 77586 8146
rect 22990 7982 23042 8034
rect 28590 7982 28642 8034
rect 41022 7982 41074 8034
rect 43822 7982 43874 8034
rect 45054 7982 45106 8034
rect 50654 7982 50706 8034
rect 55470 7982 55522 8034
rect 55918 7982 55970 8034
rect 56366 7982 56418 8034
rect 56814 7982 56866 8034
rect 57262 7982 57314 8034
rect 59054 7982 59106 8034
rect 59502 7982 59554 8034
rect 60622 7982 60674 8034
rect 61518 7982 61570 8034
rect 62302 7982 62354 8034
rect 63310 7982 63362 8034
rect 63422 7982 63474 8034
rect 65326 7982 65378 8034
rect 67342 7982 67394 8034
rect 75518 7982 75570 8034
rect 77982 7982 78034 8034
rect 20534 7814 20586 7866
rect 20638 7814 20690 7866
rect 20742 7814 20794 7866
rect 39854 7814 39906 7866
rect 39958 7814 40010 7866
rect 40062 7814 40114 7866
rect 59174 7814 59226 7866
rect 59278 7814 59330 7866
rect 59382 7814 59434 7866
rect 78494 7814 78546 7866
rect 78598 7814 78650 7866
rect 78702 7814 78754 7866
rect 7758 7646 7810 7698
rect 9998 7646 10050 7698
rect 10670 7646 10722 7698
rect 17726 7646 17778 7698
rect 24670 7646 24722 7698
rect 26798 7646 26850 7698
rect 29262 7646 29314 7698
rect 29822 7646 29874 7698
rect 30158 7646 30210 7698
rect 30606 7646 30658 7698
rect 38446 7646 38498 7698
rect 38558 7646 38610 7698
rect 38670 7646 38722 7698
rect 41134 7646 41186 7698
rect 41582 7646 41634 7698
rect 43822 7646 43874 7698
rect 44270 7646 44322 7698
rect 47854 7646 47906 7698
rect 48078 7646 48130 7698
rect 48974 7646 49026 7698
rect 53902 7646 53954 7698
rect 54350 7646 54402 7698
rect 54798 7646 54850 7698
rect 55470 7646 55522 7698
rect 56590 7646 56642 7698
rect 58606 7646 58658 7698
rect 66670 7646 66722 7698
rect 6078 7534 6130 7586
rect 7310 7534 7362 7586
rect 8766 7534 8818 7586
rect 23662 7534 23714 7586
rect 25342 7534 25394 7586
rect 25902 7534 25954 7586
rect 26350 7534 26402 7586
rect 27246 7534 27298 7586
rect 31950 7534 32002 7586
rect 33518 7534 33570 7586
rect 35758 7534 35810 7586
rect 36654 7534 36706 7586
rect 42926 7534 42978 7586
rect 45726 7534 45778 7586
rect 47182 7534 47234 7586
rect 48750 7534 48802 7586
rect 52334 7534 52386 7586
rect 53454 7534 53506 7586
rect 54462 7534 54514 7586
rect 55806 7534 55858 7586
rect 56926 7534 56978 7586
rect 57262 7534 57314 7586
rect 58382 7534 58434 7586
rect 59278 7534 59330 7586
rect 59726 7534 59778 7586
rect 60174 7534 60226 7586
rect 70814 7590 70866 7642
rect 77086 7646 77138 7698
rect 60958 7534 61010 7586
rect 62862 7534 62914 7586
rect 65326 7534 65378 7586
rect 65886 7534 65938 7586
rect 67342 7534 67394 7586
rect 70030 7534 70082 7586
rect 71486 7534 71538 7586
rect 72382 7534 72434 7586
rect 74398 7534 74450 7586
rect 77758 7534 77810 7586
rect 5854 7422 5906 7474
rect 6974 7422 7026 7474
rect 8094 7422 8146 7474
rect 8878 7422 8930 7474
rect 9662 7422 9714 7474
rect 10446 7422 10498 7474
rect 13134 7422 13186 7474
rect 16494 7422 16546 7474
rect 21758 7422 21810 7474
rect 24110 7422 24162 7474
rect 25678 7422 25730 7474
rect 26574 7422 26626 7474
rect 34078 7422 34130 7474
rect 34414 7422 34466 7474
rect 36206 7422 36258 7474
rect 36430 7422 36482 7474
rect 39006 7422 39058 7474
rect 39454 7422 39506 7474
rect 39902 7422 39954 7474
rect 46622 7422 46674 7474
rect 46734 7422 46786 7474
rect 46846 7422 46898 7474
rect 47518 7422 47570 7474
rect 48190 7422 48242 7474
rect 49086 7422 49138 7474
rect 49310 7422 49362 7474
rect 53006 7422 53058 7474
rect 55134 7422 55186 7474
rect 57486 7422 57538 7474
rect 57710 7422 57762 7474
rect 64542 7422 64594 7474
rect 66334 7422 66386 7474
rect 66894 7422 66946 7474
rect 71150 7422 71202 7474
rect 77310 7422 77362 7474
rect 77982 7422 78034 7474
rect 5518 7310 5570 7362
rect 6526 7310 6578 7362
rect 18846 7310 18898 7362
rect 26798 7310 26850 7362
rect 28366 7310 28418 7362
rect 30942 7310 30994 7362
rect 33182 7310 33234 7362
rect 38222 7310 38274 7362
rect 40350 7310 40402 7362
rect 41918 7310 41970 7362
rect 44718 7310 44770 7362
rect 47854 7310 47906 7362
rect 50094 7310 50146 7362
rect 58494 7310 58546 7362
rect 59166 7310 59218 7362
rect 61518 7310 61570 7362
rect 63534 7310 63586 7362
rect 64878 7310 64930 7362
rect 68462 7310 68514 7362
rect 69022 7310 69074 7362
rect 73726 7310 73778 7362
rect 76526 7310 76578 7362
rect 11230 7198 11282 7250
rect 14142 7198 14194 7250
rect 26014 7198 26066 7250
rect 59054 7198 59106 7250
rect 63422 7198 63474 7250
rect 63758 7198 63810 7250
rect 63870 7198 63922 7250
rect 10874 7030 10926 7082
rect 10978 7030 11030 7082
rect 11082 7030 11134 7082
rect 30194 7030 30246 7082
rect 30298 7030 30350 7082
rect 30402 7030 30454 7082
rect 49514 7030 49566 7082
rect 49618 7030 49670 7082
rect 49722 7030 49774 7082
rect 68834 7030 68886 7082
rect 68938 7030 68990 7082
rect 69042 7030 69094 7082
rect 14366 6862 14418 6914
rect 20078 6862 20130 6914
rect 26462 6862 26514 6914
rect 9886 6750 9938 6802
rect 16046 6750 16098 6802
rect 20414 6750 20466 6802
rect 5742 6638 5794 6690
rect 6302 6638 6354 6690
rect 7086 6638 7138 6690
rect 7758 6638 7810 6690
rect 12462 6638 12514 6690
rect 13918 6638 13970 6690
rect 14702 6638 14754 6690
rect 15262 6638 15314 6690
rect 15710 6638 15762 6690
rect 18846 6638 18898 6690
rect 19518 6638 19570 6690
rect 21198 6638 21250 6690
rect 21646 6638 21698 6690
rect 21758 6638 21810 6690
rect 23550 6638 23602 6690
rect 24558 6638 24610 6690
rect 25118 6638 25170 6690
rect 25678 6638 25730 6690
rect 4734 6526 4786 6578
rect 5070 6526 5122 6578
rect 6638 6526 6690 6578
rect 11342 6526 11394 6578
rect 13694 6526 13746 6578
rect 18174 6526 18226 6578
rect 19294 6526 19346 6578
rect 22990 6526 23042 6578
rect 24782 6526 24834 6578
rect 25566 6526 25618 6578
rect 4510 6414 4562 6466
rect 5966 6414 6018 6466
rect 20302 6414 20354 6466
rect 21534 6414 21586 6466
rect 22654 6414 22706 6466
rect 23102 6414 23154 6466
rect 23326 6414 23378 6466
rect 40686 6862 40738 6914
rect 41358 6862 41410 6914
rect 42030 6862 42082 6914
rect 43150 6862 43202 6914
rect 45166 6862 45218 6914
rect 45502 6862 45554 6914
rect 26910 6750 26962 6802
rect 27134 6750 27186 6802
rect 29374 6750 29426 6802
rect 34078 6750 34130 6802
rect 40014 6750 40066 6802
rect 40910 6750 40962 6802
rect 45950 6750 46002 6802
rect 49198 6750 49250 6802
rect 29598 6638 29650 6690
rect 31166 6638 31218 6690
rect 36094 6638 36146 6690
rect 36990 6638 37042 6690
rect 37998 6638 38050 6690
rect 39118 6638 39170 6690
rect 39790 6638 39842 6690
rect 40238 6638 40290 6690
rect 40350 6638 40402 6690
rect 50318 6862 50370 6914
rect 52558 6862 52610 6914
rect 52782 6862 52834 6914
rect 55694 6862 55746 6914
rect 59614 6862 59666 6914
rect 75630 6862 75682 6914
rect 50206 6750 50258 6802
rect 51774 6750 51826 6802
rect 40462 6638 40514 6690
rect 41806 6638 41858 6690
rect 42254 6638 42306 6690
rect 42814 6638 42866 6690
rect 43710 6638 43762 6690
rect 44046 6638 44098 6690
rect 45614 6638 45666 6690
rect 50094 6638 50146 6690
rect 28142 6526 28194 6578
rect 29150 6526 29202 6578
rect 38222 6526 38274 6578
rect 38894 6526 38946 6578
rect 39566 6526 39618 6578
rect 41582 6526 41634 6578
rect 42478 6526 42530 6578
rect 52110 6750 52162 6802
rect 52894 6750 52946 6802
rect 58718 6750 58770 6802
rect 60734 6750 60786 6802
rect 61518 6750 61570 6802
rect 63422 6750 63474 6802
rect 65662 6750 65714 6802
rect 69806 6750 69858 6802
rect 72830 6750 72882 6802
rect 77646 6750 77698 6802
rect 50766 6638 50818 6690
rect 51102 6638 51154 6690
rect 51438 6638 51490 6690
rect 58942 6638 58994 6690
rect 63310 6638 63362 6690
rect 66558 6638 66610 6690
rect 67678 6638 67730 6690
rect 43038 6526 43090 6578
rect 47070 6526 47122 6578
rect 48078 6526 48130 6578
rect 50206 6526 50258 6578
rect 55358 6526 55410 6578
rect 58158 6526 58210 6578
rect 58606 6526 58658 6578
rect 59502 6526 59554 6578
rect 62862 6526 62914 6578
rect 63982 6526 64034 6578
rect 64542 6526 64594 6578
rect 66670 6526 66722 6578
rect 68574 6526 68626 6578
rect 70366 6526 70418 6578
rect 73502 6526 73554 6578
rect 76302 6526 76354 6578
rect 26462 6414 26514 6466
rect 26574 6414 26626 6466
rect 31950 6414 32002 6466
rect 38110 6414 38162 6466
rect 42030 6414 42082 6466
rect 44942 6414 44994 6466
rect 49870 6414 49922 6466
rect 50318 6414 50370 6466
rect 50990 6414 51042 6466
rect 51550 6414 51602 6466
rect 59726 6414 59778 6466
rect 59950 6414 60002 6466
rect 61070 6414 61122 6466
rect 63534 6414 63586 6466
rect 63758 6414 63810 6466
rect 67454 6414 67506 6466
rect 77982 6414 78034 6466
rect 20534 6246 20586 6298
rect 20638 6246 20690 6298
rect 20742 6246 20794 6298
rect 39854 6246 39906 6298
rect 39958 6246 40010 6298
rect 40062 6246 40114 6298
rect 59174 6246 59226 6298
rect 59278 6246 59330 6298
rect 59382 6246 59434 6298
rect 78494 6246 78546 6298
rect 78598 6246 78650 6298
rect 78702 6246 78754 6298
rect 9662 6078 9714 6130
rect 17614 6078 17666 6130
rect 18510 6078 18562 6130
rect 19518 6078 19570 6130
rect 24334 6078 24386 6130
rect 33854 6078 33906 6130
rect 40238 6078 40290 6130
rect 40910 6078 40962 6130
rect 41694 6078 41746 6130
rect 42926 6078 42978 6130
rect 43934 6078 43986 6130
rect 52334 6078 52386 6130
rect 53902 6078 53954 6130
rect 56702 6078 56754 6130
rect 77646 6078 77698 6130
rect 10334 5966 10386 6018
rect 10558 5966 10610 6018
rect 17726 5966 17778 6018
rect 18174 5966 18226 6018
rect 18846 5966 18898 6018
rect 21982 5966 22034 6018
rect 23214 5966 23266 6018
rect 25342 5966 25394 6018
rect 27470 5966 27522 6018
rect 27806 5966 27858 6018
rect 29374 5966 29426 6018
rect 33182 5966 33234 6018
rect 33294 5966 33346 6018
rect 33406 5966 33458 6018
rect 40014 5966 40066 6018
rect 40350 5966 40402 6018
rect 42254 5966 42306 6018
rect 43150 5966 43202 6018
rect 44382 5966 44434 6018
rect 46510 5966 46562 6018
rect 51326 5966 51378 6018
rect 54238 5966 54290 6018
rect 54574 5966 54626 6018
rect 55470 5966 55522 6018
rect 57262 5966 57314 6018
rect 58046 5966 58098 6018
rect 58718 5966 58770 6018
rect 61742 5966 61794 6018
rect 62750 5966 62802 6018
rect 64542 5966 64594 6018
rect 65102 5966 65154 6018
rect 67790 5966 67842 6018
rect 68350 5966 68402 6018
rect 71038 5966 71090 6018
rect 72382 5966 72434 6018
rect 75182 5966 75234 6018
rect 77870 5966 77922 6018
rect 5966 5854 6018 5906
rect 8990 5854 9042 5906
rect 9998 5854 10050 5906
rect 11790 5854 11842 5906
rect 16382 5854 16434 5906
rect 17390 5854 17442 5906
rect 19294 5854 19346 5906
rect 22766 5854 22818 5906
rect 23326 5854 23378 5906
rect 23438 5854 23490 5906
rect 24670 5854 24722 5906
rect 25678 5854 25730 5906
rect 25902 5854 25954 5906
rect 26574 5854 26626 5906
rect 27694 5854 27746 5906
rect 29934 5854 29986 5906
rect 36878 5854 36930 5906
rect 39342 5854 39394 5906
rect 41134 5854 41186 5906
rect 41806 5854 41858 5906
rect 15150 5742 15202 5794
rect 19854 5742 19906 5794
rect 5070 5630 5122 5682
rect 7982 5630 8034 5682
rect 12798 5630 12850 5682
rect 23886 5630 23938 5682
rect 27358 5630 27410 5682
rect 42142 5854 42194 5906
rect 42590 5854 42642 5906
rect 42814 5854 42866 5906
rect 43374 5854 43426 5906
rect 47294 5854 47346 5906
rect 47630 5854 47682 5906
rect 48862 5854 48914 5906
rect 53230 5854 53282 5906
rect 54798 5854 54850 5906
rect 55806 5854 55858 5906
rect 56030 5854 56082 5906
rect 58942 5854 58994 5906
rect 59502 5854 59554 5906
rect 63086 5854 63138 5906
rect 63758 5854 63810 5906
rect 71262 5854 71314 5906
rect 78094 5854 78146 5906
rect 28142 5742 28194 5794
rect 44830 5742 44882 5794
rect 45390 5742 45442 5794
rect 48190 5742 48242 5794
rect 49310 5742 49362 5794
rect 50206 5742 50258 5794
rect 51886 5742 51938 5794
rect 52782 5742 52834 5794
rect 55918 5742 55970 5794
rect 57598 5742 57650 5794
rect 59950 5742 60002 5794
rect 60174 5742 60226 5794
rect 60398 5742 60450 5794
rect 62414 5742 62466 5794
rect 62862 5742 62914 5794
rect 67342 5742 67394 5794
rect 70590 5742 70642 5794
rect 74510 5742 74562 5794
rect 30942 5630 30994 5682
rect 34526 5630 34578 5682
rect 37438 5630 37490 5682
rect 43822 5630 43874 5682
rect 44270 5630 44322 5682
rect 52110 5630 52162 5682
rect 52670 5630 52722 5682
rect 59390 5630 59442 5682
rect 10874 5462 10926 5514
rect 10978 5462 11030 5514
rect 11082 5462 11134 5514
rect 30194 5462 30246 5514
rect 30298 5462 30350 5514
rect 30402 5462 30454 5514
rect 49514 5462 49566 5514
rect 49618 5462 49670 5514
rect 49722 5462 49774 5514
rect 68834 5462 68886 5514
rect 68938 5462 68990 5514
rect 69042 5462 69094 5514
rect 6750 5294 6802 5346
rect 17278 5294 17330 5346
rect 21310 5294 21362 5346
rect 22766 5294 22818 5346
rect 25790 5294 25842 5346
rect 37774 5294 37826 5346
rect 45390 5294 45442 5346
rect 47182 5294 47234 5346
rect 47630 5294 47682 5346
rect 52670 5294 52722 5346
rect 56254 5294 56306 5346
rect 60398 5294 60450 5346
rect 61070 5294 61122 5346
rect 2494 5182 2546 5234
rect 3838 5182 3890 5234
rect 5966 5182 6018 5234
rect 6190 5182 6242 5234
rect 7086 5182 7138 5234
rect 9214 5182 9266 5234
rect 14478 5182 14530 5234
rect 16606 5182 16658 5234
rect 26910 5182 26962 5234
rect 27358 5182 27410 5234
rect 30494 5182 30546 5234
rect 32958 5182 33010 5234
rect 35198 5182 35250 5234
rect 37886 5182 37938 5234
rect 39454 5182 39506 5234
rect 42702 5182 42754 5234
rect 44046 5182 44098 5234
rect 46510 5182 46562 5234
rect 46846 5182 46898 5234
rect 52110 5182 52162 5234
rect 53230 5182 53282 5234
rect 53454 5182 53506 5234
rect 59726 5182 59778 5234
rect 60622 5182 60674 5234
rect 61518 5182 61570 5234
rect 66110 5182 66162 5234
rect 70590 5182 70642 5234
rect 71262 5182 71314 5234
rect 74062 5182 74114 5234
rect 76190 5182 76242 5234
rect 2942 5070 2994 5122
rect 3390 5070 3442 5122
rect 4622 5070 4674 5122
rect 5070 5070 5122 5122
rect 6414 5070 6466 5122
rect 9886 5070 9938 5122
rect 12574 5070 12626 5122
rect 13694 5070 13746 5122
rect 16942 5070 16994 5122
rect 19966 5070 20018 5122
rect 20750 5070 20802 5122
rect 21422 5070 21474 5122
rect 21646 5070 21698 5122
rect 21982 5070 22034 5122
rect 22318 5070 22370 5122
rect 23102 5070 23154 5122
rect 23438 5070 23490 5122
rect 24670 5070 24722 5122
rect 25006 5070 25058 5122
rect 25230 5070 25282 5122
rect 25342 5070 25394 5122
rect 29262 5070 29314 5122
rect 29822 5070 29874 5122
rect 30606 5070 30658 5122
rect 31390 5070 31442 5122
rect 35982 5070 36034 5122
rect 37214 5070 37266 5122
rect 38446 5070 38498 5122
rect 41358 5070 41410 5122
rect 42254 5070 42306 5122
rect 42926 5070 42978 5122
rect 44830 5070 44882 5122
rect 45054 5070 45106 5122
rect 45950 5070 46002 5122
rect 48302 5070 48354 5122
rect 48638 5070 48690 5122
rect 50318 5070 50370 5122
rect 53006 5070 53058 5122
rect 59390 5070 59442 5122
rect 59502 5070 59554 5122
rect 59950 5070 60002 5122
rect 61070 5070 61122 5122
rect 22206 4958 22258 5010
rect 23326 4958 23378 5010
rect 24334 4958 24386 5010
rect 28254 4958 28306 5010
rect 29150 4958 29202 5010
rect 43486 4958 43538 5010
rect 45614 4958 45666 5010
rect 47966 4958 48018 5010
rect 48974 4958 49026 5010
rect 51102 4958 51154 5010
rect 55918 4958 55970 5010
rect 58382 4958 58434 5010
rect 62638 4958 62690 5010
rect 65662 4958 65714 5010
rect 67230 4958 67282 5010
rect 68462 4958 68514 5010
rect 73166 4958 73218 5010
rect 74958 4958 75010 5010
rect 77534 4958 77586 5010
rect 2046 4846 2098 4898
rect 4286 4846 4338 4898
rect 11902 4846 11954 4898
rect 17166 4846 17218 4898
rect 17726 4846 17778 4898
rect 23886 4846 23938 4898
rect 26350 4846 26402 4898
rect 38782 4846 38834 4898
rect 42478 4846 42530 4898
rect 42702 4846 42754 4898
rect 43710 4846 43762 4898
rect 43934 4846 43986 4898
rect 44046 4846 44098 4898
rect 45838 4846 45890 4898
rect 47294 4846 47346 4898
rect 49422 4846 49474 4898
rect 49870 4846 49922 4898
rect 59726 4846 59778 4898
rect 63198 4846 63250 4898
rect 77982 4846 78034 4898
rect 20534 4678 20586 4730
rect 20638 4678 20690 4730
rect 20742 4678 20794 4730
rect 39854 4678 39906 4730
rect 39958 4678 40010 4730
rect 40062 4678 40114 4730
rect 59174 4678 59226 4730
rect 59278 4678 59330 4730
rect 59382 4678 59434 4730
rect 78494 4678 78546 4730
rect 78598 4678 78650 4730
rect 78702 4678 78754 4730
rect 2494 4510 2546 4562
rect 10670 4510 10722 4562
rect 17838 4510 17890 4562
rect 24222 4510 24274 4562
rect 27694 4510 27746 4562
rect 44158 4510 44210 4562
rect 44830 4510 44882 4562
rect 48638 4510 48690 4562
rect 51662 4510 51714 4562
rect 51774 4510 51826 4562
rect 52334 4510 52386 4562
rect 54350 4510 54402 4562
rect 72158 4510 72210 4562
rect 13022 4398 13074 4450
rect 17390 4398 17442 4450
rect 17614 4398 17666 4450
rect 18958 4398 19010 4450
rect 22206 4398 22258 4450
rect 22542 4398 22594 4450
rect 23326 4398 23378 4450
rect 23438 4398 23490 4450
rect 25902 4398 25954 4450
rect 26798 4398 26850 4450
rect 29150 4398 29202 4450
rect 33182 4398 33234 4450
rect 34526 4398 34578 4450
rect 47966 4398 48018 4450
rect 50990 4398 51042 4450
rect 52222 4398 52274 4450
rect 55470 4398 55522 4450
rect 55806 4398 55858 4450
rect 56814 4398 56866 4450
rect 57038 4398 57090 4450
rect 58606 4398 58658 4450
rect 61742 4398 61794 4450
rect 62526 4398 62578 4450
rect 64542 4398 64594 4450
rect 67678 4398 67730 4450
rect 71038 4398 71090 4450
rect 74286 4398 74338 4450
rect 75182 4398 75234 4450
rect 77870 4398 77922 4450
rect 78206 4398 78258 4450
rect 2270 4286 2322 4338
rect 5630 4286 5682 4338
rect 8990 4286 9042 4338
rect 9550 4286 9602 4338
rect 13694 4286 13746 4338
rect 16718 4286 16770 4338
rect 18062 4286 18114 4338
rect 18734 4286 18786 4338
rect 21534 4286 21586 4338
rect 23102 4286 23154 4338
rect 24558 4286 24610 4338
rect 26126 4286 26178 4338
rect 26350 4286 26402 4338
rect 26574 4286 26626 4338
rect 29934 4286 29986 4338
rect 33966 4286 34018 4338
rect 34862 4286 34914 4338
rect 40350 4286 40402 4338
rect 43038 4286 43090 4338
rect 43822 4286 43874 4338
rect 44046 4286 44098 4338
rect 44270 4286 44322 4338
rect 44382 4286 44434 4338
rect 45054 4286 45106 4338
rect 45390 4286 45442 4338
rect 52110 4286 52162 4338
rect 52782 4286 52834 4338
rect 53342 4286 53394 4338
rect 53902 4286 53954 4338
rect 54798 4286 54850 4338
rect 55246 4286 55298 4338
rect 1934 4174 1986 4226
rect 3278 4174 3330 4226
rect 4846 4174 4898 4226
rect 7870 4174 7922 4226
rect 10894 4174 10946 4226
rect 15710 4174 15762 4226
rect 25678 4174 25730 4226
rect 26686 4174 26738 4226
rect 27246 4174 27298 4226
rect 28142 4174 28194 4226
rect 32174 4174 32226 4226
rect 33630 4174 33682 4226
rect 36206 4174 36258 4226
rect 38334 4174 38386 4226
rect 44942 4174 44994 4226
rect 52558 4174 52610 4226
rect 56702 4174 56754 4226
rect 57598 4174 57650 4226
rect 63870 4174 63922 4226
rect 66670 4174 66722 4226
rect 69470 4174 69522 4226
rect 70254 4174 70306 4226
rect 77310 4174 77362 4226
rect 9774 4062 9826 4114
rect 10110 4062 10162 4114
rect 19518 4062 19570 4114
rect 23886 4062 23938 4114
rect 41134 4062 41186 4114
rect 45614 4062 45666 4114
rect 53566 4062 53618 4114
rect 55022 4062 55074 4114
rect 59278 4062 59330 4114
rect 10874 3894 10926 3946
rect 10978 3894 11030 3946
rect 11082 3894 11134 3946
rect 30194 3894 30246 3946
rect 30298 3894 30350 3946
rect 30402 3894 30454 3946
rect 49514 3894 49566 3946
rect 49618 3894 49670 3946
rect 49722 3894 49774 3946
rect 68834 3894 68886 3946
rect 68938 3894 68990 3946
rect 69042 3894 69094 3946
rect 26126 3726 26178 3778
rect 27358 3726 27410 3778
rect 32510 3726 32562 3778
rect 43710 3726 43762 3778
rect 44606 3726 44658 3778
rect 59166 3726 59218 3778
rect 59390 3726 59442 3778
rect 65326 3726 65378 3778
rect 66334 3726 66386 3778
rect 4958 3614 5010 3666
rect 7758 3614 7810 3666
rect 11566 3614 11618 3666
rect 17614 3614 17666 3666
rect 21870 3614 21922 3666
rect 27582 3614 27634 3666
rect 31390 3614 31442 3666
rect 32398 3614 32450 3666
rect 34414 3614 34466 3666
rect 40686 3614 40738 3666
rect 44158 3614 44210 3666
rect 46510 3614 46562 3666
rect 48414 3614 48466 3666
rect 51886 3614 51938 3666
rect 52222 3614 52274 3666
rect 52558 3614 52610 3666
rect 52670 3614 52722 3666
rect 53230 3614 53282 3666
rect 53678 3614 53730 3666
rect 55470 3614 55522 3666
rect 55918 3614 55970 3666
rect 56926 3614 56978 3666
rect 57598 3614 57650 3666
rect 61070 3614 61122 3666
rect 72606 3614 72658 3666
rect 2270 3502 2322 3554
rect 3614 3502 3666 3554
rect 4062 3502 4114 3554
rect 4510 3502 4562 3554
rect 5630 3502 5682 3554
rect 8766 3502 8818 3554
rect 9326 3502 9378 3554
rect 12574 3502 12626 3554
rect 13134 3502 13186 3554
rect 16270 3502 16322 3554
rect 19742 3502 19794 3554
rect 20750 3502 20802 3554
rect 23662 3502 23714 3554
rect 25006 3502 25058 3554
rect 25566 3502 25618 3554
rect 25902 3502 25954 3554
rect 26350 3502 26402 3554
rect 26574 3502 26626 3554
rect 26910 3502 26962 3554
rect 27134 3502 27186 3554
rect 27806 3502 27858 3554
rect 28590 3502 28642 3554
rect 29038 3502 29090 3554
rect 35086 3502 35138 3554
rect 38782 3502 38834 3554
rect 42590 3502 42642 3554
rect 43934 3502 43986 3554
rect 45166 3502 45218 3554
rect 46174 3502 46226 3554
rect 46846 3502 46898 3554
rect 47406 3502 47458 3554
rect 50430 3502 50482 3554
rect 52894 3502 52946 3554
rect 53566 3502 53618 3554
rect 55358 3502 55410 3554
rect 55694 3502 55746 3554
rect 56254 3502 56306 3554
rect 57934 3502 57986 3554
rect 59614 3502 59666 3554
rect 59950 3502 60002 3554
rect 60174 3502 60226 3554
rect 60398 3502 60450 3554
rect 60622 3502 60674 3554
rect 60958 3502 61010 3554
rect 61182 3502 61234 3554
rect 61406 3502 61458 3554
rect 65774 3502 65826 3554
rect 69470 3502 69522 3554
rect 77086 3502 77138 3554
rect 78094 3502 78146 3554
rect 1934 3390 1986 3442
rect 2494 3390 2546 3442
rect 2830 3390 2882 3442
rect 14814 3390 14866 3442
rect 23998 3390 24050 3442
rect 25342 3390 25394 3442
rect 28366 3390 28418 3442
rect 32286 3390 32338 3442
rect 35982 3390 36034 3442
rect 36318 3390 36370 3442
rect 37662 3390 37714 3442
rect 46286 3390 46338 3442
rect 47742 3390 47794 3442
rect 49646 3390 49698 3442
rect 51214 3390 51266 3442
rect 51998 3390 52050 3442
rect 55022 3390 55074 3442
rect 56702 3390 56754 3442
rect 57374 3390 57426 3442
rect 60286 3390 60338 3442
rect 62862 3390 62914 3442
rect 65550 3390 65602 3442
rect 68462 3390 68514 3442
rect 70366 3390 70418 3442
rect 73502 3390 73554 3442
rect 73950 3390 74002 3442
rect 76078 3390 76130 3442
rect 76862 3390 76914 3442
rect 77870 3390 77922 3442
rect 3166 3278 3218 3330
rect 5854 3278 5906 3330
rect 9662 3278 9714 3330
rect 13470 3278 13522 3330
rect 17054 3278 17106 3330
rect 24670 3278 24722 3330
rect 26686 3278 26738 3330
rect 27918 3278 27970 3330
rect 40014 3278 40066 3330
rect 44718 3278 44770 3330
rect 44942 3278 44994 3330
rect 45726 3278 45778 3330
rect 45838 3278 45890 3330
rect 46958 3278 47010 3330
rect 50206 3278 50258 3330
rect 51550 3278 51602 3330
rect 54574 3278 54626 3330
rect 56030 3278 56082 3330
rect 56814 3278 56866 3330
rect 59502 3278 59554 3330
rect 61966 3278 62018 3330
rect 69246 3278 69298 3330
rect 73166 3278 73218 3330
rect 20534 3110 20586 3162
rect 20638 3110 20690 3162
rect 20742 3110 20794 3162
rect 39854 3110 39906 3162
rect 39958 3110 40010 3162
rect 40062 3110 40114 3162
rect 59174 3110 59226 3162
rect 59278 3110 59330 3162
rect 59382 3110 59434 3162
rect 78494 3110 78546 3162
rect 78598 3110 78650 3162
rect 78702 3110 78754 3162
rect 25454 2942 25506 2994
rect 29150 2942 29202 2994
rect 43374 2942 43426 2994
rect 47182 2942 47234 2994
rect 67454 2942 67506 2994
rect 68014 2942 68066 2994
rect 38894 2830 38946 2882
rect 40238 2830 40290 2882
rect 61406 2830 61458 2882
rect 67342 2830 67394 2882
rect 42926 2718 42978 2770
rect 45502 2718 45554 2770
rect 46286 2718 46338 2770
rect 62750 2718 62802 2770
rect 65998 2718 66050 2770
rect 68462 2718 68514 2770
rect 42814 2606 42866 2658
rect 43710 2606 43762 2658
rect 66110 2606 66162 2658
rect 70254 2606 70306 2658
rect 43262 2494 43314 2546
rect 44382 2494 44434 2546
rect 45390 2494 45442 2546
rect 54350 2494 54402 2546
rect 46062 2382 46114 2434
rect 54574 2382 54626 2434
rect 45726 2270 45778 2322
rect 50878 2270 50930 2322
rect 61630 1822 61682 1874
rect 64430 1822 64482 1874
rect 42366 926 42418 978
rect 45838 926 45890 978
<< metal2 >>
rect 10872 36876 11136 36886
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 10872 36810 11136 36820
rect 30192 36876 30456 36886
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30192 36810 30456 36820
rect 49512 36876 49776 36886
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49512 36810 49776 36820
rect 68832 36876 69096 36886
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 68832 36810 69096 36820
rect 20532 36092 20796 36102
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20532 36026 20796 36036
rect 39852 36092 40116 36102
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 39852 36026 40116 36036
rect 59172 36092 59436 36102
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59172 36026 59436 36036
rect 78492 36092 78756 36102
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78492 36026 78756 36036
rect 10872 35308 11136 35318
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 10872 35242 11136 35252
rect 30192 35308 30456 35318
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30192 35242 30456 35252
rect 49512 35308 49776 35318
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49512 35242 49776 35252
rect 68832 35308 69096 35318
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 68832 35242 69096 35252
rect 20532 34524 20796 34534
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20532 34458 20796 34468
rect 39852 34524 40116 34534
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 39852 34458 40116 34468
rect 59172 34524 59436 34534
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59172 34458 59436 34468
rect 78492 34524 78756 34534
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78492 34458 78756 34468
rect 10872 33740 11136 33750
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 10872 33674 11136 33684
rect 30192 33740 30456 33750
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30192 33674 30456 33684
rect 49512 33740 49776 33750
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49512 33674 49776 33684
rect 68832 33740 69096 33750
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 68832 33674 69096 33684
rect 20532 32956 20796 32966
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20532 32890 20796 32900
rect 39852 32956 40116 32966
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 39852 32890 40116 32900
rect 59172 32956 59436 32966
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59172 32890 59436 32900
rect 78492 32956 78756 32966
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78492 32890 78756 32900
rect 10872 32172 11136 32182
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 10872 32106 11136 32116
rect 30192 32172 30456 32182
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30192 32106 30456 32116
rect 49512 32172 49776 32182
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49512 32106 49776 32116
rect 68832 32172 69096 32182
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 68832 32106 69096 32116
rect 20532 31388 20796 31398
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20532 31322 20796 31332
rect 39852 31388 40116 31398
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 39852 31322 40116 31332
rect 59172 31388 59436 31398
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59172 31322 59436 31332
rect 78492 31388 78756 31398
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78492 31322 78756 31332
rect 10872 30604 11136 30614
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 10872 30538 11136 30548
rect 30192 30604 30456 30614
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30192 30538 30456 30548
rect 49512 30604 49776 30614
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49512 30538 49776 30548
rect 68832 30604 69096 30614
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 68832 30538 69096 30548
rect 20532 29820 20796 29830
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20532 29754 20796 29764
rect 39852 29820 40116 29830
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 39852 29754 40116 29764
rect 59172 29820 59436 29830
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59172 29754 59436 29764
rect 78492 29820 78756 29830
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78492 29754 78756 29764
rect 10872 29036 11136 29046
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 10872 28970 11136 28980
rect 30192 29036 30456 29046
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30192 28970 30456 28980
rect 49512 29036 49776 29046
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49512 28970 49776 28980
rect 68832 29036 69096 29046
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 68832 28970 69096 28980
rect 20532 28252 20796 28262
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20532 28186 20796 28196
rect 39852 28252 40116 28262
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 39852 28186 40116 28196
rect 59172 28252 59436 28262
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59172 28186 59436 28196
rect 78492 28252 78756 28262
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78492 28186 78756 28196
rect 10872 27468 11136 27478
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 10872 27402 11136 27412
rect 30192 27468 30456 27478
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30192 27402 30456 27412
rect 49512 27468 49776 27478
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49512 27402 49776 27412
rect 68832 27468 69096 27478
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 68832 27402 69096 27412
rect 20532 26684 20796 26694
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20532 26618 20796 26628
rect 39852 26684 40116 26694
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 39852 26618 40116 26628
rect 59172 26684 59436 26694
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59172 26618 59436 26628
rect 78492 26684 78756 26694
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78492 26618 78756 26628
rect 10872 25900 11136 25910
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 10872 25834 11136 25844
rect 30192 25900 30456 25910
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30192 25834 30456 25844
rect 49512 25900 49776 25910
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49512 25834 49776 25844
rect 68832 25900 69096 25910
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 68832 25834 69096 25844
rect 20532 25116 20796 25126
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20532 25050 20796 25060
rect 39852 25116 40116 25126
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 39852 25050 40116 25060
rect 59172 25116 59436 25126
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59172 25050 59436 25060
rect 78492 25116 78756 25126
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78492 25050 78756 25060
rect 10872 24332 11136 24342
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 10872 24266 11136 24276
rect 30192 24332 30456 24342
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30192 24266 30456 24276
rect 49512 24332 49776 24342
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49512 24266 49776 24276
rect 68832 24332 69096 24342
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 68832 24266 69096 24276
rect 20532 23548 20796 23558
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20532 23482 20796 23492
rect 39852 23548 40116 23558
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 39852 23482 40116 23492
rect 59172 23548 59436 23558
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59172 23482 59436 23492
rect 78492 23548 78756 23558
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78492 23482 78756 23492
rect 10872 22764 11136 22774
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 10872 22698 11136 22708
rect 30192 22764 30456 22774
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30192 22698 30456 22708
rect 49512 22764 49776 22774
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49512 22698 49776 22708
rect 68832 22764 69096 22774
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 68832 22698 69096 22708
rect 20532 21980 20796 21990
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20532 21914 20796 21924
rect 39852 21980 40116 21990
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 39852 21914 40116 21924
rect 59172 21980 59436 21990
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59172 21914 59436 21924
rect 78492 21980 78756 21990
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78492 21914 78756 21924
rect 10872 21196 11136 21206
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 10872 21130 11136 21140
rect 30192 21196 30456 21206
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30192 21130 30456 21140
rect 49512 21196 49776 21206
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49512 21130 49776 21140
rect 68832 21196 69096 21206
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 68832 21130 69096 21140
rect 20532 20412 20796 20422
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20532 20346 20796 20356
rect 39852 20412 40116 20422
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 39852 20346 40116 20356
rect 59172 20412 59436 20422
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59172 20346 59436 20356
rect 78492 20412 78756 20422
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78492 20346 78756 20356
rect 10872 19628 11136 19638
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 10872 19562 11136 19572
rect 30192 19628 30456 19638
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30192 19562 30456 19572
rect 49512 19628 49776 19638
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49512 19562 49776 19572
rect 68832 19628 69096 19638
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 68832 19562 69096 19572
rect 20532 18844 20796 18854
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20532 18778 20796 18788
rect 39852 18844 40116 18854
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 39852 18778 40116 18788
rect 59172 18844 59436 18854
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59172 18778 59436 18788
rect 78492 18844 78756 18854
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78492 18778 78756 18788
rect 16716 18564 16772 18574
rect 16604 18508 16716 18564
rect 10872 18060 11136 18070
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 10872 17994 11136 18004
rect 4844 17444 4900 17454
rect 4732 6578 4788 6590
rect 4732 6526 4734 6578
rect 4786 6526 4788 6578
rect 4508 6468 4564 6478
rect 4732 6468 4788 6526
rect 4508 6466 4788 6468
rect 4508 6414 4510 6466
rect 4562 6414 4788 6466
rect 4508 6412 4788 6414
rect 4508 6402 4564 6412
rect 3836 5572 3892 5582
rect 2492 5292 2884 5348
rect 2492 5234 2548 5292
rect 2492 5182 2494 5234
rect 2546 5182 2548 5234
rect 2492 5170 2548 5182
rect 2604 5124 2660 5134
rect 2044 4898 2100 4910
rect 2044 4846 2046 4898
rect 2098 4846 2100 4898
rect 2044 4340 2100 4846
rect 2492 4564 2548 4574
rect 2604 4564 2660 5068
rect 2492 4562 2660 4564
rect 2492 4510 2494 4562
rect 2546 4510 2660 4562
rect 2492 4508 2660 4510
rect 2492 4498 2548 4508
rect 2268 4340 2324 4350
rect 2044 4284 2268 4340
rect 2268 4246 2324 4284
rect 1932 4228 1988 4238
rect 1932 4226 2100 4228
rect 1932 4174 1934 4226
rect 1986 4174 2100 4226
rect 1932 4172 2100 4174
rect 1932 4162 1988 4172
rect 2044 3556 2100 4172
rect 2492 3780 2548 3790
rect 2268 3556 2324 3566
rect 2044 3500 2268 3556
rect 2268 3462 2324 3500
rect 1932 3444 1988 3454
rect 1932 3350 1988 3388
rect 2492 3442 2548 3724
rect 2492 3390 2494 3442
rect 2546 3390 2548 3442
rect 2492 3378 2548 3390
rect 2828 3442 2884 5292
rect 3836 5234 3892 5516
rect 4732 5460 4788 6412
rect 4732 5394 4788 5404
rect 3836 5182 3838 5234
rect 3890 5182 3892 5234
rect 3836 5170 3892 5182
rect 2940 5122 2996 5134
rect 2940 5070 2942 5122
rect 2994 5070 2996 5122
rect 2940 3668 2996 5070
rect 3388 5122 3444 5134
rect 3388 5070 3390 5122
rect 3442 5070 3444 5122
rect 3388 4900 3444 5070
rect 4620 5122 4676 5134
rect 4620 5070 4622 5122
rect 4674 5070 4676 5122
rect 3388 4834 3444 4844
rect 4284 4898 4340 4910
rect 4284 4846 4286 4898
rect 4338 4846 4340 4898
rect 4284 4452 4340 4846
rect 4620 4900 4676 5070
rect 4844 5012 4900 17388
rect 10872 16492 11136 16502
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 10872 16426 11136 16436
rect 4956 15316 5012 15326
rect 4956 5348 5012 15260
rect 6412 15204 6468 15214
rect 16604 15148 16660 18508
rect 16716 18498 16772 18508
rect 54572 18564 54628 18574
rect 30192 18060 30456 18070
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30192 17994 30456 18004
rect 49512 18060 49776 18070
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49512 17994 49776 18004
rect 20532 17276 20796 17286
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 39852 17276 40116 17286
rect 20532 17210 20796 17220
rect 37772 17220 37828 17230
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 39852 17210 40116 17220
rect 6300 8036 6356 8046
rect 6188 8034 6356 8036
rect 6188 7982 6302 8034
rect 6354 7982 6356 8034
rect 6188 7980 6356 7982
rect 6076 7588 6132 7598
rect 6076 7494 6132 7532
rect 5852 7474 5908 7486
rect 5852 7422 5854 7474
rect 5906 7422 5908 7474
rect 5516 7362 5572 7374
rect 5516 7310 5518 7362
rect 5570 7310 5572 7362
rect 5068 6916 5124 6926
rect 5068 6578 5124 6860
rect 5516 6692 5572 7310
rect 5852 7364 5908 7422
rect 5852 7298 5908 7308
rect 5740 6692 5796 6702
rect 5516 6690 5796 6692
rect 5516 6638 5742 6690
rect 5794 6638 5796 6690
rect 5516 6636 5796 6638
rect 5068 6526 5070 6578
rect 5122 6526 5124 6578
rect 5068 6514 5124 6526
rect 5068 5684 5124 5694
rect 5068 5590 5124 5628
rect 5628 5348 5684 5358
rect 4956 5292 5236 5348
rect 5068 5122 5124 5134
rect 5068 5070 5070 5122
rect 5122 5070 5124 5122
rect 5068 5012 5124 5070
rect 4844 4956 5124 5012
rect 5180 4900 5236 5292
rect 4620 4834 4676 4844
rect 4956 4844 5236 4900
rect 4284 4386 4340 4396
rect 3276 4226 3332 4238
rect 3276 4174 3278 4226
rect 3330 4174 3332 4226
rect 3276 3892 3332 4174
rect 4844 4226 4900 4238
rect 4844 4174 4846 4226
rect 4898 4174 4900 4226
rect 4844 4116 4900 4174
rect 4844 4050 4900 4060
rect 3500 3892 3556 3902
rect 3276 3826 3332 3836
rect 3388 3836 3500 3892
rect 2940 3602 2996 3612
rect 3388 3556 3444 3836
rect 3500 3826 3556 3836
rect 4956 3666 5012 4844
rect 5628 4338 5684 5292
rect 5740 5012 5796 6636
rect 5964 6468 6020 6478
rect 5852 6466 6020 6468
rect 5852 6414 5966 6466
rect 6018 6414 6020 6466
rect 5852 6412 6020 6414
rect 5852 5236 5908 6412
rect 5964 6402 6020 6412
rect 6076 6244 6132 6254
rect 5964 6132 6020 6142
rect 5964 5906 6020 6076
rect 5964 5854 5966 5906
rect 6018 5854 6020 5906
rect 5964 5842 6020 5854
rect 5852 5170 5908 5180
rect 5964 5236 6020 5246
rect 6076 5236 6132 6188
rect 6188 6132 6244 7980
rect 6300 7970 6356 7980
rect 6300 6692 6356 6702
rect 6300 6598 6356 6636
rect 6412 6356 6468 15148
rect 16044 15092 16660 15148
rect 20188 17108 20244 17118
rect 10872 14924 11136 14934
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 10872 14858 11136 14868
rect 10444 13748 10500 13758
rect 9548 12964 9604 12974
rect 9548 10610 9604 12908
rect 10108 12964 10164 12974
rect 10108 12870 10164 12908
rect 9772 12404 9828 12414
rect 9548 10558 9550 10610
rect 9602 10558 9604 10610
rect 9548 10546 9604 10558
rect 9660 12348 9772 12404
rect 9548 10052 9604 10062
rect 9436 9940 9492 9950
rect 9548 9940 9604 9996
rect 8988 9938 9604 9940
rect 8988 9886 9438 9938
rect 9490 9886 9604 9938
rect 8988 9884 9604 9886
rect 6748 9492 6804 9502
rect 6524 7364 6580 7374
rect 6524 6804 6580 7308
rect 6524 6738 6580 6748
rect 6636 6692 6692 6702
rect 6636 6578 6692 6636
rect 6636 6526 6638 6578
rect 6690 6526 6692 6578
rect 6636 6514 6692 6526
rect 6188 6066 6244 6076
rect 6300 6300 6468 6356
rect 5964 5234 6132 5236
rect 5964 5182 5966 5234
rect 6018 5182 6132 5234
rect 5964 5180 6132 5182
rect 6188 5236 6244 5246
rect 5964 5170 6020 5180
rect 6188 5142 6244 5180
rect 5740 4946 5796 4956
rect 5628 4286 5630 4338
rect 5682 4286 5684 4338
rect 5628 4274 5684 4286
rect 4956 3614 4958 3666
rect 5010 3614 5012 3666
rect 4956 3602 5012 3614
rect 5628 4004 5684 4014
rect 5628 3668 5684 3948
rect 3388 3490 3444 3500
rect 3612 3556 3668 3566
rect 3612 3462 3668 3500
rect 4060 3554 4116 3566
rect 4060 3502 4062 3554
rect 4114 3502 4116 3554
rect 2828 3390 2830 3442
rect 2882 3390 2884 3442
rect 2828 2548 2884 3390
rect 3164 3330 3220 3342
rect 3164 3278 3166 3330
rect 3218 3278 3220 3330
rect 2940 2548 2996 2558
rect 2828 2492 2940 2548
rect 2940 2482 2996 2492
rect 3164 2436 3220 3278
rect 4060 2660 4116 3502
rect 4508 3554 4564 3566
rect 4508 3502 4510 3554
rect 4562 3502 4564 3554
rect 4508 3444 4564 3502
rect 5628 3554 5684 3612
rect 5628 3502 5630 3554
rect 5682 3502 5684 3554
rect 5628 3490 5684 3502
rect 4508 3378 4564 3388
rect 4060 2594 4116 2604
rect 5852 3330 5908 3342
rect 5852 3278 5854 3330
rect 5906 3278 5908 3330
rect 3164 2370 3220 2380
rect 5852 1092 5908 3278
rect 5852 1026 5908 1036
rect 6300 800 6356 6300
rect 6748 5346 6804 9436
rect 8540 8930 8596 8942
rect 8540 8878 8542 8930
rect 8594 8878 8596 8930
rect 8540 8372 8596 8878
rect 8204 8316 8540 8372
rect 8092 8148 8148 8158
rect 7980 8146 8148 8148
rect 7980 8094 8094 8146
rect 8146 8094 8148 8146
rect 7980 8092 8148 8094
rect 7420 8036 7476 8046
rect 7868 8036 7924 8046
rect 7196 8034 7476 8036
rect 7196 7982 7422 8034
rect 7474 7982 7476 8034
rect 7196 7980 7476 7982
rect 6972 7476 7028 7486
rect 7196 7476 7252 7980
rect 7420 7970 7476 7980
rect 7644 8034 7924 8036
rect 7644 7982 7870 8034
rect 7922 7982 7924 8034
rect 7644 7980 7924 7982
rect 6972 7474 7252 7476
rect 6972 7422 6974 7474
rect 7026 7422 7252 7474
rect 6972 7420 7252 7422
rect 7308 7586 7364 7598
rect 7308 7534 7310 7586
rect 7362 7534 7364 7586
rect 6972 6356 7028 7420
rect 7084 6690 7140 6702
rect 7084 6638 7086 6690
rect 7138 6638 7140 6690
rect 7084 6580 7140 6638
rect 7140 6524 7252 6580
rect 7084 6514 7140 6524
rect 7084 6356 7140 6366
rect 6972 6300 7084 6356
rect 7084 6290 7140 6300
rect 7196 6244 7252 6524
rect 7196 6178 7252 6188
rect 6748 5294 6750 5346
rect 6802 5294 6804 5346
rect 6748 5282 6804 5294
rect 6860 5684 6916 5694
rect 6412 5124 6468 5134
rect 6412 5030 6468 5068
rect 6524 4900 6580 4910
rect 6524 800 6580 4844
rect 6860 2884 6916 5628
rect 7084 5684 7140 5694
rect 7084 5348 7140 5628
rect 7084 5234 7140 5292
rect 7084 5182 7086 5234
rect 7138 5182 7140 5234
rect 7084 5170 7140 5182
rect 7308 4564 7364 7534
rect 7644 6244 7700 7980
rect 7868 7970 7924 7980
rect 7756 7700 7812 7710
rect 7980 7700 8036 8092
rect 8092 8082 8148 8092
rect 7756 7698 8036 7700
rect 7756 7646 7758 7698
rect 7810 7646 8036 7698
rect 7756 7644 8036 7646
rect 7756 7634 7812 7644
rect 8092 7476 8148 7486
rect 8204 7476 8260 8316
rect 8540 8306 8596 8316
rect 8988 8260 9044 9884
rect 9436 9874 9492 9884
rect 9100 8930 9156 8942
rect 9100 8878 9102 8930
rect 9154 8878 9156 8930
rect 9100 8484 9156 8878
rect 9100 8428 9604 8484
rect 9100 8260 9156 8270
rect 8988 8258 9156 8260
rect 8988 8206 9102 8258
rect 9154 8206 9156 8258
rect 8988 8204 9156 8206
rect 9100 8148 9156 8204
rect 9100 8092 9268 8148
rect 8428 8036 8484 8046
rect 8428 8034 9156 8036
rect 8428 7982 8430 8034
rect 8482 7982 9156 8034
rect 8428 7980 9156 7982
rect 8428 7970 8484 7980
rect 8092 7474 8260 7476
rect 8092 7422 8094 7474
rect 8146 7422 8260 7474
rect 8092 7420 8260 7422
rect 8764 7586 8820 7598
rect 8764 7534 8766 7586
rect 8818 7534 8820 7586
rect 8092 7410 8148 7420
rect 7756 6692 7812 6702
rect 7756 6598 7812 6636
rect 7644 6178 7700 6188
rect 8652 6356 8708 6366
rect 7980 5682 8036 5694
rect 7980 5630 7982 5682
rect 8034 5630 8036 5682
rect 7756 5460 7812 5470
rect 7308 4498 7364 4508
rect 7420 5012 7476 5022
rect 6748 2828 6916 2884
rect 6972 3556 7028 3566
rect 6748 800 6804 2828
rect 6972 800 7028 3500
rect 7196 3444 7252 3454
rect 7196 800 7252 3388
rect 7420 800 7476 4956
rect 7756 4004 7812 5404
rect 7868 4228 7924 4238
rect 7868 4134 7924 4172
rect 7756 3948 7924 4004
rect 7756 3666 7812 3678
rect 7756 3614 7758 3666
rect 7810 3614 7812 3666
rect 7756 3444 7812 3614
rect 7756 3378 7812 3388
rect 7868 800 7924 3948
rect 7980 3388 8036 5630
rect 8316 4340 8372 4350
rect 7980 3332 8148 3388
rect 8092 800 8148 3332
rect 8316 800 8372 4284
rect 8652 3388 8708 6300
rect 8764 5684 8820 7534
rect 8876 7474 8932 7486
rect 8876 7422 8878 7474
rect 8930 7422 8932 7474
rect 8876 6020 8932 7422
rect 8876 5954 8932 5964
rect 8988 5908 9044 5918
rect 8988 5814 9044 5852
rect 8764 5618 8820 5628
rect 8988 5684 9044 5694
rect 8764 4900 8820 4910
rect 8764 3554 8820 4844
rect 8988 4338 9044 5628
rect 9100 5236 9156 7980
rect 9212 6580 9268 8092
rect 9548 7476 9604 8428
rect 9660 8036 9716 12348
rect 9772 12338 9828 12348
rect 10332 10498 10388 10510
rect 10332 10446 10334 10498
rect 10386 10446 10388 10498
rect 10220 9716 10276 9726
rect 10332 9716 10388 10446
rect 10220 9714 10388 9716
rect 10220 9662 10222 9714
rect 10274 9662 10388 9714
rect 10220 9660 10388 9662
rect 10220 9650 10276 9660
rect 9996 9604 10052 9614
rect 9884 9602 10052 9604
rect 9884 9550 9998 9602
rect 10050 9550 10052 9602
rect 9884 9548 10052 9550
rect 9772 9044 9828 9054
rect 9884 9044 9940 9548
rect 9996 9538 10052 9548
rect 9772 9042 9940 9044
rect 9772 8990 9774 9042
rect 9826 8990 9940 9042
rect 9772 8988 9940 8990
rect 9996 9154 10052 9166
rect 9996 9102 9998 9154
rect 10050 9102 10052 9154
rect 9772 8484 9828 8988
rect 9996 8820 10052 9102
rect 9996 8754 10052 8764
rect 10332 9154 10388 9166
rect 10332 9102 10334 9154
rect 10386 9102 10388 9154
rect 9772 8428 10164 8484
rect 9884 8260 9940 8298
rect 10108 8260 10164 8428
rect 10332 8260 10388 9102
rect 10444 8820 10500 13692
rect 13244 13634 13300 13646
rect 13244 13582 13246 13634
rect 13298 13582 13300 13634
rect 10872 13356 11136 13366
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 10872 13290 11136 13300
rect 12908 13074 12964 13086
rect 12908 13022 12910 13074
rect 12962 13022 12964 13074
rect 10780 12852 10836 12862
rect 10780 12850 11284 12852
rect 10780 12798 10782 12850
rect 10834 12798 11284 12850
rect 10780 12796 11284 12798
rect 10780 12786 10836 12796
rect 11228 12402 11284 12796
rect 11228 12350 11230 12402
rect 11282 12350 11284 12402
rect 11228 12338 11284 12350
rect 12908 12290 12964 13022
rect 12908 12238 12910 12290
rect 12962 12238 12964 12290
rect 11564 12180 11620 12190
rect 12012 12180 12068 12190
rect 11564 12178 12068 12180
rect 11564 12126 11566 12178
rect 11618 12126 12014 12178
rect 12066 12126 12068 12178
rect 11564 12124 12068 12126
rect 11564 12114 11620 12124
rect 12012 12114 12068 12124
rect 12348 11954 12404 11966
rect 12348 11902 12350 11954
rect 12402 11902 12404 11954
rect 11676 11844 11732 11854
rect 10872 11788 11136 11798
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 10872 11722 11136 11732
rect 10872 10220 11136 10230
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 10872 10154 11136 10164
rect 11564 9826 11620 9838
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 10556 9716 10612 9726
rect 11228 9716 11284 9726
rect 10556 9714 11284 9716
rect 10556 9662 10558 9714
rect 10610 9662 11230 9714
rect 11282 9662 11284 9714
rect 10556 9660 11284 9662
rect 10556 9650 10612 9660
rect 11228 9650 11284 9660
rect 11452 9716 11508 9726
rect 10668 9044 10724 9054
rect 11116 9044 11172 9054
rect 10668 9042 11172 9044
rect 10668 8990 10670 9042
rect 10722 8990 11118 9042
rect 11170 8990 11172 9042
rect 10668 8988 11172 8990
rect 10668 8978 10724 8988
rect 11116 8978 11172 8988
rect 11452 9042 11508 9660
rect 11564 9604 11620 9774
rect 11564 9538 11620 9548
rect 11452 8990 11454 9042
rect 11506 8990 11508 9042
rect 11452 8978 11508 8990
rect 10444 8764 10724 8820
rect 10108 8204 10276 8260
rect 9884 8194 9940 8204
rect 9660 7980 10052 8036
rect 9996 7698 10052 7980
rect 9996 7646 9998 7698
rect 10050 7646 10052 7698
rect 9996 7634 10052 7646
rect 9660 7476 9716 7486
rect 9548 7474 9716 7476
rect 9548 7422 9662 7474
rect 9714 7422 9716 7474
rect 9548 7420 9716 7422
rect 9212 6514 9268 6524
rect 9436 6804 9492 6814
rect 9324 5572 9380 5582
rect 9212 5236 9268 5246
rect 9100 5234 9268 5236
rect 9100 5182 9214 5234
rect 9266 5182 9268 5234
rect 9100 5180 9268 5182
rect 9212 5170 9268 5180
rect 8988 4286 8990 4338
rect 9042 4286 9044 4338
rect 8988 4274 9044 4286
rect 8764 3502 8766 3554
rect 8818 3502 8820 3554
rect 8764 3490 8820 3502
rect 8876 4228 8932 4238
rect 8876 3388 8932 4172
rect 9324 4004 9380 5516
rect 9212 3892 9268 3902
rect 8652 3332 8820 3388
rect 8876 3332 9044 3388
rect 8764 800 8820 3332
rect 8988 800 9044 3332
rect 9212 800 9268 3836
rect 9324 3554 9380 3948
rect 9324 3502 9326 3554
rect 9378 3502 9380 3554
rect 9324 3490 9380 3502
rect 9436 2772 9492 6748
rect 9548 6356 9604 7420
rect 9660 7410 9716 7420
rect 9884 6804 9940 6814
rect 9772 6802 9940 6804
rect 9772 6750 9886 6802
rect 9938 6750 9940 6802
rect 9772 6748 9940 6750
rect 9548 6290 9604 6300
rect 9660 6468 9716 6478
rect 9660 6130 9716 6412
rect 9660 6078 9662 6130
rect 9714 6078 9716 6130
rect 9660 6066 9716 6078
rect 9772 5684 9828 6748
rect 9884 6738 9940 6748
rect 9772 5618 9828 5628
rect 9884 6580 9940 6590
rect 9548 5236 9604 5246
rect 9548 4338 9604 5180
rect 9884 5124 9940 6524
rect 9996 6244 10052 6254
rect 9996 5906 10052 6188
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9996 5842 10052 5854
rect 9884 5030 9940 5068
rect 9548 4286 9550 4338
rect 9602 4286 9604 4338
rect 9548 4274 9604 4286
rect 9772 4114 9828 4126
rect 9772 4062 9774 4114
rect 9826 4062 9828 4114
rect 9772 3780 9828 4062
rect 9772 3714 9828 3724
rect 9884 4116 9940 4126
rect 9660 3330 9716 3342
rect 9660 3278 9662 3330
rect 9714 3278 9716 3330
rect 9660 2996 9716 3278
rect 9660 2930 9716 2940
rect 9436 2716 9716 2772
rect 9660 800 9716 2716
rect 9884 800 9940 4060
rect 10108 4114 10164 4126
rect 10108 4062 10110 4114
rect 10162 4062 10164 4114
rect 10108 1204 10164 4062
rect 10220 3388 10276 8204
rect 10332 8194 10388 8204
rect 10444 7700 10500 7710
rect 10444 7474 10500 7644
rect 10668 7698 10724 8764
rect 10872 8652 11136 8662
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 10872 8586 11136 8596
rect 10668 7646 10670 7698
rect 10722 7646 10724 7698
rect 10668 7634 10724 7646
rect 10444 7422 10446 7474
rect 10498 7422 10500 7474
rect 10444 7410 10500 7422
rect 11228 7250 11284 7262
rect 11228 7198 11230 7250
rect 11282 7198 11284 7250
rect 10872 7084 11136 7094
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 10872 7018 11136 7028
rect 10332 6020 10388 6030
rect 10332 5926 10388 5964
rect 10556 6018 10612 6030
rect 10556 5966 10558 6018
rect 10610 5966 10612 6018
rect 10556 5684 10612 5966
rect 10556 5618 10612 5628
rect 10872 5516 11136 5526
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 10872 5450 11136 5460
rect 10892 5348 10948 5358
rect 10668 4564 10724 4574
rect 10668 4470 10724 4508
rect 10892 4226 10948 5292
rect 10892 4174 10894 4226
rect 10946 4174 10948 4226
rect 10892 4162 10948 4174
rect 10872 3948 11136 3958
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 10872 3882 11136 3892
rect 11228 3780 11284 7198
rect 11676 6692 11732 11788
rect 12124 11284 12180 11294
rect 12124 9826 12180 11228
rect 12236 11170 12292 11182
rect 12236 11118 12238 11170
rect 12290 11118 12292 11170
rect 12236 10500 12292 11118
rect 12348 11172 12404 11902
rect 12908 11844 12964 12238
rect 13244 12964 13300 13582
rect 14924 13524 14980 13534
rect 14812 13468 14924 13524
rect 12908 11778 12964 11788
rect 13132 12178 13188 12190
rect 13132 12126 13134 12178
rect 13186 12126 13188 12178
rect 13132 11284 13188 12126
rect 13132 11218 13188 11228
rect 12348 11106 12404 11116
rect 12236 10434 12292 10444
rect 12460 10498 12516 10510
rect 12460 10446 12462 10498
rect 12514 10446 12516 10498
rect 12124 9774 12126 9826
rect 12178 9774 12180 9826
rect 12012 9154 12068 9166
rect 12012 9102 12014 9154
rect 12066 9102 12068 9154
rect 12012 8370 12068 9102
rect 12124 9044 12180 9774
rect 12348 9716 12404 9726
rect 12460 9716 12516 10446
rect 12908 10498 12964 10510
rect 12908 10446 12910 10498
rect 12962 10446 12964 10498
rect 12908 10164 12964 10446
rect 13244 10164 13300 12908
rect 13580 12962 13636 12974
rect 13580 12910 13582 12962
rect 13634 12910 13636 12962
rect 13580 11956 13636 12910
rect 13804 12740 13860 12750
rect 13804 12738 14420 12740
rect 13804 12686 13806 12738
rect 13858 12686 14420 12738
rect 13804 12684 14420 12686
rect 13804 12674 13860 12684
rect 14364 12290 14420 12684
rect 14364 12238 14366 12290
rect 14418 12238 14420 12290
rect 14364 12226 14420 12238
rect 13692 12180 13748 12190
rect 13692 12086 13748 12124
rect 13580 11900 14196 11956
rect 14140 11618 14196 11900
rect 14140 11566 14142 11618
rect 14194 11566 14196 11618
rect 14140 11554 14196 11566
rect 14476 11394 14532 11406
rect 14476 11342 14478 11394
rect 14530 11342 14532 11394
rect 13580 11172 13636 11182
rect 12908 10108 13244 10164
rect 13244 10098 13300 10108
rect 13356 10498 13412 10510
rect 13356 10446 13358 10498
rect 13410 10446 13412 10498
rect 13356 9716 13412 10446
rect 13580 10276 13636 11116
rect 14476 10724 14532 11342
rect 14700 11284 14756 11294
rect 14700 11190 14756 11228
rect 14476 10658 14532 10668
rect 14028 10500 14084 10510
rect 14028 10406 14084 10444
rect 13580 10210 13636 10220
rect 12348 9714 12628 9716
rect 12348 9662 12350 9714
rect 12402 9662 12628 9714
rect 12348 9660 12628 9662
rect 12348 9650 12404 9660
rect 12124 8950 12180 8988
rect 12012 8318 12014 8370
rect 12066 8318 12068 8370
rect 11788 7700 11844 7710
rect 11844 7644 11956 7700
rect 11788 7634 11844 7644
rect 11676 6636 11844 6692
rect 11340 6580 11396 6590
rect 11340 6578 11732 6580
rect 11340 6526 11342 6578
rect 11394 6526 11732 6578
rect 11340 6524 11732 6526
rect 11340 6514 11396 6524
rect 10780 3724 11284 3780
rect 11452 6356 11508 6366
rect 10220 3332 10612 3388
rect 10108 1138 10164 1148
rect 10556 800 10612 3332
rect 10780 800 10836 3724
rect 11452 800 11508 6300
rect 11564 3668 11620 3678
rect 11564 3574 11620 3612
rect 11676 800 11732 6524
rect 11788 5906 11844 6636
rect 11788 5854 11790 5906
rect 11842 5854 11844 5906
rect 11788 5842 11844 5854
rect 11900 5684 11956 7644
rect 12012 6692 12068 8318
rect 12460 8258 12516 8270
rect 12460 8206 12462 8258
rect 12514 8206 12516 8258
rect 12460 6916 12516 8206
rect 12460 6850 12516 6860
rect 12460 6692 12516 6702
rect 12012 6690 12516 6692
rect 12012 6638 12462 6690
rect 12514 6638 12516 6690
rect 12012 6636 12516 6638
rect 12460 6626 12516 6636
rect 11788 5628 11956 5684
rect 11788 3332 11844 5628
rect 12572 5122 12628 9660
rect 13356 9650 13412 9660
rect 14364 9714 14420 9726
rect 14364 9662 14366 9714
rect 14418 9662 14420 9714
rect 12908 9604 12964 9614
rect 13580 9604 13636 9614
rect 12908 8932 12964 9548
rect 13468 9602 13636 9604
rect 13468 9550 13582 9602
rect 13634 9550 13636 9602
rect 13468 9548 13636 9550
rect 13356 9042 13412 9054
rect 13356 8990 13358 9042
rect 13410 8990 13412 9042
rect 12908 8866 12964 8876
rect 13020 8932 13076 8942
rect 13356 8932 13412 8990
rect 13020 8930 13412 8932
rect 13020 8878 13022 8930
rect 13074 8878 13412 8930
rect 13020 8876 13412 8878
rect 13020 8866 13076 8876
rect 12684 8036 12740 8046
rect 12684 8034 13076 8036
rect 12684 7982 12686 8034
rect 12738 7982 13076 8034
rect 12684 7980 13076 7982
rect 12684 7970 12740 7980
rect 12572 5070 12574 5122
rect 12626 5070 12628 5122
rect 12572 5058 12628 5070
rect 12684 5796 12740 5806
rect 11900 4900 11956 4910
rect 11900 4898 12404 4900
rect 11900 4846 11902 4898
rect 11954 4846 12404 4898
rect 11900 4844 12404 4846
rect 11900 4834 11956 4844
rect 11788 3276 12180 3332
rect 12124 800 12180 3276
rect 12348 800 12404 4844
rect 12572 3556 12628 3566
rect 12684 3556 12740 5740
rect 12572 3554 12740 3556
rect 12572 3502 12574 3554
rect 12626 3502 12740 3554
rect 12572 3500 12740 3502
rect 12796 5682 12852 5694
rect 12796 5630 12798 5682
rect 12850 5630 12852 5682
rect 12572 3490 12628 3500
rect 12796 3388 12852 5630
rect 13020 4450 13076 7980
rect 13132 7474 13188 7486
rect 13132 7422 13134 7474
rect 13186 7422 13188 7474
rect 13132 6580 13188 7422
rect 13356 7140 13412 8876
rect 13468 7700 13524 9548
rect 13580 9538 13636 9548
rect 14140 9604 14196 9614
rect 14364 9604 14420 9662
rect 14700 9716 14756 9726
rect 14812 9716 14868 13468
rect 14924 13458 14980 13468
rect 15260 12180 15316 12190
rect 15148 11284 15204 11294
rect 15148 11190 15204 11228
rect 14700 9714 14868 9716
rect 14700 9662 14702 9714
rect 14754 9662 14868 9714
rect 14700 9660 14868 9662
rect 15036 10498 15092 10510
rect 15036 10446 15038 10498
rect 15090 10446 15092 10498
rect 14700 9650 14756 9660
rect 14140 9602 14420 9604
rect 14140 9550 14142 9602
rect 14194 9550 14420 9602
rect 14140 9548 14420 9550
rect 14140 9538 14196 9548
rect 13580 9154 13636 9166
rect 13580 9102 13582 9154
rect 13634 9102 13636 9154
rect 13580 8484 13636 9102
rect 14028 9044 14084 9054
rect 13580 8418 13636 8428
rect 13916 8930 13972 8942
rect 13916 8878 13918 8930
rect 13970 8878 13972 8930
rect 13804 8148 13860 8158
rect 13804 8054 13860 8092
rect 13468 7634 13524 7644
rect 13916 7140 13972 8878
rect 14028 8370 14084 8988
rect 14028 8318 14030 8370
rect 14082 8318 14084 8370
rect 14028 8306 14084 8318
rect 14140 7250 14196 7262
rect 14140 7198 14142 7250
rect 14194 7198 14196 7250
rect 13356 7084 13524 7140
rect 13916 7084 14084 7140
rect 13132 6514 13188 6524
rect 13468 6356 13524 7084
rect 13916 6690 13972 6702
rect 13916 6638 13918 6690
rect 13970 6638 13972 6690
rect 13692 6580 13748 6590
rect 13468 6300 13636 6356
rect 13020 4398 13022 4450
rect 13074 4398 13076 4450
rect 13020 4386 13076 4398
rect 13132 4452 13188 4462
rect 13132 3556 13188 4396
rect 13132 3462 13188 3500
rect 12796 3332 13076 3388
rect 12796 2548 12852 2558
rect 12796 800 12852 2492
rect 13020 800 13076 3332
rect 13468 3332 13524 3342
rect 13468 3238 13524 3276
rect 13580 3108 13636 6300
rect 13692 5348 13748 6524
rect 13916 6020 13972 6638
rect 13916 5954 13972 5964
rect 13916 5796 13972 5806
rect 14028 5796 14084 7084
rect 13972 5740 14084 5796
rect 13916 5730 13972 5740
rect 13692 5282 13748 5292
rect 13692 5124 13748 5134
rect 13692 4338 13748 5068
rect 13692 4286 13694 4338
rect 13746 4286 13748 4338
rect 13692 4274 13748 4286
rect 14140 4116 14196 7198
rect 13468 3052 13636 3108
rect 13692 4060 14196 4116
rect 13468 800 13524 3052
rect 13692 800 13748 4060
rect 13804 3332 13860 3342
rect 13804 1428 13860 3276
rect 14252 2212 14308 9548
rect 14588 8036 14644 8046
rect 14588 7942 14644 7980
rect 14364 7028 14420 7038
rect 14364 6914 14420 6972
rect 15036 7028 15092 10446
rect 15260 10052 15316 12124
rect 15820 11170 15876 11182
rect 15820 11118 15822 11170
rect 15874 11118 15876 11170
rect 15820 10724 15876 11118
rect 15820 10658 15876 10668
rect 15260 9828 15316 9996
rect 15372 9828 15428 9838
rect 15260 9826 15428 9828
rect 15260 9774 15374 9826
rect 15426 9774 15428 9826
rect 15260 9772 15428 9774
rect 15372 9762 15428 9772
rect 16044 9156 16100 15092
rect 19292 13972 19348 13982
rect 17948 13188 18004 13198
rect 17500 12180 17556 12190
rect 17500 12086 17556 12124
rect 16492 12066 16548 12078
rect 16492 12014 16494 12066
rect 16546 12014 16548 12066
rect 16492 11284 16548 12014
rect 16380 10500 16436 10510
rect 16380 10406 16436 10444
rect 16268 10164 16324 10174
rect 16156 9716 16212 9726
rect 16156 9622 16212 9660
rect 16044 9100 16212 9156
rect 16044 8930 16100 8942
rect 16044 8878 16046 8930
rect 16098 8878 16100 8930
rect 15148 8258 15204 8270
rect 15148 8206 15150 8258
rect 15202 8206 15204 8258
rect 15148 8036 15204 8206
rect 15372 8260 15428 8270
rect 15372 8146 15428 8204
rect 15372 8094 15374 8146
rect 15426 8094 15428 8146
rect 15372 8082 15428 8094
rect 15820 8258 15876 8270
rect 15820 8206 15822 8258
rect 15874 8206 15876 8258
rect 15260 8036 15316 8046
rect 15148 7980 15260 8036
rect 15036 6962 15092 6972
rect 15260 7476 15316 7980
rect 14364 6862 14366 6914
rect 14418 6862 14420 6914
rect 14364 6850 14420 6862
rect 14700 6692 14756 6702
rect 14700 6598 14756 6636
rect 15260 6690 15316 7420
rect 15260 6638 15262 6690
rect 15314 6638 15316 6690
rect 15260 6626 15316 6638
rect 15708 6690 15764 6702
rect 15708 6638 15710 6690
rect 15762 6638 15764 6690
rect 14476 6468 14532 6478
rect 14476 5234 14532 6412
rect 15708 6020 15764 6638
rect 15820 6244 15876 8206
rect 15820 6178 15876 6188
rect 15932 8148 15988 8158
rect 14476 5182 14478 5234
rect 14530 5182 14532 5234
rect 14476 5170 14532 5182
rect 15148 5794 15204 5806
rect 15148 5742 15150 5794
rect 15202 5742 15204 5794
rect 14924 4452 14980 4462
rect 13804 1362 13860 1372
rect 14140 2156 14308 2212
rect 14364 3444 14420 3454
rect 14140 800 14196 2156
rect 14364 800 14420 3388
rect 14812 3444 14868 3482
rect 14812 3378 14868 3388
rect 14924 2212 14980 4396
rect 15148 3444 15204 5742
rect 15708 5348 15764 5964
rect 15708 5282 15764 5292
rect 15708 4226 15764 4238
rect 15708 4174 15710 4226
rect 15762 4174 15764 4226
rect 14812 2156 14980 2212
rect 15036 3388 15204 3444
rect 15484 3780 15540 3790
rect 14812 800 14868 2156
rect 15036 800 15092 3388
rect 15484 800 15540 3724
rect 15708 800 15764 4174
rect 15932 3388 15988 8092
rect 16044 8034 16100 8878
rect 16044 7982 16046 8034
rect 16098 7982 16100 8034
rect 16044 7970 16100 7982
rect 16044 6802 16100 6814
rect 16044 6750 16046 6802
rect 16098 6750 16100 6802
rect 16044 5908 16100 6750
rect 16044 5124 16100 5852
rect 16156 6356 16212 9100
rect 16156 5684 16212 6300
rect 16268 5908 16324 10108
rect 16380 8258 16436 8270
rect 16380 8206 16382 8258
rect 16434 8206 16436 8258
rect 16380 8148 16436 8206
rect 16380 8082 16436 8092
rect 16492 7474 16548 11228
rect 16940 11620 16996 11630
rect 16940 10834 16996 11564
rect 17724 11172 17780 11182
rect 16940 10782 16942 10834
rect 16994 10782 16996 10834
rect 16828 10500 16884 10510
rect 16828 9042 16884 10444
rect 16828 8990 16830 9042
rect 16882 8990 16884 9042
rect 16492 7422 16494 7474
rect 16546 7422 16548 7474
rect 16492 7410 16548 7422
rect 16604 8148 16660 8158
rect 16604 6804 16660 8092
rect 16604 6738 16660 6748
rect 16716 8034 16772 8046
rect 16716 7982 16718 8034
rect 16770 7982 16772 8034
rect 16716 6468 16772 7982
rect 16828 7364 16884 8990
rect 16940 8258 16996 10782
rect 16940 8206 16942 8258
rect 16994 8206 16996 8258
rect 16940 8194 16996 8206
rect 17276 11170 17780 11172
rect 17276 11118 17726 11170
rect 17778 11118 17780 11170
rect 17276 11116 17780 11118
rect 16828 7298 16884 7308
rect 17164 8146 17220 8158
rect 17164 8094 17166 8146
rect 17218 8094 17220 8146
rect 16716 6402 16772 6412
rect 16828 6356 16884 6366
rect 16716 6132 16772 6142
rect 16380 5908 16436 5918
rect 16268 5906 16436 5908
rect 16268 5854 16382 5906
rect 16434 5854 16436 5906
rect 16268 5852 16436 5854
rect 16380 5842 16436 5852
rect 16156 5618 16212 5628
rect 16604 5236 16660 5246
rect 16044 5058 16100 5068
rect 16268 5180 16604 5236
rect 16156 5012 16212 5022
rect 15932 3332 16100 3388
rect 16044 2884 16100 3332
rect 16044 2818 16100 2828
rect 16156 800 16212 4956
rect 16268 3554 16324 5180
rect 16604 5142 16660 5180
rect 16716 4338 16772 6076
rect 16716 4286 16718 4338
rect 16770 4286 16772 4338
rect 16716 4274 16772 4286
rect 16268 3502 16270 3554
rect 16322 3502 16324 3554
rect 16268 3490 16324 3502
rect 16380 3668 16436 3678
rect 16380 800 16436 3612
rect 16828 800 16884 6300
rect 17164 5460 17220 8094
rect 17276 7028 17332 11116
rect 17724 11106 17780 11116
rect 17948 10836 18004 13132
rect 18284 12740 18340 12750
rect 17724 10834 18004 10836
rect 17724 10782 17950 10834
rect 18002 10782 18004 10834
rect 17724 10780 18004 10782
rect 17500 10500 17556 10510
rect 17500 10406 17556 10444
rect 17500 9716 17556 9726
rect 17500 9266 17556 9660
rect 17500 9214 17502 9266
rect 17554 9214 17556 9266
rect 17500 9202 17556 9214
rect 17724 9154 17780 10780
rect 17948 10770 18004 10780
rect 18172 12066 18228 12078
rect 18172 12014 18174 12066
rect 18226 12014 18228 12066
rect 18172 11284 18228 12014
rect 18172 10164 18228 11228
rect 18284 11170 18340 12684
rect 18844 11172 18900 11182
rect 18284 11118 18286 11170
rect 18338 11118 18340 11170
rect 18284 10500 18340 11118
rect 18620 11116 18844 11172
rect 18284 10434 18340 10444
rect 18508 10498 18564 10510
rect 18508 10446 18510 10498
rect 18562 10446 18564 10498
rect 18172 10098 18228 10108
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17724 9090 17780 9102
rect 18284 9938 18340 9950
rect 18284 9886 18286 9938
rect 18338 9886 18340 9938
rect 17388 9042 17444 9054
rect 17388 8990 17390 9042
rect 17442 8990 17444 9042
rect 17388 8148 17444 8990
rect 17836 9042 17892 9054
rect 17836 8990 17838 9042
rect 17890 8990 17892 9042
rect 17836 8482 17892 8990
rect 17836 8430 17838 8482
rect 17890 8430 17892 8482
rect 17836 8418 17892 8430
rect 17500 8260 17556 8270
rect 17836 8260 17892 8270
rect 17556 8204 17668 8260
rect 17500 8166 17556 8204
rect 17388 8082 17444 8092
rect 17612 7364 17668 8204
rect 17836 8258 18004 8260
rect 17836 8206 17838 8258
rect 17890 8206 18004 8258
rect 17836 8204 18004 8206
rect 17836 8194 17892 8204
rect 17724 7700 17780 7710
rect 17724 7606 17780 7644
rect 17612 7308 17780 7364
rect 17276 6972 17444 7028
rect 17164 5394 17220 5404
rect 17276 6804 17332 6814
rect 17276 5346 17332 6748
rect 17388 6356 17444 6972
rect 17388 6290 17444 6300
rect 17500 6244 17556 6254
rect 17556 6188 17668 6244
rect 17500 6178 17556 6188
rect 17612 6130 17668 6188
rect 17612 6078 17614 6130
rect 17666 6078 17668 6130
rect 17612 6066 17668 6078
rect 17724 6018 17780 7308
rect 17948 7252 18004 8204
rect 18172 8034 18228 8046
rect 18172 7982 18174 8034
rect 18226 7982 18228 8034
rect 18172 7476 18228 7982
rect 18172 7410 18228 7420
rect 18284 7252 18340 9886
rect 18508 8372 18564 10446
rect 18396 8316 18564 8372
rect 18396 7924 18452 8316
rect 18508 8148 18564 8158
rect 18620 8148 18676 11116
rect 18844 11078 18900 11116
rect 18732 10052 18788 10062
rect 18732 9938 18788 9996
rect 18732 9886 18734 9938
rect 18786 9886 18788 9938
rect 18732 9874 18788 9886
rect 19180 9604 19236 9614
rect 18956 9602 19236 9604
rect 18956 9550 19182 9602
rect 19234 9550 19236 9602
rect 18956 9548 19236 9550
rect 18844 9268 18900 9278
rect 18844 9174 18900 9212
rect 18508 8146 18676 8148
rect 18508 8094 18510 8146
rect 18562 8094 18676 8146
rect 18508 8092 18676 8094
rect 18508 8082 18564 8092
rect 18396 7868 18564 7924
rect 17948 7196 18340 7252
rect 18172 6580 18228 6590
rect 17724 5966 17726 6018
rect 17778 5966 17780 6018
rect 17724 5954 17780 5966
rect 17836 6578 18228 6580
rect 17836 6526 18174 6578
rect 18226 6526 18228 6578
rect 17836 6524 18228 6526
rect 17388 5908 17444 5946
rect 17388 5842 17444 5852
rect 17724 5684 17780 5694
rect 17276 5294 17278 5346
rect 17330 5294 17332 5346
rect 17276 5282 17332 5294
rect 17612 5572 17668 5582
rect 16940 5124 16996 5134
rect 16940 5030 16996 5068
rect 17164 4898 17220 4910
rect 17164 4846 17166 4898
rect 17218 4846 17220 4898
rect 17164 4452 17220 4846
rect 17388 4452 17444 4462
rect 17164 4450 17444 4452
rect 17164 4398 17390 4450
rect 17442 4398 17444 4450
rect 17164 4396 17444 4398
rect 17388 4386 17444 4396
rect 17612 4450 17668 5516
rect 17724 4898 17780 5628
rect 17724 4846 17726 4898
rect 17778 4846 17780 4898
rect 17724 4834 17780 4846
rect 17836 4562 17892 6524
rect 18172 6514 18228 6524
rect 18172 6018 18228 6030
rect 18172 5966 18174 6018
rect 18226 5966 18228 6018
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 18060 5124 18116 5134
rect 17612 4398 17614 4450
rect 17666 4398 17668 4450
rect 17612 4386 17668 4398
rect 18060 4338 18116 5068
rect 18060 4286 18062 4338
rect 18114 4286 18116 4338
rect 18060 4274 18116 4286
rect 17836 3892 17892 3902
rect 17612 3666 17668 3678
rect 17612 3614 17614 3666
rect 17666 3614 17668 3666
rect 17612 3388 17668 3614
rect 17052 3332 17108 3342
rect 16940 3330 17108 3332
rect 16940 3278 17054 3330
rect 17106 3278 17108 3330
rect 16940 3276 17108 3278
rect 16940 1092 16996 3276
rect 17052 3266 17108 3276
rect 17164 3332 17668 3388
rect 17164 1764 17220 3332
rect 17836 1876 17892 3836
rect 18172 3780 18228 5966
rect 18284 4564 18340 7196
rect 18508 6130 18564 7868
rect 18844 7364 18900 7374
rect 18844 6690 18900 7308
rect 18844 6638 18846 6690
rect 18898 6638 18900 6690
rect 18844 6626 18900 6638
rect 18508 6078 18510 6130
rect 18562 6078 18564 6130
rect 18508 5012 18564 6078
rect 18844 6020 18900 6030
rect 18508 4946 18564 4956
rect 18732 6018 18900 6020
rect 18732 5966 18846 6018
rect 18898 5966 18900 6018
rect 18732 5964 18900 5966
rect 18732 4676 18788 5964
rect 18844 5954 18900 5964
rect 18956 4788 19012 9548
rect 19180 9538 19236 9548
rect 19068 8932 19124 8942
rect 19068 8930 19236 8932
rect 19068 8878 19070 8930
rect 19122 8878 19236 8930
rect 19068 8876 19236 8878
rect 19068 8866 19124 8876
rect 19180 8258 19236 8876
rect 19180 8206 19182 8258
rect 19234 8206 19236 8258
rect 19180 6132 19236 8206
rect 19292 7028 19348 13916
rect 19404 12964 19460 12974
rect 19404 12962 19572 12964
rect 19404 12910 19406 12962
rect 19458 12910 19572 12962
rect 19404 12908 19572 12910
rect 19404 12898 19460 12908
rect 19516 11618 19572 12908
rect 19628 12738 19684 12750
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19628 12292 19684 12686
rect 19628 12226 19684 12236
rect 19516 11566 19518 11618
rect 19570 11566 19572 11618
rect 19516 11554 19572 11566
rect 19852 11396 19908 11406
rect 19852 11302 19908 11340
rect 19964 10610 20020 10622
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19852 9602 19908 9614
rect 19852 9550 19854 9602
rect 19906 9550 19908 9602
rect 19852 9492 19908 9550
rect 19852 9426 19908 9436
rect 19404 8372 19460 8382
rect 19404 8370 19908 8372
rect 19404 8318 19406 8370
rect 19458 8318 19908 8370
rect 19404 8316 19908 8318
rect 19404 8306 19460 8316
rect 19852 8258 19908 8316
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 19516 8148 19572 8158
rect 19572 8092 19684 8148
rect 19516 8054 19572 8092
rect 19516 7476 19572 7486
rect 19292 6972 19460 7028
rect 19292 6804 19348 6814
rect 19292 6578 19348 6748
rect 19292 6526 19294 6578
rect 19346 6526 19348 6578
rect 19292 6514 19348 6526
rect 19180 6066 19236 6076
rect 19292 6356 19348 6366
rect 19292 5906 19348 6300
rect 19404 6132 19460 6972
rect 19516 6690 19572 7420
rect 19628 7364 19684 8092
rect 19964 8036 20020 10558
rect 20188 9268 20244 17052
rect 27580 17108 27636 17118
rect 23772 16884 23828 16894
rect 20532 15708 20796 15718
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20532 15642 20796 15652
rect 23772 15148 23828 16828
rect 27356 15876 27412 15886
rect 23772 15092 24052 15148
rect 20532 14140 20796 14150
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20532 14074 20796 14084
rect 20860 12740 20916 12750
rect 21756 12740 21812 12750
rect 20860 12646 20916 12684
rect 21644 12738 21812 12740
rect 21644 12686 21758 12738
rect 21810 12686 21812 12738
rect 21644 12684 21812 12686
rect 20532 12572 20796 12582
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20532 12506 20796 12516
rect 20300 12292 20356 12302
rect 20300 12198 20356 12236
rect 20972 12178 21028 12190
rect 20972 12126 20974 12178
rect 21026 12126 21028 12178
rect 20972 12068 21028 12126
rect 21532 12068 21588 12078
rect 20972 12066 21588 12068
rect 20972 12014 21534 12066
rect 21586 12014 21588 12066
rect 20972 12012 21588 12014
rect 20636 11396 20692 11406
rect 20636 11394 20916 11396
rect 20636 11342 20638 11394
rect 20690 11342 20916 11394
rect 20636 11340 20916 11342
rect 20636 11330 20692 11340
rect 20412 11284 20468 11294
rect 20412 11190 20468 11228
rect 20532 11004 20796 11014
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20532 10938 20796 10948
rect 20300 10052 20356 10062
rect 20300 9938 20356 9996
rect 20300 9886 20302 9938
rect 20354 9886 20356 9938
rect 20300 9874 20356 9886
rect 20860 9828 20916 11340
rect 20972 10724 21028 12012
rect 21532 12002 21588 12012
rect 21644 11844 21700 12684
rect 21756 12674 21812 12684
rect 22540 12740 22596 12750
rect 22540 12402 22596 12684
rect 22876 12740 22932 12750
rect 23660 12740 23716 12750
rect 22876 12738 23044 12740
rect 22876 12686 22878 12738
rect 22930 12686 23044 12738
rect 22876 12684 23044 12686
rect 22876 12674 22932 12684
rect 22540 12350 22542 12402
rect 22594 12350 22596 12402
rect 22540 12338 22596 12350
rect 21308 11788 21700 11844
rect 22204 12066 22260 12078
rect 22204 12014 22206 12066
rect 22258 12014 22260 12066
rect 22204 11788 22260 12014
rect 22652 11844 22708 11854
rect 21084 10724 21140 10734
rect 20972 10722 21140 10724
rect 20972 10670 21086 10722
rect 21138 10670 21140 10722
rect 20972 10668 21140 10670
rect 20972 10052 21028 10668
rect 21084 10658 21140 10668
rect 21308 10164 21364 11788
rect 22204 11732 22372 11788
rect 21756 11508 21812 11518
rect 21420 11396 21476 11406
rect 21420 11172 21476 11340
rect 21420 11170 21588 11172
rect 21420 11118 21422 11170
rect 21474 11118 21588 11170
rect 21420 11116 21588 11118
rect 21420 11106 21476 11116
rect 21308 10098 21364 10108
rect 20972 9986 21028 9996
rect 21420 10052 21476 10062
rect 20860 9772 21364 9828
rect 20860 9604 20916 9614
rect 20860 9510 20916 9548
rect 20532 9436 20796 9446
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20532 9370 20796 9380
rect 19852 7980 20020 8036
rect 20076 9156 20132 9166
rect 19852 7700 19908 7980
rect 20076 7924 20132 9100
rect 20188 8258 20244 9212
rect 21196 8930 21252 8942
rect 21196 8878 21198 8930
rect 21250 8878 21252 8930
rect 21196 8484 21252 8878
rect 20300 8428 21252 8484
rect 20300 8370 20356 8428
rect 20300 8318 20302 8370
rect 20354 8318 20356 8370
rect 20300 8306 20356 8318
rect 21308 8372 21364 9772
rect 21420 9826 21476 9996
rect 21420 9774 21422 9826
rect 21474 9774 21476 9826
rect 21420 9762 21476 9774
rect 21532 8932 21588 11116
rect 21532 8866 21588 8876
rect 21644 8372 21700 8382
rect 21308 8316 21644 8372
rect 20188 8206 20190 8258
rect 20242 8206 20244 8258
rect 20188 8194 20244 8206
rect 20524 8260 20580 8270
rect 20524 8258 21252 8260
rect 20524 8206 20526 8258
rect 20578 8206 21252 8258
rect 20524 8204 21252 8206
rect 20524 8194 20580 8204
rect 19852 7634 19908 7644
rect 19964 7868 20132 7924
rect 21196 8148 21252 8204
rect 21644 8258 21700 8316
rect 21644 8206 21646 8258
rect 21698 8206 21700 8258
rect 21644 8194 21700 8206
rect 21308 8148 21364 8158
rect 21196 8146 21364 8148
rect 21196 8094 21310 8146
rect 21362 8094 21364 8146
rect 21196 8092 21364 8094
rect 20532 7868 20796 7878
rect 19628 7298 19684 7308
rect 19964 7252 20020 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20532 7802 20796 7812
rect 19740 7196 20020 7252
rect 20076 7364 20132 7374
rect 19516 6638 19518 6690
rect 19570 6638 19572 6690
rect 19516 6626 19572 6638
rect 19628 7140 19684 7150
rect 19516 6132 19572 6142
rect 19404 6130 19572 6132
rect 19404 6078 19518 6130
rect 19570 6078 19572 6130
rect 19404 6076 19572 6078
rect 19516 6066 19572 6076
rect 19292 5854 19294 5906
rect 19346 5854 19348 5906
rect 19292 5842 19348 5854
rect 18508 4620 18788 4676
rect 18844 4732 19012 4788
rect 18396 4564 18452 4574
rect 18284 4508 18396 4564
rect 18396 4498 18452 4508
rect 18172 3714 18228 3724
rect 16940 1026 16996 1036
rect 17052 1708 17220 1764
rect 17500 1820 17892 1876
rect 17948 3668 18004 3678
rect 17052 800 17108 1708
rect 17500 800 17556 1820
rect 17948 1764 18004 3612
rect 17724 1708 18004 1764
rect 18172 3556 18228 3566
rect 17724 800 17780 1708
rect 18172 800 18228 3500
rect 18396 3444 18452 3454
rect 18396 800 18452 3388
rect 18508 3388 18564 4620
rect 18732 4340 18788 4350
rect 18844 4340 18900 4732
rect 18732 4338 18900 4340
rect 18732 4286 18734 4338
rect 18786 4286 18900 4338
rect 18732 4284 18900 4286
rect 18732 4274 18788 4284
rect 18508 3332 18676 3388
rect 18620 2772 18676 3332
rect 18620 2706 18676 2716
rect 18844 800 18900 4284
rect 18956 4450 19012 4462
rect 18956 4398 18958 4450
rect 19010 4398 19012 4450
rect 18956 980 19012 4398
rect 19516 4116 19572 4126
rect 18956 914 19012 924
rect 19068 4114 19572 4116
rect 19068 4062 19518 4114
rect 19570 4062 19572 4114
rect 19068 4060 19572 4062
rect 19068 800 19124 4060
rect 19516 4050 19572 4060
rect 19628 3388 19684 7084
rect 19740 3554 19796 7196
rect 20076 6914 20132 7308
rect 20076 6862 20078 6914
rect 20130 6862 20132 6914
rect 20076 6850 20132 6862
rect 20412 6802 20468 6814
rect 20412 6750 20414 6802
rect 20466 6750 20468 6802
rect 20412 6692 20468 6750
rect 20412 6626 20468 6636
rect 20524 6804 20580 6814
rect 20300 6466 20356 6478
rect 20524 6468 20580 6748
rect 21196 6690 21252 8092
rect 21308 8082 21364 8092
rect 21644 8036 21700 8046
rect 21196 6638 21198 6690
rect 21250 6638 21252 6690
rect 21196 6468 21252 6638
rect 20300 6414 20302 6466
rect 20354 6414 20356 6466
rect 19852 5796 19908 5806
rect 20300 5796 20356 6414
rect 19852 5794 20356 5796
rect 19852 5742 19854 5794
rect 19906 5742 20356 5794
rect 19852 5740 20356 5742
rect 20412 6412 20580 6468
rect 20972 6412 21252 6468
rect 21308 7924 21364 7934
rect 19852 4900 19908 5740
rect 19964 5124 20020 5134
rect 19964 5030 20020 5068
rect 19852 4834 19908 4844
rect 19740 3502 19742 3554
rect 19794 3502 19796 3554
rect 19740 3490 19796 3502
rect 19628 3332 19796 3388
rect 19740 800 19796 3332
rect 20300 1428 20356 1438
rect 20300 1092 20356 1372
rect 20300 1026 20356 1036
rect 20412 800 20468 6412
rect 20532 6300 20796 6310
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20532 6234 20796 6244
rect 20748 5908 20804 5918
rect 20748 5122 20804 5852
rect 20748 5070 20750 5122
rect 20802 5070 20804 5122
rect 20748 5058 20804 5070
rect 20860 5124 20916 5134
rect 20972 5124 21028 6412
rect 21308 5572 21364 7868
rect 21532 7364 21588 7374
rect 21420 7308 21532 7364
rect 21420 5684 21476 7308
rect 21532 7298 21588 7308
rect 21644 6690 21700 7980
rect 21756 7924 21812 11452
rect 22204 11284 22260 11294
rect 22204 11190 22260 11228
rect 21868 11172 21924 11182
rect 21868 11170 22148 11172
rect 21868 11118 21870 11170
rect 21922 11118 22148 11170
rect 21868 11116 22148 11118
rect 21868 11106 21924 11116
rect 21980 10164 22036 10174
rect 21868 10052 21924 10062
rect 21868 9042 21924 9996
rect 21868 8990 21870 9042
rect 21922 8990 21924 9042
rect 21868 8978 21924 8990
rect 21756 7858 21812 7868
rect 21868 8260 21924 8270
rect 21756 7700 21812 7710
rect 21756 7474 21812 7644
rect 21756 7422 21758 7474
rect 21810 7422 21812 7474
rect 21756 7410 21812 7422
rect 21644 6638 21646 6690
rect 21698 6638 21700 6690
rect 21644 6626 21700 6638
rect 21756 6692 21812 6702
rect 21756 6598 21812 6636
rect 21532 6466 21588 6478
rect 21532 6414 21534 6466
rect 21586 6414 21588 6466
rect 21532 6132 21588 6414
rect 21868 6356 21924 8204
rect 21980 6916 22036 10108
rect 22092 9938 22148 11116
rect 22092 9886 22094 9938
rect 22146 9886 22148 9938
rect 22092 9874 22148 9886
rect 22316 11060 22372 11732
rect 22316 9716 22372 11004
rect 22092 9660 22372 9716
rect 22540 11284 22596 11294
rect 22092 8260 22148 9660
rect 22540 9266 22596 11228
rect 22540 9214 22542 9266
rect 22594 9214 22596 9266
rect 22540 9202 22596 9214
rect 22652 8932 22708 11788
rect 22764 11172 22820 11182
rect 22764 11078 22820 11116
rect 22876 10276 22932 10286
rect 22876 9828 22932 10220
rect 22092 8194 22148 8204
rect 22204 8876 22708 8932
rect 22764 9772 22932 9828
rect 21980 6580 22036 6860
rect 22092 8034 22148 8046
rect 22092 7982 22094 8034
rect 22146 7982 22148 8034
rect 22092 6804 22148 7982
rect 22092 6738 22148 6748
rect 21980 6524 22148 6580
rect 21868 6290 21924 6300
rect 21532 6076 22036 6132
rect 21980 6018 22036 6076
rect 21980 5966 21982 6018
rect 22034 5966 22036 6018
rect 21980 5954 22036 5966
rect 22092 5796 22148 6524
rect 21980 5740 22148 5796
rect 21420 5628 21812 5684
rect 21308 5516 21588 5572
rect 20916 5068 21028 5124
rect 21084 5460 21140 5470
rect 21084 5124 21140 5404
rect 21308 5348 21364 5358
rect 21308 5254 21364 5292
rect 21420 5124 21476 5134
rect 21084 5122 21476 5124
rect 21084 5070 21422 5122
rect 21474 5070 21476 5122
rect 21084 5068 21476 5070
rect 20860 5058 20916 5068
rect 21420 5058 21476 5068
rect 21084 4788 21140 4798
rect 20532 4732 20796 4742
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20532 4666 20796 4676
rect 20748 4564 20804 4574
rect 20748 3554 20804 4508
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 20532 3164 20796 3174
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20532 3098 20796 3108
rect 21084 800 21140 4732
rect 21532 4338 21588 5516
rect 21644 5236 21700 5246
rect 21644 5122 21700 5180
rect 21644 5070 21646 5122
rect 21698 5070 21700 5122
rect 21644 5058 21700 5070
rect 21532 4286 21534 4338
rect 21586 4286 21588 4338
rect 21532 4274 21588 4286
rect 21756 800 21812 5628
rect 21980 5122 22036 5740
rect 22204 5236 22260 8876
rect 22316 8708 22372 8718
rect 22316 6356 22372 8652
rect 22764 8484 22820 9772
rect 22876 9604 22932 9614
rect 22876 8818 22932 9548
rect 22876 8766 22878 8818
rect 22930 8766 22932 8818
rect 22876 8708 22932 8766
rect 22876 8642 22932 8652
rect 22316 6290 22372 6300
rect 22428 8428 22820 8484
rect 21980 5070 21982 5122
rect 22034 5070 22036 5122
rect 21980 5058 22036 5070
rect 22092 5180 22260 5236
rect 22428 5236 22484 8428
rect 22764 8260 22820 8270
rect 22988 8260 23044 12684
rect 23660 12738 23828 12740
rect 23660 12686 23662 12738
rect 23714 12686 23828 12738
rect 23660 12684 23828 12686
rect 23660 12674 23716 12684
rect 23548 12290 23604 12302
rect 23548 12238 23550 12290
rect 23602 12238 23604 12290
rect 23100 12068 23156 12078
rect 23100 12066 23268 12068
rect 23100 12014 23102 12066
rect 23154 12014 23268 12066
rect 23100 12012 23268 12014
rect 23100 12002 23156 12012
rect 23100 11172 23156 11182
rect 23100 10052 23156 11116
rect 23100 9986 23156 9996
rect 22092 4452 22148 5180
rect 22428 5170 22484 5180
rect 22540 8090 22596 8102
rect 22540 8038 22542 8090
rect 22594 8038 22596 8090
rect 22316 5124 22372 5134
rect 22316 5030 22372 5068
rect 22204 5012 22260 5022
rect 22204 4918 22260 4956
rect 22540 4676 22596 8038
rect 22652 6466 22708 6478
rect 22652 6414 22654 6466
rect 22706 6414 22708 6466
rect 22652 5124 22708 6414
rect 22764 5908 22820 8204
rect 22876 8204 23044 8260
rect 23100 9156 23156 9166
rect 22876 7588 22932 8204
rect 22876 7140 22932 7532
rect 22988 8034 23044 8046
rect 22988 7982 22990 8034
rect 23042 7982 23044 8034
rect 22988 7364 23044 7982
rect 22988 7298 23044 7308
rect 22876 7074 22932 7084
rect 23100 6804 23156 9100
rect 23212 7812 23268 12012
rect 23436 11508 23492 11518
rect 23548 11508 23604 12238
rect 23492 11452 23604 11508
rect 23660 12178 23716 12190
rect 23660 12126 23662 12178
rect 23714 12126 23716 12178
rect 23436 11414 23492 11452
rect 23324 11284 23380 11294
rect 23324 10052 23380 11228
rect 23324 9996 23604 10052
rect 23436 9268 23492 9278
rect 23436 9154 23492 9212
rect 23436 9102 23438 9154
rect 23490 9102 23492 9154
rect 23436 9090 23492 9102
rect 23548 9044 23604 9996
rect 23548 8258 23604 8988
rect 23660 9042 23716 12126
rect 23660 8990 23662 9042
rect 23714 8990 23716 9042
rect 23660 8372 23716 8990
rect 23660 8306 23716 8316
rect 23772 9716 23828 12684
rect 23548 8206 23550 8258
rect 23602 8206 23604 8258
rect 23548 8194 23604 8206
rect 23212 7756 23492 7812
rect 22764 5814 22820 5852
rect 22876 6748 23156 6804
rect 23212 7140 23268 7150
rect 22764 5348 22820 5358
rect 22764 5254 22820 5292
rect 22876 5236 22932 6748
rect 22988 6580 23044 6618
rect 22988 6514 23044 6524
rect 23100 6466 23156 6478
rect 23100 6414 23102 6466
rect 23154 6414 23156 6466
rect 22988 6356 23044 6366
rect 22988 5796 23044 6300
rect 23100 6132 23156 6414
rect 23100 6066 23156 6076
rect 23212 6018 23268 7084
rect 23436 6580 23492 7756
rect 23660 7586 23716 7598
rect 23660 7534 23662 7586
rect 23714 7534 23716 7586
rect 23436 6514 23492 6524
rect 23548 6690 23604 6702
rect 23548 6638 23550 6690
rect 23602 6638 23604 6690
rect 23324 6468 23380 6478
rect 23324 6374 23380 6412
rect 23212 5966 23214 6018
rect 23266 5966 23268 6018
rect 23212 5954 23268 5966
rect 23324 5906 23380 5918
rect 23324 5854 23326 5906
rect 23378 5854 23380 5906
rect 22988 5740 23156 5796
rect 22876 5180 23044 5236
rect 22652 5068 22932 5124
rect 22876 4900 22932 5068
rect 22876 4834 22932 4844
rect 22428 4620 22596 4676
rect 22204 4452 22260 4462
rect 22148 4450 22260 4452
rect 22148 4398 22206 4450
rect 22258 4398 22260 4450
rect 22148 4396 22260 4398
rect 22092 4358 22148 4396
rect 22204 4386 22260 4396
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 22428 800 22484 4620
rect 22540 4450 22596 4462
rect 22540 4398 22542 4450
rect 22594 4398 22596 4450
rect 22540 3556 22596 4398
rect 22540 3490 22596 3500
rect 22988 3388 23044 5180
rect 23100 5122 23156 5740
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 23100 5058 23156 5070
rect 23324 5012 23380 5854
rect 23324 4564 23380 4956
rect 23324 4450 23380 4508
rect 23324 4398 23326 4450
rect 23378 4398 23380 4450
rect 23324 4386 23380 4398
rect 23436 5906 23492 5918
rect 23436 5854 23438 5906
rect 23490 5854 23492 5906
rect 23436 5124 23492 5854
rect 23548 5572 23604 6638
rect 23660 5796 23716 7534
rect 23660 5730 23716 5740
rect 23548 5506 23604 5516
rect 23772 5236 23828 9660
rect 23884 8372 23940 8382
rect 23884 8278 23940 8316
rect 23884 7588 23940 7598
rect 23884 6020 23940 7532
rect 23996 7140 24052 15092
rect 24108 12740 24164 12750
rect 24164 12684 24388 12740
rect 24108 12646 24164 12684
rect 24220 12404 24276 12414
rect 24220 12178 24276 12348
rect 24220 12126 24222 12178
rect 24274 12126 24276 12178
rect 24220 12114 24276 12126
rect 24220 9938 24276 9950
rect 24220 9886 24222 9938
rect 24274 9886 24276 9938
rect 24220 9268 24276 9886
rect 24220 9202 24276 9212
rect 24108 9156 24164 9166
rect 24108 9062 24164 9100
rect 24220 8932 24276 8942
rect 24108 8148 24164 8158
rect 24108 7476 24164 8092
rect 24220 7588 24276 8876
rect 24332 8260 24388 12684
rect 24444 12738 24500 12750
rect 25004 12740 25060 12750
rect 24444 12686 24446 12738
rect 24498 12686 24500 12738
rect 24444 11172 24500 12686
rect 24780 12684 25004 12740
rect 24444 11106 24500 11116
rect 24556 11954 24612 11966
rect 24556 11902 24558 11954
rect 24610 11902 24612 11954
rect 24556 10724 24612 11902
rect 24556 10658 24612 10668
rect 24332 8166 24388 8204
rect 24444 10052 24500 10062
rect 24444 9828 24500 9996
rect 24220 7522 24276 7532
rect 24332 7924 24388 7934
rect 24108 7382 24164 7420
rect 23996 7074 24052 7084
rect 23884 5954 23940 5964
rect 24220 6916 24276 6926
rect 24108 5796 24164 5806
rect 23884 5684 23940 5694
rect 23884 5682 24052 5684
rect 23884 5630 23886 5682
rect 23938 5630 24052 5682
rect 23884 5628 24052 5630
rect 23884 5618 23940 5628
rect 23436 4450 23492 5068
rect 23436 4398 23438 4450
rect 23490 4398 23492 4450
rect 23436 4386 23492 4398
rect 23548 5180 23828 5236
rect 23100 4340 23156 4350
rect 23100 4246 23156 4284
rect 23548 3556 23604 5180
rect 23772 4900 23828 4910
rect 23660 3556 23716 3566
rect 23548 3554 23716 3556
rect 23548 3502 23662 3554
rect 23714 3502 23716 3554
rect 23548 3500 23716 3502
rect 23660 3490 23716 3500
rect 22988 3332 23156 3388
rect 23100 800 23156 3332
rect 23772 800 23828 4844
rect 23884 4898 23940 4910
rect 23884 4846 23886 4898
rect 23938 4846 23940 4898
rect 23884 4340 23940 4846
rect 23884 4274 23940 4284
rect 23884 4116 23940 4126
rect 23884 4022 23940 4060
rect 23996 3780 24052 5628
rect 24108 4788 24164 5740
rect 24220 5684 24276 6860
rect 24332 6132 24388 7868
rect 24444 7028 24500 9772
rect 24556 9154 24612 9166
rect 24556 9102 24558 9154
rect 24610 9102 24612 9154
rect 24556 7252 24612 9102
rect 24668 8260 24724 8270
rect 24668 7698 24724 8204
rect 24668 7646 24670 7698
rect 24722 7646 24724 7698
rect 24668 7634 24724 7646
rect 24556 7186 24612 7196
rect 24444 6972 24612 7028
rect 24556 6916 24612 6972
rect 24556 6850 24612 6860
rect 24332 6038 24388 6076
rect 24444 6804 24500 6814
rect 24780 6804 24836 12684
rect 25004 12646 25060 12684
rect 25340 12738 25396 12750
rect 25340 12686 25342 12738
rect 25394 12686 25396 12738
rect 25340 11844 25396 12686
rect 25900 12740 25956 12750
rect 26684 12740 26740 12750
rect 25900 12646 25956 12684
rect 26348 12738 26740 12740
rect 26348 12686 26686 12738
rect 26738 12686 26740 12738
rect 26348 12684 26740 12686
rect 25452 12404 25508 12414
rect 25452 12310 25508 12348
rect 25340 11778 25396 11788
rect 25788 12066 25844 12078
rect 25788 12014 25790 12066
rect 25842 12014 25844 12066
rect 25788 11956 25844 12014
rect 26236 12068 26292 12078
rect 26236 11974 26292 12012
rect 25564 11282 25620 11294
rect 25564 11230 25566 11282
rect 25618 11230 25620 11282
rect 25564 10834 25620 11230
rect 25564 10782 25566 10834
rect 25618 10782 25620 10834
rect 25564 10770 25620 10782
rect 25228 10724 25284 10734
rect 25228 10630 25284 10668
rect 25788 10276 25844 11900
rect 26124 11508 26180 11518
rect 26012 11452 26124 11508
rect 25788 10210 25844 10220
rect 25900 10722 25956 10734
rect 25900 10670 25902 10722
rect 25954 10670 25956 10722
rect 25228 10164 25284 10174
rect 24220 5618 24276 5628
rect 24332 5124 24388 5134
rect 24332 5010 24388 5068
rect 24332 4958 24334 5010
rect 24386 4958 24388 5010
rect 24332 4946 24388 4958
rect 24108 4722 24164 4732
rect 24220 4564 24276 4574
rect 24220 4470 24276 4508
rect 23996 3714 24052 3724
rect 24108 4228 24164 4238
rect 23996 3444 24052 3454
rect 24108 3444 24164 4172
rect 23996 3442 24164 3444
rect 23996 3390 23998 3442
rect 24050 3390 24164 3442
rect 23996 3388 24164 3390
rect 23996 3378 24052 3388
rect 24444 800 24500 6748
rect 24668 6748 24836 6804
rect 24892 9602 24948 9614
rect 24892 9550 24894 9602
rect 24946 9550 24948 9602
rect 24556 6690 24612 6702
rect 24556 6638 24558 6690
rect 24610 6638 24612 6690
rect 24556 4564 24612 6638
rect 24668 6356 24724 6748
rect 24668 6290 24724 6300
rect 24780 6578 24836 6590
rect 24780 6526 24782 6578
rect 24834 6526 24836 6578
rect 24668 5908 24724 5918
rect 24668 5814 24724 5852
rect 24668 5684 24724 5694
rect 24668 5124 24724 5628
rect 24780 5348 24836 6526
rect 24780 5282 24836 5292
rect 24668 5122 24836 5124
rect 24668 5070 24670 5122
rect 24722 5070 24836 5122
rect 24668 5068 24836 5070
rect 24668 5058 24724 5068
rect 24556 4508 24724 4564
rect 24556 4338 24612 4350
rect 24556 4286 24558 4338
rect 24610 4286 24612 4338
rect 24556 3780 24612 4286
rect 24668 4228 24724 4508
rect 24668 4162 24724 4172
rect 24780 4004 24836 5068
rect 24892 4788 24948 9550
rect 25004 8484 25060 8494
rect 25004 6692 25060 8428
rect 25116 8372 25172 8382
rect 25116 8278 25172 8316
rect 25228 6804 25284 10108
rect 25900 10164 25956 10670
rect 25900 10098 25956 10108
rect 25340 9602 25396 9614
rect 25340 9550 25342 9602
rect 25394 9550 25396 9602
rect 25340 9268 25396 9550
rect 25788 9604 25844 9614
rect 25788 9510 25844 9548
rect 26012 9492 26068 11452
rect 26124 11442 26180 11452
rect 26236 11394 26292 11406
rect 26236 11342 26238 11394
rect 26290 11342 26292 11394
rect 26236 11172 26292 11342
rect 26236 10500 26292 11116
rect 26236 10434 26292 10444
rect 25340 9202 25396 9212
rect 25900 9436 26068 9492
rect 25676 9156 25732 9166
rect 25564 8818 25620 8830
rect 25564 8766 25566 8818
rect 25618 8766 25620 8818
rect 25228 6738 25284 6748
rect 25340 7586 25396 7598
rect 25340 7534 25342 7586
rect 25394 7534 25396 7586
rect 25116 6692 25172 6702
rect 25004 6690 25172 6692
rect 25004 6638 25118 6690
rect 25170 6638 25172 6690
rect 25004 6636 25172 6638
rect 25116 6626 25172 6636
rect 25116 6356 25172 6366
rect 25004 6244 25060 6254
rect 25004 5122 25060 6188
rect 25004 5070 25006 5122
rect 25058 5070 25060 5122
rect 25004 5058 25060 5070
rect 25116 5684 25172 6300
rect 25340 6356 25396 7534
rect 25564 7140 25620 8766
rect 25676 7474 25732 9100
rect 25900 9044 25956 9436
rect 26348 9380 26404 12684
rect 26684 12674 26740 12684
rect 27132 12738 27188 12750
rect 27132 12686 27134 12738
rect 27186 12686 27188 12738
rect 26684 12066 26740 12078
rect 26684 12014 26686 12066
rect 26738 12014 26740 12066
rect 26684 11956 26740 12014
rect 26684 11890 26740 11900
rect 26796 12068 26852 12078
rect 26796 11170 26852 12012
rect 27132 11788 27188 12686
rect 27356 12402 27412 15820
rect 27580 12740 27636 17052
rect 28812 16996 28868 17006
rect 27356 12350 27358 12402
rect 27410 12350 27412 12402
rect 27356 12338 27412 12350
rect 27468 12738 27636 12740
rect 27468 12686 27582 12738
rect 27634 12686 27636 12738
rect 27468 12684 27636 12686
rect 27132 11732 27412 11788
rect 27244 11172 27300 11182
rect 26796 11118 26798 11170
rect 26850 11118 26852 11170
rect 26796 10500 26852 11118
rect 26684 10498 26852 10500
rect 26684 10446 26798 10498
rect 26850 10446 26852 10498
rect 26684 10444 26852 10446
rect 26460 10276 26516 10286
rect 26516 10220 26628 10276
rect 26460 10210 26516 10220
rect 26236 9324 26404 9380
rect 26460 9714 26516 9726
rect 26460 9662 26462 9714
rect 26514 9662 26516 9714
rect 26012 9268 26068 9278
rect 26068 9212 26180 9268
rect 26012 9202 26068 9212
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 7410 25732 7422
rect 25788 8988 25956 9044
rect 25788 7252 25844 8988
rect 25900 8820 25956 8830
rect 25900 8818 26068 8820
rect 25900 8766 25902 8818
rect 25954 8766 26068 8818
rect 25900 8764 26068 8766
rect 25900 8754 25956 8764
rect 25900 7588 25956 7598
rect 25900 7494 25956 7532
rect 26012 7476 26068 8764
rect 26012 7410 26068 7420
rect 25564 7074 25620 7084
rect 25676 7196 25844 7252
rect 25900 7252 25956 7262
rect 25676 6916 25732 7196
rect 25900 7140 25956 7196
rect 25564 6860 25732 6916
rect 25788 7084 25956 7140
rect 26012 7250 26068 7262
rect 26012 7198 26014 7250
rect 26066 7198 26068 7250
rect 25564 6578 25620 6860
rect 25564 6526 25566 6578
rect 25618 6526 25620 6578
rect 25564 6514 25620 6526
rect 25676 6690 25732 6702
rect 25676 6638 25678 6690
rect 25730 6638 25732 6690
rect 25340 6290 25396 6300
rect 25676 6356 25732 6638
rect 25676 6290 25732 6300
rect 24892 4722 24948 4732
rect 25116 4004 25172 5628
rect 24780 3938 24836 3948
rect 25004 3948 25172 4004
rect 25228 6132 25284 6142
rect 25228 5122 25284 6076
rect 25340 6018 25396 6030
rect 25340 5966 25342 6018
rect 25394 5966 25396 6018
rect 25340 5684 25396 5966
rect 25676 5908 25732 5918
rect 25564 5906 25732 5908
rect 25564 5854 25678 5906
rect 25730 5854 25732 5906
rect 25564 5852 25732 5854
rect 25340 5628 25508 5684
rect 25228 5070 25230 5122
rect 25282 5070 25284 5122
rect 25004 3780 25060 3948
rect 24556 3724 25060 3780
rect 24892 3556 24948 3566
rect 24668 3444 24724 3454
rect 24668 3330 24724 3388
rect 24668 3278 24670 3330
rect 24722 3278 24724 3330
rect 24668 3266 24724 3278
rect 24892 1316 24948 3500
rect 25004 3554 25060 3724
rect 25004 3502 25006 3554
rect 25058 3502 25060 3554
rect 25004 3490 25060 3502
rect 25116 3668 25172 3678
rect 24892 1250 24948 1260
rect 25116 800 25172 3612
rect 25228 3444 25284 5070
rect 25340 5460 25396 5470
rect 25340 5122 25396 5404
rect 25340 5070 25342 5122
rect 25394 5070 25396 5122
rect 25340 5058 25396 5070
rect 25340 3444 25396 3454
rect 25228 3442 25396 3444
rect 25228 3390 25342 3442
rect 25394 3390 25396 3442
rect 25228 3388 25396 3390
rect 25340 3378 25396 3388
rect 25452 2994 25508 5628
rect 25564 3554 25620 5852
rect 25676 5842 25732 5852
rect 25788 5346 25844 7084
rect 25900 6468 25956 6478
rect 25900 5906 25956 6412
rect 25900 5854 25902 5906
rect 25954 5854 25956 5906
rect 25900 5842 25956 5854
rect 25788 5294 25790 5346
rect 25842 5294 25844 5346
rect 25788 5282 25844 5294
rect 26012 5012 26068 7198
rect 26012 4946 26068 4956
rect 25788 4788 25844 4798
rect 25564 3502 25566 3554
rect 25618 3502 25620 3554
rect 25564 3490 25620 3502
rect 25676 4226 25732 4238
rect 25676 4174 25678 4226
rect 25730 4174 25732 4226
rect 25452 2942 25454 2994
rect 25506 2942 25508 2994
rect 25452 2930 25508 2942
rect 25676 2548 25732 4174
rect 25676 2482 25732 2492
rect 25788 800 25844 4732
rect 26124 4564 26180 9212
rect 26012 4508 26180 4564
rect 25900 4452 25956 4462
rect 25900 4358 25956 4396
rect 25900 4228 25956 4238
rect 25900 3556 25956 4172
rect 25900 3490 25956 3500
rect 26012 3388 26068 4508
rect 26124 4338 26180 4350
rect 26124 4286 26126 4338
rect 26178 4286 26180 4338
rect 26124 4228 26180 4286
rect 26124 4162 26180 4172
rect 26124 3780 26180 3790
rect 26124 3686 26180 3724
rect 26236 3444 26292 9324
rect 26460 9266 26516 9662
rect 26460 9214 26462 9266
rect 26514 9214 26516 9266
rect 26460 9202 26516 9214
rect 26348 9156 26404 9166
rect 26348 9062 26404 9100
rect 26572 9044 26628 10220
rect 26684 9156 26740 10444
rect 26796 10434 26852 10444
rect 27132 11116 27244 11172
rect 27132 10276 27188 11116
rect 27244 11078 27300 11116
rect 26684 9090 26740 9100
rect 26796 10220 27188 10276
rect 27244 10500 27300 10510
rect 26460 8988 26628 9044
rect 26460 8932 26516 8988
rect 26348 8876 26516 8932
rect 26348 7700 26404 8876
rect 26572 8820 26628 8830
rect 26572 8818 26740 8820
rect 26572 8766 26574 8818
rect 26626 8766 26740 8818
rect 26572 8764 26740 8766
rect 26572 8754 26628 8764
rect 26348 7586 26404 7644
rect 26348 7534 26350 7586
rect 26402 7534 26404 7586
rect 26348 7522 26404 7534
rect 26572 7700 26628 7710
rect 26572 7474 26628 7644
rect 26572 7422 26574 7474
rect 26626 7422 26628 7474
rect 26460 7364 26516 7374
rect 26460 6914 26516 7308
rect 26460 6862 26462 6914
rect 26514 6862 26516 6914
rect 26460 6850 26516 6862
rect 26572 6692 26628 7422
rect 26572 6626 26628 6636
rect 26460 6468 26516 6478
rect 26348 6466 26516 6468
rect 26348 6414 26462 6466
rect 26514 6414 26516 6466
rect 26348 6412 26516 6414
rect 26348 5124 26404 6412
rect 26460 6402 26516 6412
rect 26572 6466 26628 6478
rect 26572 6414 26574 6466
rect 26626 6414 26628 6466
rect 26572 5906 26628 6414
rect 26572 5854 26574 5906
rect 26626 5854 26628 5906
rect 26572 5842 26628 5854
rect 26572 5572 26628 5582
rect 26348 5068 26516 5124
rect 26348 4900 26404 4910
rect 26348 4806 26404 4844
rect 26348 4340 26404 4350
rect 26348 4246 26404 4284
rect 26460 3668 26516 5068
rect 26572 4338 26628 5516
rect 26684 5236 26740 8764
rect 26796 8148 26852 10220
rect 26796 8082 26852 8092
rect 26908 9940 26964 9950
rect 26796 7924 26852 7934
rect 26796 7698 26852 7868
rect 26796 7646 26798 7698
rect 26850 7646 26852 7698
rect 26796 7634 26852 7646
rect 26796 7362 26852 7374
rect 26796 7310 26798 7362
rect 26850 7310 26852 7362
rect 26796 6692 26852 7310
rect 26908 6802 26964 9884
rect 27020 9044 27076 9054
rect 27244 9044 27300 10444
rect 27020 9042 27300 9044
rect 27020 8990 27022 9042
rect 27074 8990 27300 9042
rect 27020 8988 27300 8990
rect 27020 8978 27076 8988
rect 27132 8372 27188 8382
rect 27020 8148 27076 8158
rect 27020 7700 27076 8092
rect 27020 7634 27076 7644
rect 26908 6750 26910 6802
rect 26962 6750 26964 6802
rect 26908 6738 26964 6750
rect 27132 6802 27188 8316
rect 27244 8370 27300 8382
rect 27244 8318 27246 8370
rect 27298 8318 27300 8370
rect 27244 8260 27300 8318
rect 27244 7812 27300 8204
rect 27244 7746 27300 7756
rect 27244 7588 27300 7598
rect 27244 7494 27300 7532
rect 27356 7252 27412 11732
rect 27468 8820 27524 12684
rect 27580 12674 27636 12684
rect 28252 15652 28308 15662
rect 27916 12066 27972 12078
rect 27916 12014 27918 12066
rect 27970 12014 27972 12066
rect 27804 11170 27860 11182
rect 27804 11118 27806 11170
rect 27858 11118 27860 11170
rect 27804 10724 27860 11118
rect 27804 10658 27860 10668
rect 27692 10500 27748 10510
rect 27692 10498 27860 10500
rect 27692 10446 27694 10498
rect 27746 10446 27860 10498
rect 27692 10444 27860 10446
rect 27692 10434 27748 10444
rect 27580 9940 27636 9950
rect 27580 9846 27636 9884
rect 27692 8930 27748 8942
rect 27692 8878 27694 8930
rect 27746 8878 27748 8930
rect 27468 8764 27636 8820
rect 27356 7028 27412 7196
rect 27580 7252 27636 8764
rect 27692 8260 27748 8878
rect 27692 8194 27748 8204
rect 27692 8036 27748 8046
rect 27804 8036 27860 10444
rect 27916 10052 27972 12014
rect 28252 11508 28308 15596
rect 28252 11414 28308 11452
rect 28364 12066 28420 12078
rect 28364 12014 28366 12066
rect 28418 12014 28420 12066
rect 28028 10498 28084 10510
rect 28028 10446 28030 10498
rect 28082 10446 28084 10498
rect 28028 10164 28084 10446
rect 28028 10098 28084 10108
rect 27916 9986 27972 9996
rect 28140 9828 28196 9838
rect 28140 9734 28196 9772
rect 28364 8484 28420 12014
rect 28812 12066 28868 16940
rect 30192 16492 30456 16502
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30192 16426 30456 16436
rect 31836 15876 31892 15886
rect 31276 15540 31332 15550
rect 31276 15148 31332 15484
rect 31836 15148 31892 15820
rect 31948 15764 32004 15774
rect 31948 15540 32004 15708
rect 32508 15652 32564 15662
rect 31948 15474 32004 15484
rect 32396 15596 32508 15652
rect 30716 15092 31332 15148
rect 31388 15092 31892 15148
rect 30192 14924 30456 14934
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30192 14858 30456 14868
rect 28812 12014 28814 12066
rect 28866 12014 28868 12066
rect 28588 11172 28644 11182
rect 28588 11078 28644 11116
rect 28700 10052 28756 10062
rect 28700 9938 28756 9996
rect 28700 9886 28702 9938
rect 28754 9886 28756 9938
rect 28700 9874 28756 9886
rect 28252 8428 28420 8484
rect 28700 9268 28756 9278
rect 27916 8372 27972 8382
rect 27916 8258 27972 8316
rect 27916 8206 27918 8258
rect 27970 8206 27972 8258
rect 27916 8194 27972 8206
rect 27748 7980 27860 8036
rect 28028 8146 28084 8158
rect 28028 8094 28030 8146
rect 28082 8094 28084 8146
rect 27692 7970 27748 7980
rect 28028 7588 28084 8094
rect 27804 7532 28084 7588
rect 28140 8148 28196 8158
rect 27580 7186 27636 7196
rect 27692 7476 27748 7486
rect 27356 6972 27636 7028
rect 27132 6750 27134 6802
rect 27186 6750 27188 6802
rect 27132 6738 27188 6750
rect 26796 6626 26852 6636
rect 26908 6468 26964 6478
rect 26796 6356 26852 6366
rect 26796 5796 26852 6300
rect 26796 5730 26852 5740
rect 26684 5170 26740 5180
rect 26908 5234 26964 6412
rect 27356 6356 27412 6366
rect 27356 6020 27412 6300
rect 27468 6020 27524 6030
rect 27356 6018 27524 6020
rect 27356 5966 27470 6018
rect 27522 5966 27524 6018
rect 27356 5964 27524 5966
rect 27468 5954 27524 5964
rect 27356 5682 27412 5694
rect 27356 5630 27358 5682
rect 27410 5630 27412 5682
rect 26908 5182 26910 5234
rect 26962 5182 26964 5234
rect 26908 5170 26964 5182
rect 27244 5236 27300 5246
rect 26796 4900 26852 4910
rect 26796 4450 26852 4844
rect 26796 4398 26798 4450
rect 26850 4398 26852 4450
rect 26796 4386 26852 4398
rect 26908 4676 26964 4686
rect 26572 4286 26574 4338
rect 26626 4286 26628 4338
rect 26572 4274 26628 4286
rect 26684 4228 26740 4238
rect 26684 4134 26740 4172
rect 26460 3602 26516 3612
rect 26572 4004 26628 4014
rect 26348 3554 26404 3566
rect 26348 3502 26350 3554
rect 26402 3502 26404 3554
rect 26348 3444 26404 3502
rect 26572 3554 26628 3948
rect 26572 3502 26574 3554
rect 26626 3502 26628 3554
rect 26572 3490 26628 3502
rect 26908 3554 26964 4620
rect 27244 4226 27300 5180
rect 27356 5234 27412 5630
rect 27580 5572 27636 6972
rect 27692 5906 27748 7420
rect 27804 6692 27860 7532
rect 28140 7364 28196 8092
rect 28028 7308 28196 7364
rect 27804 6626 27860 6636
rect 27916 7252 27972 7262
rect 27804 6020 27860 6030
rect 27804 5926 27860 5964
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 27692 5842 27748 5854
rect 27916 5572 27972 7196
rect 28028 6916 28084 7308
rect 28028 6850 28084 6860
rect 28140 7140 28196 7150
rect 28028 6692 28084 6702
rect 28028 6132 28084 6636
rect 28140 6578 28196 7084
rect 28140 6526 28142 6578
rect 28194 6526 28196 6578
rect 28140 6514 28196 6526
rect 28028 6066 28084 6076
rect 27580 5506 27636 5516
rect 27692 5516 27972 5572
rect 28140 5794 28196 5806
rect 28140 5742 28142 5794
rect 28194 5742 28196 5794
rect 27356 5182 27358 5234
rect 27410 5182 27412 5234
rect 27356 5170 27412 5182
rect 27692 4788 27748 5516
rect 27804 5348 27860 5358
rect 28140 5348 28196 5742
rect 27860 5292 28196 5348
rect 27804 5282 27860 5292
rect 28252 5236 28308 8428
rect 28364 8260 28420 8270
rect 28364 7362 28420 8204
rect 28364 7310 28366 7362
rect 28418 7310 28420 7362
rect 28364 7298 28420 7310
rect 28588 8034 28644 8046
rect 28588 7982 28590 8034
rect 28642 7982 28644 8034
rect 28476 7140 28532 7150
rect 27244 4174 27246 4226
rect 27298 4174 27300 4226
rect 27244 4162 27300 4174
rect 27580 4732 27748 4788
rect 28028 5180 28308 5236
rect 28364 6916 28420 6926
rect 28364 5460 28420 6860
rect 28476 6468 28532 7084
rect 28588 6916 28644 7982
rect 28588 6850 28644 6860
rect 28476 6412 28644 6468
rect 28588 6356 28644 6412
rect 28588 6290 28644 6300
rect 27356 4116 27412 4126
rect 27356 3778 27412 4060
rect 27580 4004 27636 4732
rect 27692 4564 27748 4602
rect 27692 4498 27748 4508
rect 27580 3938 27636 3948
rect 27692 4340 27748 4350
rect 27356 3726 27358 3778
rect 27410 3726 27412 3778
rect 27356 3714 27412 3726
rect 27580 3668 27636 3678
rect 27580 3574 27636 3612
rect 26908 3502 26910 3554
rect 26962 3502 26964 3554
rect 26908 3490 26964 3502
rect 27132 3556 27188 3566
rect 27132 3462 27188 3500
rect 26236 3388 26404 3444
rect 25900 3332 26068 3388
rect 25900 980 25956 3332
rect 26348 2324 26404 3388
rect 26684 3332 26740 3342
rect 26684 3238 26740 3276
rect 26348 2258 26404 2268
rect 27692 1316 27748 4284
rect 27804 3556 27860 3566
rect 28028 3556 28084 5180
rect 28140 5012 28196 5022
rect 28140 4226 28196 4956
rect 28140 4174 28142 4226
rect 28194 4174 28196 4226
rect 28140 4162 28196 4174
rect 28252 5010 28308 5022
rect 28252 4958 28254 5010
rect 28306 4958 28308 5010
rect 27804 3554 28084 3556
rect 27804 3502 27806 3554
rect 27858 3502 28084 3554
rect 27804 3500 28084 3502
rect 27804 3490 27860 3500
rect 27916 3330 27972 3342
rect 27916 3278 27918 3330
rect 27970 3278 27972 3330
rect 27916 3220 27972 3278
rect 27916 3154 27972 3164
rect 27692 1260 27860 1316
rect 27132 980 27188 990
rect 25900 924 26516 980
rect 26460 800 26516 924
rect 27132 800 27188 924
rect 27804 800 27860 1260
rect 28028 980 28084 3500
rect 28252 3332 28308 4958
rect 28364 3442 28420 5404
rect 28364 3390 28366 3442
rect 28418 3390 28420 3442
rect 28364 3378 28420 3390
rect 28476 6244 28532 6254
rect 28252 3266 28308 3276
rect 28028 914 28084 924
rect 28476 800 28532 6188
rect 28700 4340 28756 9212
rect 28700 4274 28756 4284
rect 28588 3892 28644 3902
rect 28588 3554 28644 3836
rect 28812 3668 28868 12014
rect 28924 13748 28980 13758
rect 28924 8372 28980 13692
rect 30192 13356 30456 13366
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30192 13290 30456 13300
rect 30492 12738 30548 12750
rect 30492 12686 30494 12738
rect 30546 12686 30548 12738
rect 29372 12290 29428 12302
rect 29372 12238 29374 12290
rect 29426 12238 29428 12290
rect 29372 11506 29428 12238
rect 29372 11454 29374 11506
rect 29426 11454 29428 11506
rect 29372 11442 29428 11454
rect 30044 12292 30100 12302
rect 29484 11282 29540 11294
rect 29484 11230 29486 11282
rect 29538 11230 29540 11282
rect 29260 11172 29316 11182
rect 29260 11078 29316 11116
rect 29148 10836 29204 10846
rect 28924 8306 28980 8316
rect 29036 8596 29092 8606
rect 28924 7812 28980 7822
rect 28924 4228 28980 7756
rect 29036 7140 29092 8540
rect 29148 7700 29204 10780
rect 29260 10500 29316 10510
rect 29260 9826 29316 10444
rect 29260 9774 29262 9826
rect 29314 9774 29316 9826
rect 29260 9762 29316 9774
rect 29484 8820 29540 11230
rect 29932 11284 29988 11294
rect 29932 11170 29988 11228
rect 29932 11118 29934 11170
rect 29986 11118 29988 11170
rect 29932 10836 29988 11118
rect 29484 8754 29540 8764
rect 29596 10780 29988 10836
rect 29596 9268 29652 10780
rect 29820 10612 29876 10622
rect 29820 10164 29876 10556
rect 29820 9716 29876 10108
rect 29932 9940 29988 9950
rect 29932 9846 29988 9884
rect 29820 9660 29988 9716
rect 29596 8596 29652 9212
rect 29820 8932 29876 8942
rect 29820 8838 29876 8876
rect 29596 8530 29652 8540
rect 29708 8708 29764 8718
rect 29484 7924 29540 7934
rect 29260 7700 29316 7710
rect 29148 7698 29316 7700
rect 29148 7646 29262 7698
rect 29314 7646 29316 7698
rect 29148 7644 29316 7646
rect 29036 7074 29092 7084
rect 29148 6580 29204 6590
rect 29036 6578 29204 6580
rect 29036 6526 29150 6578
rect 29202 6526 29204 6578
rect 29036 6524 29204 6526
rect 29036 4452 29092 6524
rect 29148 6514 29204 6524
rect 29260 6468 29316 7644
rect 29372 6804 29428 6842
rect 29372 6738 29428 6748
rect 29260 6402 29316 6412
rect 29372 6580 29428 6590
rect 29372 6244 29428 6524
rect 29260 6188 29428 6244
rect 29260 5236 29316 6188
rect 29260 5122 29316 5180
rect 29260 5070 29262 5122
rect 29314 5070 29316 5122
rect 29260 5058 29316 5070
rect 29372 6018 29428 6030
rect 29372 5966 29374 6018
rect 29426 5966 29428 6018
rect 29148 5010 29204 5022
rect 29148 4958 29150 5010
rect 29202 4958 29204 5010
rect 29148 4676 29204 4958
rect 29148 4610 29204 4620
rect 29036 4386 29092 4396
rect 29148 4450 29204 4462
rect 29148 4398 29150 4450
rect 29202 4398 29204 4450
rect 28924 4172 29092 4228
rect 28812 3602 28868 3612
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 29036 3554 29092 4172
rect 29036 3502 29038 3554
rect 29090 3502 29092 3554
rect 29036 3490 29092 3502
rect 29148 3220 29204 4398
rect 29372 4228 29428 5966
rect 29484 5124 29540 7868
rect 29596 7028 29652 7038
rect 29596 6690 29652 6972
rect 29596 6638 29598 6690
rect 29650 6638 29652 6690
rect 29596 5684 29652 6638
rect 29708 6132 29764 8652
rect 29820 7700 29876 7710
rect 29820 7606 29876 7644
rect 29708 6066 29764 6076
rect 29932 5908 29988 9660
rect 30044 7924 30100 12236
rect 30492 12068 30548 12686
rect 30492 12002 30548 12012
rect 30604 12066 30660 12078
rect 30604 12014 30606 12066
rect 30658 12014 30660 12066
rect 30192 11788 30456 11798
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30192 11722 30456 11732
rect 30604 11284 30660 12014
rect 30156 11228 30660 11284
rect 30156 10722 30212 11228
rect 30156 10670 30158 10722
rect 30210 10670 30212 10722
rect 30156 10658 30212 10670
rect 30604 10724 30660 10734
rect 30192 10220 30456 10230
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30192 10154 30456 10164
rect 30492 10052 30548 10062
rect 30492 9154 30548 9996
rect 30492 9102 30494 9154
rect 30546 9102 30548 9154
rect 30492 9090 30548 9102
rect 30192 8652 30456 8662
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30192 8586 30456 8596
rect 30604 8484 30660 10668
rect 30492 8428 30660 8484
rect 30716 9042 30772 15092
rect 30940 14084 30996 14094
rect 30828 10610 30884 10622
rect 30828 10558 30830 10610
rect 30882 10558 30884 10610
rect 30828 10500 30884 10558
rect 30828 10434 30884 10444
rect 30940 9266 30996 14028
rect 31052 12738 31108 12750
rect 31052 12686 31054 12738
rect 31106 12686 31108 12738
rect 31052 11956 31108 12686
rect 31388 12292 31444 15092
rect 32172 13634 32228 13646
rect 32172 13582 32174 13634
rect 32226 13582 32228 13634
rect 31948 13522 32004 13534
rect 31948 13470 31950 13522
rect 32002 13470 32004 13522
rect 31948 13412 32004 13470
rect 31836 13356 32004 13412
rect 32172 13412 32228 13582
rect 31612 13300 31668 13310
rect 31276 12236 31444 12292
rect 31500 13244 31612 13300
rect 31052 11890 31108 11900
rect 31164 12180 31220 12190
rect 31164 11284 31220 12124
rect 31164 11218 31220 11228
rect 31164 10612 31220 10622
rect 31164 10518 31220 10556
rect 31276 9604 31332 12236
rect 31388 12068 31444 12078
rect 31388 11954 31444 12012
rect 31388 11902 31390 11954
rect 31442 11902 31444 11954
rect 31388 11890 31444 11902
rect 30940 9214 30942 9266
rect 30994 9214 30996 9266
rect 30940 9202 30996 9214
rect 31052 9548 31332 9604
rect 31388 10610 31444 10622
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 30716 8990 30718 9042
rect 30770 8990 30772 9042
rect 30268 8146 30324 8158
rect 30268 8094 30270 8146
rect 30322 8094 30324 8146
rect 30268 8036 30324 8094
rect 30268 7970 30324 7980
rect 30044 7700 30100 7868
rect 30156 7700 30212 7710
rect 30044 7698 30212 7700
rect 30044 7646 30158 7698
rect 30210 7646 30212 7698
rect 30044 7644 30212 7646
rect 30156 7634 30212 7644
rect 30492 7476 30548 8428
rect 30604 8260 30660 8270
rect 30604 7698 30660 8204
rect 30604 7646 30606 7698
rect 30658 7646 30660 7698
rect 30604 7634 30660 7646
rect 30716 7700 30772 8990
rect 30716 7634 30772 7644
rect 30940 8820 30996 8830
rect 30492 7420 30660 7476
rect 30604 7140 30660 7420
rect 30940 7362 30996 8764
rect 30940 7310 30942 7362
rect 30994 7310 30996 7362
rect 30940 7298 30996 7310
rect 30192 7084 30456 7094
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30192 7018 30456 7028
rect 29932 5814 29988 5852
rect 30604 5796 30660 7084
rect 31052 6244 31108 9548
rect 31388 9492 31444 10558
rect 31500 10052 31556 13244
rect 31612 13234 31668 13244
rect 31500 9986 31556 9996
rect 31612 12740 31668 12750
rect 30604 5730 30660 5740
rect 30716 6188 31108 6244
rect 31164 9436 31444 9492
rect 31164 8932 31220 9436
rect 31388 9156 31444 9166
rect 31388 9062 31444 9100
rect 31500 9044 31556 9054
rect 31500 8950 31556 8988
rect 31164 6690 31220 8876
rect 31388 8932 31444 8942
rect 31164 6638 31166 6690
rect 31218 6638 31220 6690
rect 29596 5628 29988 5684
rect 29820 5124 29876 5134
rect 29484 5068 29820 5124
rect 29820 5030 29876 5068
rect 29932 4338 29988 5628
rect 30192 5516 30456 5526
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30192 5450 30456 5460
rect 30492 5236 30548 5246
rect 30492 5142 30548 5180
rect 30604 5124 30660 5134
rect 30604 5030 30660 5068
rect 30716 4900 30772 6188
rect 31052 6020 31108 6030
rect 30940 5684 30996 5694
rect 30716 4834 30772 4844
rect 30828 5682 30996 5684
rect 30828 5630 30942 5682
rect 30994 5630 30996 5682
rect 30828 5628 30996 5630
rect 29932 4286 29934 4338
rect 29986 4286 29988 4338
rect 29932 4274 29988 4286
rect 29372 4162 29428 4172
rect 30192 3948 30456 3958
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30192 3882 30456 3892
rect 29148 3154 29204 3164
rect 29820 3444 29876 3454
rect 30828 3388 30884 5628
rect 30940 5618 30996 5628
rect 29148 2994 29204 3006
rect 29148 2942 29150 2994
rect 29202 2942 29204 2994
rect 29148 800 29204 2942
rect 29820 800 29876 3388
rect 30268 3332 30884 3388
rect 30940 4900 30996 4910
rect 30268 800 30324 3332
rect 30940 800 30996 4844
rect 31052 2436 31108 5964
rect 31164 4564 31220 6638
rect 31276 8820 31332 8830
rect 31276 6244 31332 8764
rect 31276 6178 31332 6188
rect 31388 5122 31444 8876
rect 31612 8036 31668 12684
rect 31724 12738 31780 12750
rect 31724 12686 31726 12738
rect 31778 12686 31780 12738
rect 31724 12180 31780 12686
rect 31836 12740 31892 13356
rect 32172 13346 32228 13356
rect 31948 12964 32004 12974
rect 31948 12962 32228 12964
rect 31948 12910 31950 12962
rect 32002 12910 32228 12962
rect 31948 12908 32228 12910
rect 31948 12898 32004 12908
rect 31836 12684 32004 12740
rect 31836 12292 31892 12302
rect 31836 12198 31892 12236
rect 31724 12114 31780 12124
rect 31724 11956 31780 11966
rect 31724 10722 31780 11900
rect 31836 11956 31892 11966
rect 31948 11956 32004 12684
rect 31836 11954 32004 11956
rect 31836 11902 31838 11954
rect 31890 11902 32004 11954
rect 31836 11900 32004 11902
rect 31836 11890 31892 11900
rect 31724 10670 31726 10722
rect 31778 10670 31780 10722
rect 31724 10658 31780 10670
rect 31948 10612 32004 11900
rect 32172 11844 32228 12908
rect 32284 12290 32340 12302
rect 32284 12238 32286 12290
rect 32338 12238 32340 12290
rect 32284 12180 32340 12238
rect 32396 12292 32452 15596
rect 32508 15586 32564 15596
rect 34748 15652 34804 15662
rect 34748 15202 34804 15596
rect 34748 15150 34750 15202
rect 34802 15150 34804 15202
rect 34748 15138 34804 15150
rect 35756 15426 35812 15438
rect 35756 15374 35758 15426
rect 35810 15374 35812 15426
rect 34860 14642 34916 14654
rect 34860 14590 34862 14642
rect 34914 14590 34916 14642
rect 33852 14418 33908 14430
rect 33852 14366 33854 14418
rect 33906 14366 33908 14418
rect 33404 13860 33460 13870
rect 33292 13748 33348 13758
rect 32508 13634 32564 13646
rect 33180 13636 33236 13646
rect 32508 13582 32510 13634
rect 32562 13582 32564 13634
rect 32508 13522 32564 13582
rect 32508 13470 32510 13522
rect 32562 13470 32564 13522
rect 32508 13458 32564 13470
rect 33068 13634 33236 13636
rect 33068 13582 33182 13634
rect 33234 13582 33236 13634
rect 33068 13580 33236 13582
rect 32508 12740 32564 12750
rect 32508 12738 32676 12740
rect 32508 12686 32510 12738
rect 32562 12686 32676 12738
rect 32508 12684 32676 12686
rect 32508 12674 32564 12684
rect 32508 12292 32564 12302
rect 32396 12290 32564 12292
rect 32396 12238 32510 12290
rect 32562 12238 32564 12290
rect 32396 12236 32564 12238
rect 32508 12226 32564 12236
rect 32284 12114 32340 12124
rect 32396 12068 32452 12078
rect 32396 11974 32452 12012
rect 32172 11788 32452 11844
rect 32172 11282 32228 11294
rect 32172 11230 32174 11282
rect 32226 11230 32228 11282
rect 31948 10610 32116 10612
rect 31948 10558 31950 10610
rect 32002 10558 32116 10610
rect 31948 10556 32116 10558
rect 31948 10546 32004 10556
rect 32060 9938 32116 10556
rect 32172 10052 32228 11230
rect 32284 10388 32340 10398
rect 32284 10294 32340 10332
rect 32172 9986 32228 9996
rect 32060 9886 32062 9938
rect 32114 9886 32116 9938
rect 31612 7970 31668 7980
rect 31948 8484 32004 8494
rect 31948 7586 32004 8428
rect 31948 7534 31950 7586
rect 32002 7534 32004 7586
rect 31948 7522 32004 7534
rect 32060 7252 32116 9886
rect 32396 9828 32452 11788
rect 32396 9762 32452 9772
rect 32620 9938 32676 12684
rect 32844 11396 32900 11406
rect 32844 10500 32900 11340
rect 32956 11060 33012 11070
rect 32956 10612 33012 11004
rect 33068 10836 33124 13580
rect 33180 13570 33236 13580
rect 33292 12964 33348 13692
rect 33180 12908 33348 12964
rect 33180 12180 33236 12908
rect 33292 12740 33348 12750
rect 33292 12646 33348 12684
rect 33404 12402 33460 13804
rect 33740 13634 33796 13646
rect 33740 13582 33742 13634
rect 33794 13582 33796 13634
rect 33404 12350 33406 12402
rect 33458 12350 33460 12402
rect 33404 12338 33460 12350
rect 33516 13074 33572 13086
rect 33516 13022 33518 13074
rect 33570 13022 33572 13074
rect 33516 12180 33572 13022
rect 33180 12178 33348 12180
rect 33180 12126 33182 12178
rect 33234 12126 33348 12178
rect 33180 12124 33348 12126
rect 33180 12114 33236 12124
rect 33292 10836 33348 12124
rect 33404 12124 33572 12180
rect 33404 11284 33460 12124
rect 33516 11956 33572 11966
rect 33516 11862 33572 11900
rect 33740 11788 33796 13582
rect 33852 12068 33908 14366
rect 34524 13858 34580 13870
rect 34524 13806 34526 13858
rect 34578 13806 34580 13858
rect 34524 13748 34580 13806
rect 34524 13682 34580 13692
rect 33852 12002 33908 12012
rect 34636 13634 34692 13646
rect 34636 13582 34638 13634
rect 34690 13582 34692 13634
rect 33628 11732 33796 11788
rect 34636 11844 34692 13582
rect 34636 11778 34692 11788
rect 34748 13522 34804 13534
rect 34748 13470 34750 13522
rect 34802 13470 34804 13522
rect 33516 11508 33572 11518
rect 33628 11508 33684 11732
rect 33516 11506 33684 11508
rect 33516 11454 33518 11506
rect 33570 11454 33684 11506
rect 33516 11452 33684 11454
rect 33516 11442 33572 11452
rect 33404 11228 33572 11284
rect 33404 10836 33460 10846
rect 33068 10780 33236 10836
rect 33292 10834 33460 10836
rect 33292 10782 33406 10834
rect 33458 10782 33460 10834
rect 33292 10780 33460 10782
rect 33068 10612 33124 10622
rect 32956 10610 33124 10612
rect 32956 10558 33070 10610
rect 33122 10558 33124 10610
rect 32956 10556 33124 10558
rect 33068 10546 33124 10556
rect 32844 10434 32900 10444
rect 32620 9886 32622 9938
rect 32674 9886 32676 9938
rect 32508 9042 32564 9054
rect 32508 8990 32510 9042
rect 32562 8990 32564 9042
rect 32508 8148 32564 8990
rect 32620 8932 32676 9886
rect 32620 8866 32676 8876
rect 33068 10388 33124 10398
rect 33068 9042 33124 10332
rect 33180 9156 33236 10780
rect 33404 10770 33460 10780
rect 33292 9828 33348 9838
rect 33516 9828 33572 11228
rect 33628 10836 33684 11452
rect 33628 10770 33684 10780
rect 33852 11060 33908 11070
rect 33852 10834 33908 11004
rect 33852 10782 33854 10834
rect 33906 10782 33908 10834
rect 33852 10770 33908 10782
rect 34412 10498 34468 10510
rect 34412 10446 34414 10498
rect 34466 10446 34468 10498
rect 34412 9940 34468 10446
rect 34748 10498 34804 13470
rect 34748 10446 34750 10498
rect 34802 10446 34804 10498
rect 34748 10434 34804 10446
rect 33348 9772 33460 9828
rect 33292 9762 33348 9772
rect 33180 9100 33348 9156
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 32508 8082 32564 8092
rect 33068 8036 33124 8990
rect 33068 7970 33124 7980
rect 33180 8930 33236 8942
rect 33180 8878 33182 8930
rect 33234 8878 33236 8930
rect 33180 7588 33236 8878
rect 32060 7186 32116 7196
rect 32508 7532 33236 7588
rect 31388 5070 31390 5122
rect 31442 5070 31444 5122
rect 31388 5058 31444 5070
rect 31948 6466 32004 6478
rect 31948 6414 31950 6466
rect 32002 6414 32004 6466
rect 31948 4900 32004 6414
rect 31948 4834 32004 4844
rect 31164 4498 31220 4508
rect 32172 4226 32228 4238
rect 32172 4174 32174 4226
rect 32226 4174 32228 4226
rect 31388 3666 31444 3678
rect 31388 3614 31390 3666
rect 31442 3614 31444 3666
rect 31388 3388 31444 3614
rect 31388 3332 31668 3388
rect 31052 2370 31108 2380
rect 31612 800 31668 3332
rect 32172 1316 32228 4174
rect 32396 3780 32452 3790
rect 32396 3666 32452 3724
rect 32508 3778 32564 7532
rect 33180 7364 33236 7374
rect 33068 7308 33180 7364
rect 32508 3726 32510 3778
rect 32562 3726 32564 3778
rect 32508 3714 32564 3726
rect 32956 5234 33012 5246
rect 32956 5182 32958 5234
rect 33010 5182 33012 5234
rect 32396 3614 32398 3666
rect 32450 3614 32452 3666
rect 32396 3602 32452 3614
rect 32284 3556 32340 3566
rect 32284 3442 32340 3500
rect 32284 3390 32286 3442
rect 32338 3390 32340 3442
rect 32284 3378 32340 3390
rect 32732 1540 32788 1550
rect 32172 1260 32340 1316
rect 32284 800 32340 1260
rect 32732 980 32788 1484
rect 32732 914 32788 924
rect 32956 800 33012 5182
rect 33068 4116 33124 7308
rect 33180 7270 33236 7308
rect 33292 7140 33348 9100
rect 33404 9154 33460 9772
rect 33516 9762 33572 9772
rect 34076 9884 34412 9940
rect 33740 9380 33796 9390
rect 33404 9102 33406 9154
rect 33458 9102 33460 9154
rect 33404 8932 33460 9102
rect 33516 9268 33572 9278
rect 33516 9042 33572 9212
rect 33516 8990 33518 9042
rect 33570 8990 33572 9042
rect 33516 8978 33572 8990
rect 33404 8866 33460 8876
rect 33628 8372 33684 8382
rect 33516 8148 33572 8158
rect 33516 7586 33572 8092
rect 33516 7534 33518 7586
rect 33570 7534 33572 7586
rect 33516 7522 33572 7534
rect 33628 7700 33684 8316
rect 33180 7084 33348 7140
rect 33180 6020 33236 7084
rect 33180 5926 33236 5964
rect 33292 6692 33348 6702
rect 33292 6018 33348 6636
rect 33628 6132 33684 7644
rect 33292 5966 33294 6018
rect 33346 5966 33348 6018
rect 33292 5954 33348 5966
rect 33404 6076 33684 6132
rect 33404 6018 33460 6076
rect 33404 5966 33406 6018
rect 33458 5966 33460 6018
rect 33404 5954 33460 5966
rect 33068 4050 33124 4060
rect 33180 4450 33236 4462
rect 33180 4398 33182 4450
rect 33234 4398 33236 4450
rect 33180 3444 33236 4398
rect 33628 4340 33684 4350
rect 33628 4226 33684 4284
rect 33628 4174 33630 4226
rect 33682 4174 33684 4226
rect 33628 3556 33684 4174
rect 33740 4004 33796 9324
rect 34076 8932 34132 9884
rect 34412 9846 34468 9884
rect 34748 9940 34804 9950
rect 34860 9940 34916 14590
rect 35756 14084 35812 15374
rect 37772 15148 37828 17164
rect 48300 17108 48356 17118
rect 42252 16884 42308 16894
rect 39852 15708 40116 15718
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 39852 15642 40116 15652
rect 37772 15092 38052 15148
rect 37324 14418 37380 14430
rect 37324 14366 37326 14418
rect 37378 14366 37380 14418
rect 35756 14018 35812 14028
rect 37100 14306 37156 14318
rect 37100 14254 37102 14306
rect 37154 14254 37156 14306
rect 35308 13860 35364 13870
rect 35308 13766 35364 13804
rect 37100 13748 37156 14254
rect 36316 13636 36372 13646
rect 35644 13634 36372 13636
rect 35644 13582 36318 13634
rect 36370 13582 36372 13634
rect 35644 13580 36372 13582
rect 35644 13074 35700 13580
rect 36316 13570 36372 13580
rect 35644 13022 35646 13074
rect 35698 13022 35700 13074
rect 35644 13010 35700 13022
rect 36316 12964 36372 12974
rect 35420 12628 35476 12638
rect 35308 12066 35364 12078
rect 35308 12014 35310 12066
rect 35362 12014 35364 12066
rect 35308 11396 35364 12014
rect 35308 11330 35364 11340
rect 35420 11060 35476 12572
rect 35308 11004 35420 11060
rect 34748 9938 34916 9940
rect 34748 9886 34750 9938
rect 34802 9886 34916 9938
rect 34748 9884 34916 9886
rect 34972 10052 35028 10062
rect 34748 9874 34804 9884
rect 34076 7474 34132 8876
rect 34188 9716 34244 9726
rect 34188 9266 34244 9660
rect 34188 9214 34190 9266
rect 34242 9214 34244 9266
rect 34188 8372 34244 9214
rect 34636 9268 34692 9278
rect 34636 9174 34692 9212
rect 34972 8930 35028 9996
rect 34972 8878 34974 8930
rect 35026 8878 35028 8930
rect 34972 8866 35028 8878
rect 35196 8932 35252 8942
rect 34860 8820 34916 8830
rect 34748 8764 34860 8820
rect 34188 8306 34244 8316
rect 34412 8484 34468 8494
rect 34412 8260 34468 8428
rect 34412 8166 34468 8204
rect 34076 7422 34078 7474
rect 34130 7422 34132 7474
rect 34076 7410 34132 7422
rect 34412 8036 34468 8046
rect 34412 7476 34468 7980
rect 34412 7382 34468 7420
rect 33852 6804 33908 6814
rect 33852 6130 33908 6748
rect 33852 6078 33854 6130
rect 33906 6078 33908 6130
rect 33852 6066 33908 6078
rect 34076 6802 34132 6814
rect 34076 6750 34078 6802
rect 34130 6750 34132 6802
rect 33964 4564 34020 4574
rect 33964 4338 34020 4508
rect 33964 4286 33966 4338
rect 34018 4286 34020 4338
rect 33964 4274 34020 4286
rect 33740 3938 33796 3948
rect 33628 3490 33684 3500
rect 34076 3388 34132 6750
rect 34524 5684 34580 5694
rect 33180 3378 33236 3388
rect 33628 3332 34132 3388
rect 34300 5682 34580 5684
rect 34300 5630 34526 5682
rect 34578 5630 34580 5682
rect 34300 5628 34580 5630
rect 33068 1540 33124 1550
rect 33068 1092 33124 1484
rect 33068 1026 33124 1036
rect 33628 800 33684 3332
rect 34300 800 34356 5628
rect 34524 5618 34580 5628
rect 34524 4452 34580 4462
rect 34524 4358 34580 4396
rect 34748 4340 34804 8764
rect 34860 8754 34916 8764
rect 34860 8146 34916 8158
rect 34860 8094 34862 8146
rect 34914 8094 34916 8146
rect 34860 7924 34916 8094
rect 34860 7858 34916 7868
rect 34972 8146 35028 8158
rect 34972 8094 34974 8146
rect 35026 8094 35028 8146
rect 34972 6692 35028 8094
rect 35084 8146 35140 8158
rect 35084 8094 35086 8146
rect 35138 8094 35140 8146
rect 35084 7700 35140 8094
rect 35084 7634 35140 7644
rect 35196 7476 35252 8876
rect 34972 6626 35028 6636
rect 35084 7420 35252 7476
rect 34860 4340 34916 4350
rect 34748 4338 34916 4340
rect 34748 4286 34862 4338
rect 34914 4286 34916 4338
rect 34748 4284 34916 4286
rect 34860 4274 34916 4284
rect 34412 3668 34468 3678
rect 34412 3574 34468 3612
rect 35084 3554 35140 7420
rect 35084 3502 35086 3554
rect 35138 3502 35140 3554
rect 35084 3490 35140 3502
rect 35196 5234 35252 5246
rect 35196 5182 35198 5234
rect 35250 5182 35252 5234
rect 35196 3388 35252 5182
rect 34972 3332 35252 3388
rect 35308 3332 35364 11004
rect 35420 10994 35476 11004
rect 35532 12180 35588 12190
rect 35532 10724 35588 12124
rect 35980 11844 36036 11854
rect 35644 11282 35700 11294
rect 35644 11230 35646 11282
rect 35698 11230 35700 11282
rect 35644 10948 35700 11230
rect 35644 10882 35700 10892
rect 35532 10668 35700 10724
rect 35532 10500 35588 10510
rect 35532 9826 35588 10444
rect 35532 9774 35534 9826
rect 35586 9774 35588 9826
rect 35532 9762 35588 9774
rect 35532 9156 35588 9166
rect 35532 8370 35588 9100
rect 35532 8318 35534 8370
rect 35586 8318 35588 8370
rect 35532 8306 35588 8318
rect 35644 7364 35700 10668
rect 35756 10052 35812 10062
rect 35756 7586 35812 9996
rect 35868 9940 35924 9950
rect 35868 9846 35924 9884
rect 35980 9154 36036 11788
rect 36316 11396 36372 12908
rect 36988 12964 37044 12974
rect 36988 12870 37044 12908
rect 37100 11732 37156 13692
rect 37212 14306 37268 14318
rect 37212 14254 37214 14306
rect 37266 14254 37268 14306
rect 37212 12516 37268 14254
rect 37212 12450 37268 12460
rect 37324 12068 37380 14366
rect 37996 14306 38052 15092
rect 37996 14254 37998 14306
rect 38050 14254 38052 14306
rect 37324 12002 37380 12012
rect 37548 13412 37604 13422
rect 37100 11666 37156 11676
rect 36316 11302 36372 11340
rect 36988 11394 37044 11406
rect 37212 11396 37268 11406
rect 36988 11342 36990 11394
rect 37042 11342 37044 11394
rect 36092 10724 36148 10734
rect 36092 10722 36260 10724
rect 36092 10670 36094 10722
rect 36146 10670 36260 10722
rect 36092 10668 36260 10670
rect 36092 10658 36148 10668
rect 35980 9102 35982 9154
rect 36034 9102 36036 9154
rect 35980 9090 36036 9102
rect 36092 9826 36148 9838
rect 36092 9774 36094 9826
rect 36146 9774 36148 9826
rect 36092 9268 36148 9774
rect 35868 8372 35924 8382
rect 35868 8258 35924 8316
rect 35868 8206 35870 8258
rect 35922 8206 35924 8258
rect 35868 7700 35924 8206
rect 35868 7634 35924 7644
rect 35756 7534 35758 7586
rect 35810 7534 35812 7586
rect 35756 7522 35812 7534
rect 35644 7308 35924 7364
rect 34972 800 35028 3332
rect 35308 2548 35364 3276
rect 35308 2482 35364 2492
rect 35644 3668 35700 3678
rect 35644 800 35700 3612
rect 35868 3444 35924 7308
rect 36092 6690 36148 9212
rect 36204 8596 36260 10668
rect 36652 10500 36708 10510
rect 36652 10406 36708 10444
rect 36988 10164 37044 11342
rect 36764 10108 37044 10164
rect 37100 11394 37268 11396
rect 37100 11342 37214 11394
rect 37266 11342 37268 11394
rect 37100 11340 37268 11342
rect 36428 10052 36484 10062
rect 36428 9958 36484 9996
rect 36316 9044 36372 9054
rect 36652 9044 36708 9054
rect 36372 8988 36484 9044
rect 36316 8978 36372 8988
rect 36316 8596 36372 8606
rect 36204 8540 36316 8596
rect 36316 8530 36372 8540
rect 36428 8372 36484 8988
rect 36316 8370 36484 8372
rect 36316 8318 36430 8370
rect 36482 8318 36484 8370
rect 36316 8316 36484 8318
rect 36204 7476 36260 7486
rect 36204 7382 36260 7420
rect 36092 6638 36094 6690
rect 36146 6638 36148 6690
rect 36092 6626 36148 6638
rect 36316 6692 36372 8316
rect 36428 8306 36484 8316
rect 36652 7586 36708 8988
rect 36652 7534 36654 7586
rect 36706 7534 36708 7586
rect 36316 6626 36372 6636
rect 36428 7474 36484 7486
rect 36428 7422 36430 7474
rect 36482 7422 36484 7474
rect 35980 6580 36036 6590
rect 35980 5236 36036 6524
rect 36428 6580 36484 7422
rect 36428 6514 36484 6524
rect 35980 5122 36036 5180
rect 35980 5070 35982 5122
rect 36034 5070 36036 5122
rect 35980 5058 36036 5070
rect 36652 4564 36708 7534
rect 36764 7476 36820 10108
rect 37100 10052 37156 11340
rect 37212 11330 37268 11340
rect 37548 11172 37604 13356
rect 37772 13076 37828 13086
rect 37772 12982 37828 13020
rect 37660 12740 37716 12750
rect 37660 12178 37716 12684
rect 37660 12126 37662 12178
rect 37714 12126 37716 12178
rect 37660 11844 37716 12126
rect 37660 11778 37716 11788
rect 37884 11732 37940 11742
rect 37884 11394 37940 11676
rect 37884 11342 37886 11394
rect 37938 11342 37940 11394
rect 37884 11330 37940 11342
rect 37548 11170 37716 11172
rect 37548 11118 37550 11170
rect 37602 11118 37716 11170
rect 37548 11116 37716 11118
rect 37548 11106 37604 11116
rect 37548 10948 37604 10958
rect 37212 10498 37268 10510
rect 37212 10446 37214 10498
rect 37266 10446 37268 10498
rect 37212 10108 37268 10446
rect 37548 10498 37604 10892
rect 37548 10446 37550 10498
rect 37602 10446 37604 10498
rect 37548 10434 37604 10446
rect 37212 10052 37492 10108
rect 37100 9986 37156 9996
rect 37436 9938 37492 10052
rect 37436 9886 37438 9938
rect 37490 9886 37492 9938
rect 36988 9828 37044 9838
rect 36764 7410 36820 7420
rect 36876 9772 36988 9828
rect 36876 5906 36932 9772
rect 36988 9734 37044 9772
rect 37212 9716 37268 9726
rect 37212 9154 37268 9660
rect 37212 9102 37214 9154
rect 37266 9102 37268 9154
rect 37100 9042 37156 9054
rect 37100 8990 37102 9042
rect 37154 8990 37156 9042
rect 37100 8820 37156 8990
rect 37212 8932 37268 9102
rect 37436 9044 37492 9886
rect 37436 8978 37492 8988
rect 37212 8866 37268 8876
rect 37548 8932 37604 8942
rect 37548 8838 37604 8876
rect 37100 8754 37156 8764
rect 37548 8708 37604 8718
rect 37436 8372 37492 8382
rect 37436 8278 37492 8316
rect 37212 8148 37268 8158
rect 37212 8054 37268 8092
rect 37324 8148 37380 8158
rect 37548 8148 37604 8652
rect 37324 8146 37604 8148
rect 37324 8094 37326 8146
rect 37378 8094 37604 8146
rect 37324 8092 37604 8094
rect 37324 8082 37380 8092
rect 36876 5854 36878 5906
rect 36930 5854 36932 5906
rect 36876 5842 36932 5854
rect 36988 6690 37044 6702
rect 36988 6638 36990 6690
rect 37042 6638 37044 6690
rect 36652 4498 36708 4508
rect 36204 4226 36260 4238
rect 36204 4174 36206 4226
rect 36258 4174 36260 4226
rect 35980 3444 36036 3454
rect 35868 3442 36036 3444
rect 35868 3390 35982 3442
rect 36034 3390 36036 3442
rect 35868 3388 36036 3390
rect 35980 3378 36036 3388
rect 36204 1316 36260 4174
rect 36988 3780 37044 6638
rect 37436 5682 37492 5694
rect 37436 5630 37438 5682
rect 37490 5630 37492 5682
rect 37212 5236 37268 5246
rect 37212 5122 37268 5180
rect 37212 5070 37214 5122
rect 37266 5070 37268 5122
rect 37212 5058 37268 5070
rect 36988 3714 37044 3724
rect 36316 3442 36372 3454
rect 36316 3390 36318 3442
rect 36370 3390 36372 3442
rect 36316 3332 36372 3390
rect 36316 3266 36372 3276
rect 36204 1260 36372 1316
rect 36316 800 36372 1260
rect 37436 980 37492 5630
rect 37660 5572 37716 11116
rect 37996 10612 38052 14254
rect 38108 14418 38164 14430
rect 38108 14366 38110 14418
rect 38162 14366 38164 14418
rect 38108 14308 38164 14366
rect 38556 14308 38612 14318
rect 38108 14306 38612 14308
rect 38108 14254 38558 14306
rect 38610 14254 38612 14306
rect 38108 14252 38612 14254
rect 38108 13860 38164 13870
rect 38108 11506 38164 13804
rect 38108 11454 38110 11506
rect 38162 11454 38164 11506
rect 38108 11442 38164 11454
rect 38220 11284 38276 11294
rect 38220 11190 38276 11228
rect 37996 10556 38164 10612
rect 37996 10388 38052 10398
rect 37996 9940 38052 10332
rect 37884 9938 38052 9940
rect 37884 9886 37998 9938
rect 38050 9886 38052 9938
rect 37884 9884 38052 9886
rect 37772 8258 37828 8270
rect 37772 8206 37774 8258
rect 37826 8206 37828 8258
rect 37772 7364 37828 8206
rect 37884 8148 37940 9884
rect 37996 9874 38052 9884
rect 38108 9156 38164 10556
rect 38108 9090 38164 9100
rect 37996 8930 38052 8942
rect 37996 8878 37998 8930
rect 38050 8878 38052 8930
rect 37996 8820 38052 8878
rect 37996 8754 38052 8764
rect 37884 7476 37940 8092
rect 37884 7410 37940 7420
rect 38108 8596 38164 8606
rect 37772 7298 37828 7308
rect 37996 6692 38052 6702
rect 37996 6598 38052 6636
rect 37548 4340 37604 4350
rect 37660 4340 37716 5516
rect 37772 6580 37828 6590
rect 37772 5346 37828 6524
rect 38108 6466 38164 8540
rect 38332 7476 38388 14252
rect 38556 14242 38612 14252
rect 39852 14140 40116 14150
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 39852 14074 40116 14084
rect 39900 13860 39956 13870
rect 39900 13766 39956 13804
rect 38892 13634 38948 13646
rect 38892 13582 38894 13634
rect 38946 13582 38948 13634
rect 38892 13076 38948 13582
rect 40572 13636 40628 13646
rect 40236 13188 40292 13198
rect 39900 13076 39956 13086
rect 38892 13010 38948 13020
rect 39340 13074 39956 13076
rect 39340 13022 39902 13074
rect 39954 13022 39956 13074
rect 39340 13020 39956 13022
rect 38556 12516 38612 12526
rect 38612 12460 38724 12516
rect 38556 12450 38612 12460
rect 38668 10722 38724 12460
rect 38892 12068 38948 12078
rect 38668 10670 38670 10722
rect 38722 10670 38724 10722
rect 38668 10658 38724 10670
rect 38780 11170 38836 11182
rect 38780 11118 38782 11170
rect 38834 11118 38836 11170
rect 38780 10052 38836 11118
rect 38556 9996 38836 10052
rect 38556 9044 38612 9996
rect 38892 9938 38948 12012
rect 39116 11956 39172 11966
rect 38892 9886 38894 9938
rect 38946 9886 38948 9938
rect 38892 9874 38948 9886
rect 39004 10836 39060 10846
rect 38668 9604 38724 9614
rect 38668 9602 38836 9604
rect 38668 9550 38670 9602
rect 38722 9550 38836 9602
rect 38668 9548 38836 9550
rect 38668 9538 38724 9548
rect 38556 8930 38612 8988
rect 38556 8878 38558 8930
rect 38610 8878 38612 8930
rect 38556 8820 38612 8878
rect 38556 8754 38612 8764
rect 38668 8036 38724 8046
rect 38444 7812 38500 7822
rect 38444 7698 38500 7756
rect 38444 7646 38446 7698
rect 38498 7646 38500 7698
rect 38444 7634 38500 7646
rect 38556 7700 38612 7710
rect 38556 7606 38612 7644
rect 38668 7698 38724 7980
rect 38780 7812 38836 9548
rect 38892 8932 38948 8942
rect 38892 8146 38948 8876
rect 39004 8708 39060 10780
rect 39116 8930 39172 11900
rect 39340 10722 39396 13020
rect 39900 13010 39956 13020
rect 40236 12852 40292 13132
rect 39852 12572 40116 12582
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 39852 12506 40116 12516
rect 40236 12402 40292 12796
rect 40460 12738 40516 12750
rect 40460 12686 40462 12738
rect 40514 12686 40516 12738
rect 40460 12628 40516 12686
rect 40460 12562 40516 12572
rect 40572 12404 40628 13580
rect 41132 13634 41188 13646
rect 41132 13582 41134 13634
rect 41186 13582 41188 13634
rect 41132 13076 41188 13582
rect 41468 13524 41524 13534
rect 41132 13020 41412 13076
rect 41244 12850 41300 12862
rect 41244 12798 41246 12850
rect 41298 12798 41300 12850
rect 40236 12350 40238 12402
rect 40290 12350 40292 12402
rect 40236 12338 40292 12350
rect 40460 12348 40628 12404
rect 40796 12738 40852 12750
rect 40796 12686 40798 12738
rect 40850 12686 40852 12738
rect 40796 12404 40852 12686
rect 39900 12180 39956 12190
rect 40348 12180 40404 12190
rect 39900 12178 40292 12180
rect 39900 12126 39902 12178
rect 39954 12126 40292 12178
rect 39900 12124 40292 12126
rect 39900 12114 39956 12124
rect 39340 10670 39342 10722
rect 39394 10670 39396 10722
rect 39340 10164 39396 10670
rect 39564 11954 39620 11966
rect 39564 11902 39566 11954
rect 39618 11902 39620 11954
rect 39452 10388 39508 10398
rect 39452 10294 39508 10332
rect 39564 10164 39620 11902
rect 39900 11956 39956 11966
rect 39900 11862 39956 11900
rect 39676 11172 39732 11182
rect 39676 10724 39732 11116
rect 39852 11004 40116 11014
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 39852 10938 40116 10948
rect 40236 10836 40292 12124
rect 40348 12086 40404 12124
rect 40012 10780 40292 10836
rect 39788 10724 39844 10734
rect 39676 10722 39844 10724
rect 39676 10670 39790 10722
rect 39842 10670 39844 10722
rect 39676 10668 39844 10670
rect 39788 10658 39844 10668
rect 39564 10108 39732 10164
rect 39340 10098 39396 10108
rect 39564 9940 39620 9950
rect 39116 8878 39118 8930
rect 39170 8878 39172 8930
rect 39116 8866 39172 8878
rect 39228 9828 39284 9838
rect 39228 8932 39284 9772
rect 39228 8866 39284 8876
rect 39452 9604 39508 9614
rect 39004 8652 39172 8708
rect 38892 8094 38894 8146
rect 38946 8094 38948 8146
rect 38892 8082 38948 8094
rect 38780 7756 39060 7812
rect 38668 7646 38670 7698
rect 38722 7646 38724 7698
rect 38668 7634 38724 7646
rect 38892 7588 38948 7598
rect 38780 7532 38892 7588
rect 38332 7420 38500 7476
rect 38220 7364 38276 7374
rect 38276 7308 38388 7364
rect 38220 7270 38276 7308
rect 38220 6916 38276 6926
rect 38220 6578 38276 6860
rect 38220 6526 38222 6578
rect 38274 6526 38276 6578
rect 38220 6514 38276 6526
rect 38108 6414 38110 6466
rect 38162 6414 38164 6466
rect 38108 6402 38164 6414
rect 37772 5294 37774 5346
rect 37826 5294 37828 5346
rect 37772 5282 37828 5294
rect 37884 5348 37940 5358
rect 37884 5234 37940 5292
rect 37884 5182 37886 5234
rect 37938 5182 37940 5234
rect 37884 5170 37940 5182
rect 38332 5124 38388 7308
rect 38444 5908 38500 7420
rect 38780 7140 38836 7532
rect 38892 7522 38948 7532
rect 39004 7474 39060 7756
rect 39004 7422 39006 7474
rect 39058 7422 39060 7474
rect 38444 5842 38500 5852
rect 38556 7084 38836 7140
rect 38892 7140 38948 7150
rect 38444 5124 38500 5134
rect 38332 5122 38500 5124
rect 38332 5070 38446 5122
rect 38498 5070 38500 5122
rect 38332 5068 38500 5070
rect 38444 5058 38500 5068
rect 37604 4284 37716 4340
rect 37548 4274 37604 4284
rect 38332 4226 38388 4238
rect 38332 4174 38334 4226
rect 38386 4174 38388 4226
rect 36988 924 37492 980
rect 37660 3442 37716 3454
rect 37660 3390 37662 3442
rect 37714 3390 37716 3442
rect 36988 800 37044 924
rect 37660 800 37716 3390
rect 38332 800 38388 4174
rect 38556 2884 38612 7084
rect 38892 7028 38948 7084
rect 38668 6972 38948 7028
rect 38668 4900 38724 6972
rect 38892 6578 38948 6590
rect 38892 6526 38894 6578
rect 38946 6526 38948 6578
rect 38780 4900 38836 4910
rect 38668 4898 38836 4900
rect 38668 4846 38782 4898
rect 38834 4846 38836 4898
rect 38668 4844 38836 4846
rect 38780 4834 38836 4844
rect 38556 2818 38612 2828
rect 38780 3554 38836 3566
rect 38780 3502 38782 3554
rect 38834 3502 38836 3554
rect 38780 1540 38836 3502
rect 38892 2882 38948 6526
rect 39004 3892 39060 7422
rect 39116 6690 39172 8652
rect 39452 8372 39508 9548
rect 39116 6638 39118 6690
rect 39170 6638 39172 6690
rect 39116 6626 39172 6638
rect 39228 8148 39284 8158
rect 39004 3826 39060 3836
rect 39228 3332 39284 8092
rect 39340 8036 39396 8046
rect 39340 6468 39396 7980
rect 39452 7474 39508 8316
rect 39452 7422 39454 7474
rect 39506 7422 39508 7474
rect 39452 7140 39508 7422
rect 39452 7074 39508 7084
rect 39564 6804 39620 9884
rect 39676 9828 39732 10108
rect 39676 9762 39732 9772
rect 39900 9714 39956 9726
rect 39900 9662 39902 9714
rect 39954 9662 39956 9714
rect 39900 9604 39956 9662
rect 39676 9548 39956 9604
rect 40012 9604 40068 10780
rect 40124 10610 40180 10622
rect 40124 10558 40126 10610
rect 40178 10558 40180 10610
rect 40124 9716 40180 10558
rect 40348 10612 40404 10622
rect 40348 10518 40404 10556
rect 40236 10498 40292 10510
rect 40236 10446 40238 10498
rect 40290 10446 40292 10498
rect 40236 10164 40292 10446
rect 40236 10098 40292 10108
rect 40124 9650 40180 9660
rect 39676 8036 39732 9548
rect 40012 9538 40068 9548
rect 39852 9436 40116 9446
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 39852 9370 40116 9380
rect 40236 9154 40292 9166
rect 40236 9102 40238 9154
rect 40290 9102 40292 9154
rect 39900 8372 39956 8382
rect 39900 8258 39956 8316
rect 39900 8206 39902 8258
rect 39954 8206 39956 8258
rect 39900 8194 39956 8206
rect 39676 7970 39732 7980
rect 39852 7868 40116 7878
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 39852 7802 40116 7812
rect 39900 7476 39956 7486
rect 39900 7382 39956 7420
rect 40236 6916 40292 9102
rect 40348 9156 40404 9166
rect 40348 8146 40404 9100
rect 40348 8094 40350 8146
rect 40402 8094 40404 8146
rect 40348 7700 40404 8094
rect 40348 7634 40404 7644
rect 40348 7364 40404 7374
rect 40348 7270 40404 7308
rect 40236 6860 40404 6916
rect 39340 6402 39396 6412
rect 39452 6748 39620 6804
rect 40012 6804 40068 6814
rect 39452 6020 39508 6748
rect 40012 6710 40068 6748
rect 39788 6692 39844 6702
rect 39788 6598 39844 6636
rect 40236 6690 40292 6702
rect 40236 6638 40238 6690
rect 40290 6638 40292 6690
rect 39452 5954 39508 5964
rect 39564 6578 39620 6590
rect 39564 6526 39566 6578
rect 39618 6526 39620 6578
rect 39340 5908 39396 5918
rect 39340 5814 39396 5852
rect 39228 3266 39284 3276
rect 39452 5234 39508 5246
rect 39452 5182 39454 5234
rect 39506 5182 39508 5234
rect 38892 2830 38894 2882
rect 38946 2830 38948 2882
rect 38892 2818 38948 2830
rect 38780 1474 38836 1484
rect 39452 980 39508 5182
rect 39564 4452 39620 6526
rect 40236 6468 40292 6638
rect 40348 6690 40404 6860
rect 40348 6638 40350 6690
rect 40402 6638 40404 6690
rect 40348 6626 40404 6638
rect 40460 6690 40516 12348
rect 40796 12338 40852 12348
rect 41244 12292 41300 12798
rect 41356 12852 41412 13020
rect 41356 12758 41412 12796
rect 41244 12236 41412 12292
rect 40572 12180 40628 12190
rect 40572 6916 40628 12124
rect 40908 12068 40964 12078
rect 40684 12066 40964 12068
rect 40684 12014 40910 12066
rect 40962 12014 40964 12066
rect 40684 12012 40964 12014
rect 40684 8708 40740 12012
rect 40908 12002 40964 12012
rect 41244 12068 41300 12078
rect 41244 11974 41300 12012
rect 40908 11844 40964 11854
rect 40908 10610 40964 11788
rect 41020 11284 41076 11294
rect 41020 11282 41188 11284
rect 41020 11230 41022 11282
rect 41074 11230 41188 11282
rect 41020 11228 41188 11230
rect 41020 11218 41076 11228
rect 40908 10558 40910 10610
rect 40962 10558 40964 10610
rect 40796 9940 40852 9950
rect 40908 9940 40964 10558
rect 41020 10948 41076 10958
rect 41020 10052 41076 10892
rect 41020 9986 41076 9996
rect 40796 9938 40964 9940
rect 40796 9886 40798 9938
rect 40850 9886 40964 9938
rect 40796 9884 40964 9886
rect 40796 9874 40852 9884
rect 41020 9828 41076 9838
rect 40908 9604 40964 9614
rect 40908 9042 40964 9548
rect 40908 8990 40910 9042
rect 40962 8990 40964 9042
rect 40908 8978 40964 8990
rect 41020 9042 41076 9772
rect 41020 8990 41022 9042
rect 41074 8990 41076 9042
rect 41020 8978 41076 8990
rect 41132 8820 41188 11228
rect 41356 10948 41412 12236
rect 41356 10882 41412 10892
rect 41468 10724 41524 13468
rect 41580 12740 41636 12750
rect 41580 12646 41636 12684
rect 42028 12738 42084 12750
rect 42028 12686 42030 12738
rect 42082 12686 42084 12738
rect 42028 12404 42084 12686
rect 42028 12338 42084 12348
rect 41580 12180 41636 12190
rect 41636 12124 41860 12180
rect 41580 12114 41636 12124
rect 41804 12066 41860 12124
rect 41804 12014 41806 12066
rect 41858 12014 41860 12066
rect 41804 12002 41860 12014
rect 41356 10668 41524 10724
rect 41692 11394 41748 11406
rect 41692 11342 41694 11394
rect 41746 11342 41748 11394
rect 41132 8754 41188 8764
rect 41244 10276 41300 10286
rect 40684 8652 41076 8708
rect 41020 8372 41076 8652
rect 40908 8260 40964 8270
rect 40796 8204 40908 8260
rect 41020 8260 41076 8316
rect 41020 8204 41188 8260
rect 40684 6916 40740 6926
rect 40572 6914 40740 6916
rect 40572 6862 40686 6914
rect 40738 6862 40740 6914
rect 40572 6860 40740 6862
rect 40684 6850 40740 6860
rect 40460 6638 40462 6690
rect 40514 6638 40516 6690
rect 40460 6626 40516 6638
rect 39564 4386 39620 4396
rect 39676 6412 40292 6468
rect 39676 4228 39732 6412
rect 39852 6300 40116 6310
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 39852 6234 40116 6244
rect 40236 6132 40292 6142
rect 40796 6132 40852 8204
rect 40908 8194 40964 8204
rect 41020 8034 41076 8046
rect 41020 7982 41022 8034
rect 41074 7982 41076 8034
rect 40908 7476 40964 7486
rect 40908 6802 40964 7420
rect 40908 6750 40910 6802
rect 40962 6750 40964 6802
rect 40908 6738 40964 6750
rect 41020 6804 41076 7982
rect 41132 7698 41188 8204
rect 41132 7646 41134 7698
rect 41186 7646 41188 7698
rect 41132 7588 41188 7646
rect 41132 7522 41188 7532
rect 40908 6132 40964 6142
rect 40236 6038 40292 6076
rect 40348 6130 40964 6132
rect 40348 6078 40910 6130
rect 40962 6078 40964 6130
rect 40348 6076 40964 6078
rect 39788 6020 39844 6030
rect 40012 6020 40068 6030
rect 39844 6018 40068 6020
rect 39844 5966 40014 6018
rect 40066 5966 40068 6018
rect 39844 5964 40068 5966
rect 39788 5954 39844 5964
rect 40012 5954 40068 5964
rect 40348 6018 40404 6076
rect 40908 6066 40964 6076
rect 40348 5966 40350 6018
rect 40402 5966 40404 6018
rect 40348 5954 40404 5966
rect 41020 5908 41076 6748
rect 41132 7364 41188 7374
rect 41132 6244 41188 7308
rect 41132 6178 41188 6188
rect 41132 5908 41188 5918
rect 41020 5906 41188 5908
rect 41020 5854 41134 5906
rect 41186 5854 41188 5906
rect 41020 5852 41188 5854
rect 41132 5842 41188 5852
rect 39852 4732 40116 4742
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 39852 4666 40116 4676
rect 40908 4452 40964 4462
rect 40348 4340 40404 4350
rect 40348 4246 40404 4284
rect 39564 4172 39732 4228
rect 39564 2436 39620 4172
rect 39900 4116 39956 4126
rect 39564 2370 39620 2380
rect 39676 4060 39900 4116
rect 39004 924 39508 980
rect 39004 800 39060 924
rect 39676 800 39732 4060
rect 39900 4050 39956 4060
rect 40684 3666 40740 3678
rect 40684 3614 40686 3666
rect 40738 3614 40740 3666
rect 40684 3388 40740 3614
rect 40012 3332 40068 3342
rect 40348 3332 40740 3388
rect 40012 3330 40292 3332
rect 40012 3278 40014 3330
rect 40066 3278 40292 3330
rect 40012 3276 40292 3278
rect 40012 3266 40068 3276
rect 39852 3164 40116 3174
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 39852 3098 40116 3108
rect 40236 2882 40292 3276
rect 40236 2830 40238 2882
rect 40290 2830 40292 2882
rect 40236 2818 40292 2830
rect 40348 800 40404 3332
rect 40908 980 40964 4396
rect 41132 4116 41188 4126
rect 41132 4022 41188 4060
rect 40908 914 40964 924
rect 41020 3444 41076 3454
rect 41020 800 41076 3388
rect 41244 3388 41300 10220
rect 41356 9380 41412 10668
rect 41468 10500 41524 10510
rect 41692 10500 41748 11342
rect 41524 10444 41748 10500
rect 41916 11284 41972 11294
rect 41468 9938 41524 10444
rect 41468 9886 41470 9938
rect 41522 9886 41524 9938
rect 41468 9874 41524 9886
rect 41692 9716 41748 9726
rect 41356 9324 41524 9380
rect 41356 9154 41412 9166
rect 41356 9102 41358 9154
rect 41410 9102 41412 9154
rect 41356 8372 41412 9102
rect 41356 8306 41412 8316
rect 41356 7924 41412 7934
rect 41468 7924 41524 9324
rect 41692 9266 41748 9660
rect 41692 9214 41694 9266
rect 41746 9214 41748 9266
rect 41692 9202 41748 9214
rect 41580 9042 41636 9054
rect 41580 8990 41582 9042
rect 41634 8990 41636 9042
rect 41580 8708 41636 8990
rect 41804 9044 41860 9054
rect 41804 8950 41860 8988
rect 41580 8642 41636 8652
rect 41468 7868 41748 7924
rect 41356 7140 41412 7868
rect 41580 7700 41636 7710
rect 41580 7606 41636 7644
rect 41692 7476 41748 7868
rect 41356 7084 41524 7140
rect 41468 7028 41524 7084
rect 41468 6972 41636 7028
rect 41356 6914 41412 6926
rect 41356 6862 41358 6914
rect 41410 6862 41412 6914
rect 41356 5236 41412 6862
rect 41580 6748 41636 6972
rect 41356 5122 41412 5180
rect 41356 5070 41358 5122
rect 41410 5070 41412 5122
rect 41356 5058 41412 5070
rect 41468 6692 41636 6748
rect 41468 4116 41524 6692
rect 41580 6580 41636 6590
rect 41580 6486 41636 6524
rect 41692 6130 41748 7420
rect 41916 7362 41972 11228
rect 42140 11172 42196 11182
rect 42140 11078 42196 11116
rect 42028 10164 42084 10174
rect 42028 9714 42084 10108
rect 42028 9662 42030 9714
rect 42082 9662 42084 9714
rect 42028 9650 42084 9662
rect 42028 8820 42084 8830
rect 42028 8370 42084 8764
rect 42028 8318 42030 8370
rect 42082 8318 42084 8370
rect 42028 8306 42084 8318
rect 42252 8148 42308 16828
rect 46060 13972 46116 13982
rect 43372 13524 43428 13534
rect 42476 12738 42532 12750
rect 42476 12686 42478 12738
rect 42530 12686 42532 12738
rect 42364 12628 42420 12638
rect 42364 11394 42420 12572
rect 42476 12068 42532 12686
rect 42812 12738 42868 12750
rect 42812 12686 42814 12738
rect 42866 12686 42868 12738
rect 42812 12628 42868 12686
rect 42812 12562 42868 12572
rect 42476 12002 42532 12012
rect 43260 12292 43316 12302
rect 43148 11844 43204 11854
rect 42364 11342 42366 11394
rect 42418 11342 42420 11394
rect 42364 11330 42420 11342
rect 43036 11788 43148 11844
rect 42812 11282 42868 11294
rect 42812 11230 42814 11282
rect 42866 11230 42868 11282
rect 42812 11172 42868 11230
rect 42812 11106 42868 11116
rect 42476 10612 42532 10622
rect 41916 7310 41918 7362
rect 41970 7310 41972 7362
rect 41916 7298 41972 7310
rect 42028 8092 42308 8148
rect 42364 9828 42420 9838
rect 42028 6914 42084 8092
rect 42364 8036 42420 9772
rect 42028 6862 42030 6914
rect 42082 6862 42084 6914
rect 42028 6850 42084 6862
rect 42140 7980 42420 8036
rect 41804 6692 41860 6702
rect 42140 6692 42196 7980
rect 41804 6598 41860 6636
rect 41916 6636 42140 6692
rect 41692 6078 41694 6130
rect 41746 6078 41748 6130
rect 41692 6066 41748 6078
rect 41468 4050 41524 4060
rect 41804 5906 41860 5918
rect 41804 5854 41806 5906
rect 41858 5854 41860 5906
rect 41804 4228 41860 5854
rect 41916 4340 41972 6636
rect 42140 6626 42196 6636
rect 42252 7812 42308 7822
rect 42252 6690 42308 7756
rect 42476 7700 42532 10556
rect 42700 9044 42756 9054
rect 42476 7634 42532 7644
rect 42588 8930 42644 8942
rect 42588 8878 42590 8930
rect 42642 8878 42644 8930
rect 42588 7476 42644 8878
rect 42700 7924 42756 8988
rect 42700 7858 42756 7868
rect 42812 7588 42868 7598
rect 42476 7420 42644 7476
rect 42700 7532 42812 7588
rect 42252 6638 42254 6690
rect 42306 6638 42308 6690
rect 42252 6626 42308 6638
rect 42364 7364 42420 7374
rect 42028 6468 42084 6478
rect 42364 6468 42420 7308
rect 42476 7140 42532 7420
rect 42476 7074 42532 7084
rect 42588 7028 42644 7038
rect 42028 6374 42084 6412
rect 42140 6412 42420 6468
rect 42476 6578 42532 6590
rect 42476 6526 42478 6578
rect 42530 6526 42532 6578
rect 42140 6132 42196 6412
rect 42476 6356 42532 6526
rect 42364 6300 42532 6356
rect 42028 6076 42196 6132
rect 42252 6132 42308 6142
rect 42028 5236 42084 6076
rect 42252 6018 42308 6076
rect 42252 5966 42254 6018
rect 42306 5966 42308 6018
rect 42252 5954 42308 5966
rect 42140 5906 42196 5918
rect 42140 5854 42142 5906
rect 42194 5854 42196 5906
rect 42140 5684 42196 5854
rect 42140 5618 42196 5628
rect 42252 5796 42308 5806
rect 42028 5180 42196 5236
rect 41916 4274 41972 4284
rect 42028 5012 42084 5022
rect 41244 3332 41748 3388
rect 41692 800 41748 3332
rect 41804 3108 41860 4172
rect 41916 3108 41972 3118
rect 41804 3052 41916 3108
rect 41916 3042 41972 3052
rect 42028 1204 42084 4956
rect 42140 3220 42196 5180
rect 42140 3154 42196 3164
rect 42252 5122 42308 5740
rect 42252 5070 42254 5122
rect 42306 5070 42308 5122
rect 42252 1316 42308 5070
rect 42364 2884 42420 6300
rect 42476 6132 42532 6142
rect 42476 5684 42532 6076
rect 42588 5906 42644 6972
rect 42588 5854 42590 5906
rect 42642 5854 42644 5906
rect 42588 5842 42644 5854
rect 42476 5628 42644 5684
rect 42476 4900 42532 4910
rect 42476 4806 42532 4844
rect 42476 4676 42532 4686
rect 42476 3444 42532 4620
rect 42588 3554 42644 5628
rect 42700 5234 42756 7532
rect 42812 7522 42868 7532
rect 42924 7586 42980 7598
rect 42924 7534 42926 7586
rect 42978 7534 42980 7586
rect 42812 6692 42868 6702
rect 42812 6598 42868 6636
rect 42812 6468 42868 6478
rect 42812 5906 42868 6412
rect 42924 6130 42980 7534
rect 43036 7588 43092 11788
rect 43148 11778 43204 11788
rect 43260 11506 43316 12236
rect 43260 11454 43262 11506
rect 43314 11454 43316 11506
rect 43260 11442 43316 11454
rect 43148 11394 43204 11406
rect 43148 11342 43150 11394
rect 43202 11342 43204 11394
rect 43148 9716 43204 11342
rect 43372 10052 43428 13468
rect 44044 13076 44100 13086
rect 43932 12740 43988 12750
rect 43932 11508 43988 12684
rect 44044 12290 44100 13020
rect 45164 12738 45220 12750
rect 45612 12740 45668 12750
rect 45164 12686 45166 12738
rect 45218 12686 45220 12738
rect 44044 12238 44046 12290
rect 44098 12238 44100 12290
rect 44044 12226 44100 12238
rect 44268 12404 44324 12414
rect 44268 11788 44324 12348
rect 44716 12180 44772 12190
rect 45164 12180 45220 12686
rect 44716 12178 45220 12180
rect 44716 12126 44718 12178
rect 44770 12126 45220 12178
rect 44716 12124 45220 12126
rect 45500 12738 45668 12740
rect 45500 12686 45614 12738
rect 45666 12686 45668 12738
rect 45500 12684 45668 12686
rect 44268 11732 44548 11788
rect 43932 11452 44100 11508
rect 43148 9650 43204 9660
rect 43260 9996 43428 10052
rect 43484 11394 43540 11406
rect 43484 11342 43486 11394
rect 43538 11342 43540 11394
rect 43260 7700 43316 9996
rect 43484 9940 43540 11342
rect 43708 11282 43764 11294
rect 43708 11230 43710 11282
rect 43762 11230 43764 11282
rect 43708 11172 43764 11230
rect 43708 11106 43764 11116
rect 43932 11282 43988 11294
rect 43932 11230 43934 11282
rect 43986 11230 43988 11282
rect 43708 10500 43764 10510
rect 43708 10406 43764 10444
rect 43484 9884 43876 9940
rect 43708 9716 43764 9726
rect 43372 9604 43428 9614
rect 43372 8146 43428 9548
rect 43596 9156 43652 9166
rect 43372 8094 43374 8146
rect 43426 8094 43428 8146
rect 43372 8082 43428 8094
rect 43484 8820 43540 8830
rect 43260 7644 43428 7700
rect 43036 7532 43316 7588
rect 43148 7364 43204 7374
rect 42924 6078 42926 6130
rect 42978 6078 42980 6130
rect 42924 6066 42980 6078
rect 43036 7140 43092 7150
rect 43036 6578 43092 7084
rect 43148 6914 43204 7308
rect 43148 6862 43150 6914
rect 43202 6862 43204 6914
rect 43148 6850 43204 6862
rect 43036 6526 43038 6578
rect 43090 6526 43092 6578
rect 42812 5854 42814 5906
rect 42866 5854 42868 5906
rect 42812 5842 42868 5854
rect 42700 5182 42702 5234
rect 42754 5182 42756 5234
rect 42700 5170 42756 5182
rect 42924 5460 42980 5470
rect 42924 5122 42980 5404
rect 42924 5070 42926 5122
rect 42978 5070 42980 5122
rect 42924 5058 42980 5070
rect 42700 4900 42756 4910
rect 42700 4898 42980 4900
rect 42700 4846 42702 4898
rect 42754 4846 42980 4898
rect 42700 4844 42980 4846
rect 42700 4834 42756 4844
rect 42812 4676 42868 4686
rect 42588 3502 42590 3554
rect 42642 3502 42644 3554
rect 42588 3490 42644 3502
rect 42700 4228 42756 4238
rect 42476 3378 42532 3388
rect 42700 2996 42756 4172
rect 42700 2930 42756 2940
rect 42364 2818 42420 2828
rect 42812 2658 42868 4620
rect 42924 2770 42980 4844
rect 43036 4338 43092 6526
rect 43036 4286 43038 4338
rect 43090 4286 43092 4338
rect 43036 4274 43092 4286
rect 43148 6018 43204 6030
rect 43148 5966 43150 6018
rect 43202 5966 43204 6018
rect 43148 5684 43204 5966
rect 42924 2718 42926 2770
rect 42978 2718 42980 2770
rect 42924 2706 42980 2718
rect 43036 4116 43092 4126
rect 42812 2606 42814 2658
rect 42866 2606 42868 2658
rect 42812 2594 42868 2606
rect 42252 1250 42308 1260
rect 42028 1138 42084 1148
rect 42364 978 42420 990
rect 42364 926 42366 978
rect 42418 926 42420 978
rect 42364 800 42420 926
rect 43036 800 43092 4060
rect 43148 3780 43204 5628
rect 43148 3714 43204 3724
rect 43148 3444 43204 3454
rect 43148 980 43204 3388
rect 43260 2546 43316 7532
rect 43372 6468 43428 7644
rect 43372 6402 43428 6412
rect 43372 5906 43428 5918
rect 43372 5854 43374 5906
rect 43426 5854 43428 5906
rect 43372 3668 43428 5854
rect 43484 5236 43540 8764
rect 43596 7364 43652 9100
rect 43708 8482 43764 9660
rect 43820 8596 43876 9884
rect 43820 8530 43876 8540
rect 43708 8430 43710 8482
rect 43762 8430 43764 8482
rect 43708 8418 43764 8430
rect 43820 8036 43876 8046
rect 43596 7298 43652 7308
rect 43708 8034 43876 8036
rect 43708 7982 43822 8034
rect 43874 7982 43876 8034
rect 43708 7980 43876 7982
rect 43708 7140 43764 7980
rect 43820 7970 43876 7980
rect 43820 7812 43876 7822
rect 43820 7698 43876 7756
rect 43820 7646 43822 7698
rect 43874 7646 43876 7698
rect 43820 7634 43876 7646
rect 43596 7084 43764 7140
rect 43596 5684 43652 7084
rect 43596 5618 43652 5628
rect 43708 6690 43764 6702
rect 43708 6638 43710 6690
rect 43762 6638 43764 6690
rect 43708 6580 43764 6638
rect 43708 5236 43764 6524
rect 43932 6468 43988 11230
rect 44044 8258 44100 11452
rect 44380 11394 44436 11406
rect 44380 11342 44382 11394
rect 44434 11342 44436 11394
rect 44380 11284 44436 11342
rect 44380 11218 44436 11228
rect 44044 8206 44046 8258
rect 44098 8206 44100 8258
rect 44044 8194 44100 8206
rect 44156 11170 44212 11182
rect 44156 11118 44158 11170
rect 44210 11118 44212 11170
rect 44156 8148 44212 11118
rect 44380 9604 44436 9614
rect 44380 9510 44436 9548
rect 44380 8708 44436 8718
rect 44380 8258 44436 8652
rect 44380 8206 44382 8258
rect 44434 8206 44436 8258
rect 44380 8194 44436 8206
rect 44156 8082 44212 8092
rect 44044 8036 44100 8046
rect 44044 7364 44100 7980
rect 44044 7298 44100 7308
rect 44268 7812 44324 7822
rect 44268 7698 44324 7756
rect 44268 7646 44270 7698
rect 44322 7646 44324 7698
rect 44268 7028 44324 7646
rect 44268 6962 44324 6972
rect 44380 7476 44436 7486
rect 44044 6804 44100 6814
rect 44044 6690 44100 6748
rect 44044 6638 44046 6690
rect 44098 6638 44100 6690
rect 44044 6626 44100 6638
rect 44156 6692 44212 6702
rect 43820 6412 43988 6468
rect 44044 6468 44100 6478
rect 43820 6132 43876 6412
rect 43820 6066 43876 6076
rect 43932 6244 43988 6254
rect 43932 6130 43988 6188
rect 43932 6078 43934 6130
rect 43986 6078 43988 6130
rect 43932 6066 43988 6078
rect 43484 5180 43652 5236
rect 43372 3602 43428 3612
rect 43484 5010 43540 5022
rect 43484 4958 43486 5010
rect 43538 4958 43540 5010
rect 43484 3388 43540 4958
rect 43596 4676 43652 5180
rect 43708 5170 43764 5180
rect 43820 5682 43876 5694
rect 43820 5630 43822 5682
rect 43874 5630 43876 5682
rect 43596 4610 43652 4620
rect 43708 4900 43764 4910
rect 43708 4340 43764 4844
rect 43820 4676 43876 5630
rect 44044 5234 44100 6412
rect 44044 5182 44046 5234
rect 44098 5182 44100 5234
rect 44044 5170 44100 5182
rect 43932 4900 43988 4910
rect 43932 4806 43988 4844
rect 44044 4898 44100 4910
rect 44044 4846 44046 4898
rect 44098 4846 44100 4898
rect 43820 4610 43876 4620
rect 44044 4564 44100 4846
rect 44156 4788 44212 6636
rect 44380 6244 44436 7420
rect 44380 6178 44436 6188
rect 44380 6020 44436 6030
rect 44380 5926 44436 5964
rect 44268 5682 44324 5694
rect 44268 5630 44270 5682
rect 44322 5630 44324 5682
rect 44268 4900 44324 5630
rect 44268 4834 44324 4844
rect 44380 5684 44436 5694
rect 44156 4722 44212 4732
rect 43932 4508 44100 4564
rect 44156 4564 44212 4574
rect 44380 4564 44436 5628
rect 44156 4562 44436 4564
rect 44156 4510 44158 4562
rect 44210 4510 44436 4562
rect 44156 4508 44436 4510
rect 43708 4274 43764 4284
rect 43820 4338 43876 4350
rect 43820 4286 43822 4338
rect 43874 4286 43876 4338
rect 43820 4228 43876 4286
rect 43820 4162 43876 4172
rect 43708 4004 43764 4014
rect 43708 3778 43764 3948
rect 43932 3780 43988 4508
rect 44156 4498 44212 4508
rect 44044 4340 44100 4350
rect 44044 4246 44100 4284
rect 44268 4338 44324 4350
rect 44268 4286 44270 4338
rect 44322 4286 44324 4338
rect 44268 3892 44324 4286
rect 44380 4338 44436 4350
rect 44380 4286 44382 4338
rect 44434 4286 44436 4338
rect 44380 4116 44436 4286
rect 44380 4050 44436 4060
rect 44268 3836 44436 3892
rect 43708 3726 43710 3778
rect 43762 3726 43764 3778
rect 43708 3714 43764 3726
rect 43820 3724 43988 3780
rect 43820 3444 43876 3724
rect 44156 3666 44212 3678
rect 44156 3614 44158 3666
rect 44210 3614 44212 3666
rect 43260 2494 43262 2546
rect 43314 2494 43316 2546
rect 43260 2482 43316 2494
rect 43372 3332 43540 3388
rect 43708 3388 43876 3444
rect 43932 3554 43988 3566
rect 43932 3502 43934 3554
rect 43986 3502 43988 3554
rect 43932 3444 43988 3502
rect 44156 3556 44212 3614
rect 44156 3490 44212 3500
rect 44380 3444 44436 3836
rect 44492 3556 44548 11732
rect 44716 10500 44772 12124
rect 44828 11282 44884 11294
rect 44828 11230 44830 11282
rect 44882 11230 44884 11282
rect 44828 10724 44884 11230
rect 44940 11172 44996 11182
rect 45164 11172 45220 11182
rect 44940 11078 44996 11116
rect 45052 11170 45220 11172
rect 45052 11118 45166 11170
rect 45218 11118 45220 11170
rect 45052 11116 45220 11118
rect 44828 10668 44996 10724
rect 44828 10500 44884 10510
rect 44716 10444 44828 10500
rect 44828 10434 44884 10444
rect 44828 10164 44884 10174
rect 44716 8932 44772 8942
rect 44716 8838 44772 8876
rect 44828 8202 44884 10108
rect 44940 8708 44996 10668
rect 45052 8820 45108 11116
rect 45164 11106 45220 11116
rect 45388 11170 45444 11182
rect 45388 11118 45390 11170
rect 45442 11118 45444 11170
rect 45164 10500 45220 10510
rect 45164 9940 45220 10444
rect 45388 10276 45444 11118
rect 45500 11172 45556 12684
rect 45612 12674 45668 12684
rect 45612 12292 45668 12302
rect 45612 12198 45668 12236
rect 45724 11396 45780 11406
rect 45612 11172 45668 11182
rect 45500 11116 45612 11172
rect 45612 11106 45668 11116
rect 45388 10210 45444 10220
rect 45388 9940 45444 9950
rect 45164 9938 45388 9940
rect 45164 9886 45166 9938
rect 45218 9886 45388 9938
rect 45164 9884 45388 9886
rect 45164 9874 45220 9884
rect 45388 9044 45444 9884
rect 45724 9826 45780 11340
rect 45948 11284 46004 11294
rect 45724 9774 45726 9826
rect 45778 9774 45780 9826
rect 45388 9042 45668 9044
rect 45388 8990 45390 9042
rect 45442 8990 45668 9042
rect 45388 8988 45668 8990
rect 45388 8978 45444 8988
rect 45052 8764 45556 8820
rect 44940 8484 44996 8652
rect 45276 8596 45332 8606
rect 44940 8428 45108 8484
rect 45052 8370 45108 8428
rect 45052 8318 45054 8370
rect 45106 8318 45108 8370
rect 45052 8306 45108 8318
rect 45276 8372 45332 8540
rect 45276 8316 45444 8372
rect 44828 8150 44830 8202
rect 44882 8150 44884 8202
rect 44604 8036 44660 8046
rect 44604 6580 44660 7980
rect 44716 7700 44772 7710
rect 44716 7362 44772 7644
rect 44716 7310 44718 7362
rect 44770 7310 44772 7362
rect 44716 7298 44772 7310
rect 44604 6514 44660 6524
rect 44716 7028 44772 7038
rect 44604 6132 44660 6142
rect 44604 3778 44660 6076
rect 44716 4004 44772 6972
rect 44828 6132 44884 8150
rect 45164 8260 45220 8270
rect 45164 8148 45220 8204
rect 45276 8148 45332 8158
rect 45164 8146 45332 8148
rect 45164 8094 45278 8146
rect 45330 8094 45332 8146
rect 45164 8092 45332 8094
rect 45276 8082 45332 8092
rect 45052 8036 45108 8046
rect 45052 7942 45108 7980
rect 45388 7924 45444 8316
rect 45276 7868 45444 7924
rect 45052 7700 45108 7710
rect 44828 6066 44884 6076
rect 44940 6466 44996 6478
rect 44940 6414 44942 6466
rect 44994 6414 44996 6466
rect 44940 5908 44996 6414
rect 44940 5842 44996 5852
rect 44828 5796 44884 5806
rect 44828 5702 44884 5740
rect 45052 5684 45108 7644
rect 44940 5628 45108 5684
rect 45164 6914 45220 6926
rect 45164 6862 45166 6914
rect 45218 6862 45220 6914
rect 44828 5124 44884 5134
rect 44940 5124 44996 5628
rect 44828 5122 44996 5124
rect 44828 5070 44830 5122
rect 44882 5070 44996 5122
rect 44828 5068 44996 5070
rect 45052 5122 45108 5134
rect 45052 5070 45054 5122
rect 45106 5070 45108 5122
rect 44828 5012 44884 5068
rect 44828 4946 44884 4956
rect 44828 4676 44884 4686
rect 45052 4676 45108 5070
rect 44884 4620 45108 4676
rect 44828 4562 44884 4620
rect 44828 4510 44830 4562
rect 44882 4510 44884 4562
rect 44828 4498 44884 4510
rect 45052 4338 45108 4350
rect 45052 4286 45054 4338
rect 45106 4286 45108 4338
rect 44940 4226 44996 4238
rect 44940 4174 44942 4226
rect 44994 4174 44996 4226
rect 44716 3948 44884 4004
rect 44604 3726 44606 3778
rect 44658 3726 44660 3778
rect 44604 3714 44660 3726
rect 44716 3780 44772 3790
rect 44492 3490 44548 3500
rect 43932 3388 44100 3444
rect 43372 2994 43428 3332
rect 43372 2942 43374 2994
rect 43426 2942 43428 2994
rect 43372 1652 43428 2942
rect 43708 2884 43764 3388
rect 44044 3332 44100 3388
rect 44044 3266 44100 3276
rect 44268 3388 44436 3444
rect 43708 2828 43876 2884
rect 43372 1586 43428 1596
rect 43708 2658 43764 2670
rect 43708 2606 43710 2658
rect 43762 2606 43764 2658
rect 43148 914 43204 924
rect 43708 800 43764 2606
rect 43820 1316 43876 2828
rect 44268 1652 44324 3388
rect 44716 3330 44772 3724
rect 44828 3444 44884 3948
rect 44940 3668 44996 4174
rect 44940 3602 44996 3612
rect 44828 3378 44884 3388
rect 44716 3278 44718 3330
rect 44770 3278 44772 3330
rect 44716 2996 44772 3278
rect 44940 3330 44996 3342
rect 44940 3278 44942 3330
rect 44994 3278 44996 3330
rect 44940 3220 44996 3278
rect 45052 3332 45108 4286
rect 45164 3554 45220 6862
rect 45276 5796 45332 7868
rect 45500 6914 45556 8764
rect 45500 6862 45502 6914
rect 45554 6862 45556 6914
rect 45500 6850 45556 6862
rect 45612 6690 45668 8988
rect 45724 7924 45780 9774
rect 45836 9938 45892 9950
rect 45836 9886 45838 9938
rect 45890 9886 45892 9938
rect 45836 9156 45892 9886
rect 45836 9090 45892 9100
rect 45836 8932 45892 8942
rect 45836 8838 45892 8876
rect 45836 8148 45892 8158
rect 45836 8054 45892 8092
rect 45724 7868 45892 7924
rect 45724 7588 45780 7598
rect 45724 7494 45780 7532
rect 45612 6638 45614 6690
rect 45666 6638 45668 6690
rect 45612 6626 45668 6638
rect 45500 6580 45556 6590
rect 45388 5796 45444 5806
rect 45276 5794 45444 5796
rect 45276 5742 45390 5794
rect 45442 5742 45444 5794
rect 45276 5740 45444 5742
rect 45388 5730 45444 5740
rect 45500 5572 45556 6524
rect 45724 6356 45780 6366
rect 45836 6356 45892 7868
rect 45948 6802 46004 11228
rect 45948 6750 45950 6802
rect 46002 6750 46004 6802
rect 45948 6738 46004 6750
rect 45780 6300 45892 6356
rect 45724 6290 45780 6300
rect 45836 5796 45892 5806
rect 45388 5516 45556 5572
rect 45724 5740 45836 5796
rect 45276 5460 45332 5470
rect 45276 4676 45332 5404
rect 45388 5346 45444 5516
rect 45612 5460 45668 5470
rect 45388 5294 45390 5346
rect 45442 5294 45444 5346
rect 45388 5282 45444 5294
rect 45500 5404 45612 5460
rect 45276 4610 45332 4620
rect 45388 4900 45444 4910
rect 45388 4564 45444 4844
rect 45388 4498 45444 4508
rect 45388 4338 45444 4350
rect 45388 4286 45390 4338
rect 45442 4286 45444 4338
rect 45164 3502 45166 3554
rect 45218 3502 45220 3554
rect 45164 3490 45220 3502
rect 45276 4004 45332 4014
rect 45052 3266 45108 3276
rect 44940 3154 44996 3164
rect 45276 3108 45332 3948
rect 45276 3042 45332 3052
rect 45388 3892 45444 4286
rect 44716 2930 44772 2940
rect 44268 1586 44324 1596
rect 44380 2546 44436 2558
rect 44380 2494 44382 2546
rect 44434 2494 44436 2546
rect 43820 1250 43876 1260
rect 44380 800 44436 2494
rect 45052 2548 45108 2558
rect 45052 800 45108 2492
rect 45388 2546 45444 3836
rect 45500 3332 45556 5404
rect 45612 5394 45668 5404
rect 45724 5348 45780 5740
rect 45836 5730 45892 5740
rect 46060 5572 46116 13916
rect 46172 13076 46228 13086
rect 46172 12982 46228 13020
rect 47516 12850 47572 12862
rect 47516 12798 47518 12850
rect 47570 12798 47572 12850
rect 46172 12516 46228 12526
rect 46172 11506 46228 12460
rect 46396 12180 46452 12190
rect 46172 11454 46174 11506
rect 46226 11454 46228 11506
rect 46172 11396 46228 11454
rect 46172 11330 46228 11340
rect 46284 12124 46396 12180
rect 45724 5292 45892 5348
rect 45836 5124 45892 5292
rect 45948 5124 46004 5134
rect 45836 5122 46004 5124
rect 45836 5070 45950 5122
rect 46002 5070 46004 5122
rect 45836 5068 46004 5070
rect 45948 5058 46004 5068
rect 45612 5012 45668 5022
rect 45612 4918 45668 4956
rect 45836 4900 45892 4910
rect 45836 4898 46004 4900
rect 45836 4846 45838 4898
rect 45890 4846 46004 4898
rect 45836 4844 46004 4846
rect 45836 4834 45892 4844
rect 45948 4788 46004 4844
rect 45948 4564 46004 4732
rect 45948 4498 46004 4508
rect 45500 3266 45556 3276
rect 45612 4114 45668 4126
rect 45612 4062 45614 4114
rect 45666 4062 45668 4114
rect 45500 3108 45556 3118
rect 45500 2770 45556 3052
rect 45500 2718 45502 2770
rect 45554 2718 45556 2770
rect 45500 2706 45556 2718
rect 45388 2494 45390 2546
rect 45442 2494 45444 2546
rect 45388 2482 45444 2494
rect 45612 980 45668 4062
rect 46060 4004 46116 5516
rect 46172 10948 46228 10958
rect 46172 5236 46228 10892
rect 46284 5460 46340 12124
rect 46396 12114 46452 12124
rect 47516 12068 47572 12798
rect 48076 12738 48132 12750
rect 48076 12686 48078 12738
rect 48130 12686 48132 12738
rect 48076 12628 48132 12686
rect 47740 12068 47796 12078
rect 47516 12066 47796 12068
rect 47516 12014 47742 12066
rect 47794 12014 47796 12066
rect 47516 12012 47796 12014
rect 47740 12002 47796 12012
rect 47516 11620 47572 11630
rect 46956 11172 47012 11182
rect 46956 11060 47012 11116
rect 46956 11004 47236 11060
rect 46732 10610 46788 10622
rect 46732 10558 46734 10610
rect 46786 10558 46788 10610
rect 46508 10498 46564 10510
rect 46508 10446 46510 10498
rect 46562 10446 46564 10498
rect 46396 8036 46452 8046
rect 46396 7700 46452 7980
rect 46396 7634 46452 7644
rect 46508 7028 46564 10446
rect 46620 9714 46676 9726
rect 46620 9662 46622 9714
rect 46674 9662 46676 9714
rect 46620 8148 46676 9662
rect 46732 8260 46788 10558
rect 46956 10610 47012 10622
rect 46956 10558 46958 10610
rect 47010 10558 47012 10610
rect 46956 10388 47012 10558
rect 46956 10322 47012 10332
rect 47068 10164 47124 10174
rect 47068 9938 47124 10108
rect 47068 9886 47070 9938
rect 47122 9886 47124 9938
rect 47068 9828 47124 9886
rect 47068 9762 47124 9772
rect 47180 9380 47236 11004
rect 47068 9324 47236 9380
rect 46732 8194 46788 8204
rect 46844 8372 46900 8382
rect 46620 8082 46676 8092
rect 46508 6962 46564 6972
rect 46620 7474 46676 7486
rect 46620 7422 46622 7474
rect 46674 7422 46676 7474
rect 46396 6692 46452 6702
rect 46620 6692 46676 7422
rect 46452 6636 46676 6692
rect 46732 7474 46788 7486
rect 46732 7422 46734 7474
rect 46786 7422 46788 7474
rect 46396 6356 46452 6636
rect 46732 6356 46788 7422
rect 46844 7476 46900 8316
rect 47068 7700 47124 9324
rect 47180 9154 47236 9166
rect 47180 9102 47182 9154
rect 47234 9102 47236 9154
rect 47180 8708 47236 9102
rect 47180 8642 47236 8652
rect 47404 8932 47460 8942
rect 47068 7634 47124 7644
rect 47180 8148 47236 8158
rect 47180 7586 47236 8092
rect 47180 7534 47182 7586
rect 47234 7534 47236 7586
rect 47180 7522 47236 7534
rect 47292 7588 47348 7598
rect 46844 7474 47124 7476
rect 46844 7422 46846 7474
rect 46898 7422 47124 7474
rect 46844 7420 47124 7422
rect 46844 7410 46900 7420
rect 47068 6748 47124 7420
rect 47068 6692 47236 6748
rect 47068 6578 47124 6590
rect 47068 6526 47070 6578
rect 47122 6526 47124 6578
rect 47068 6468 47124 6526
rect 47068 6402 47124 6412
rect 46956 6356 47012 6366
rect 46732 6300 46900 6356
rect 46396 6290 46452 6300
rect 46396 6132 46452 6142
rect 46396 5684 46452 6076
rect 46732 6132 46788 6142
rect 46508 6018 46564 6030
rect 46508 5966 46510 6018
rect 46562 5966 46564 6018
rect 46508 5908 46564 5966
rect 46508 5842 46564 5852
rect 46732 5908 46788 6076
rect 46732 5842 46788 5852
rect 46844 5684 46900 6300
rect 46396 5628 46564 5684
rect 46284 5394 46340 5404
rect 46172 5180 46452 5236
rect 46172 4452 46228 4462
rect 46172 4116 46228 4396
rect 46172 4050 46228 4060
rect 45836 3948 46116 4004
rect 45836 3668 45892 3948
rect 46060 3668 46116 3678
rect 45836 3612 46004 3668
rect 45724 3330 45780 3342
rect 45724 3278 45726 3330
rect 45778 3278 45780 3330
rect 45724 3108 45780 3278
rect 45836 3332 45892 3370
rect 45836 3266 45892 3276
rect 45948 3108 46004 3612
rect 45724 3052 46004 3108
rect 46060 2434 46116 3612
rect 46172 3554 46228 3566
rect 46172 3502 46174 3554
rect 46226 3502 46228 3554
rect 46172 3332 46228 3502
rect 46284 3444 46340 3454
rect 46284 3350 46340 3388
rect 46172 3266 46228 3276
rect 46396 2996 46452 5180
rect 46508 5234 46564 5628
rect 46844 5618 46900 5628
rect 46732 5460 46788 5470
rect 46508 5182 46510 5234
rect 46562 5182 46564 5234
rect 46508 5170 46564 5182
rect 46620 5236 46676 5246
rect 46620 4676 46676 5180
rect 46732 4788 46788 5404
rect 46844 5236 46900 5246
rect 46956 5236 47012 6300
rect 47180 6132 47236 6692
rect 47180 5346 47236 6076
rect 47292 5906 47348 7532
rect 47292 5854 47294 5906
rect 47346 5854 47348 5906
rect 47292 5842 47348 5854
rect 47180 5294 47182 5346
rect 47234 5294 47236 5346
rect 47180 5282 47236 5294
rect 46900 5180 47012 5236
rect 46844 5142 46900 5180
rect 47292 4898 47348 4910
rect 47292 4846 47294 4898
rect 47346 4846 47348 4898
rect 46732 4732 46900 4788
rect 46620 4610 46676 4620
rect 46844 4564 46900 4732
rect 46844 4498 46900 4508
rect 46620 4452 46676 4462
rect 46620 4340 46676 4396
rect 46508 4284 46676 4340
rect 46844 4340 46900 4350
rect 47180 4340 47236 4350
rect 46900 4284 47180 4340
rect 46508 3666 46564 4284
rect 46844 4274 46900 4284
rect 47180 4274 47236 4284
rect 46508 3614 46510 3666
rect 46562 3614 46564 3666
rect 46508 3602 46564 3614
rect 46732 4004 46788 4014
rect 46732 3332 46788 3948
rect 47068 4004 47124 4014
rect 46732 3266 46788 3276
rect 46844 3554 46900 3566
rect 46844 3502 46846 3554
rect 46898 3502 46900 3554
rect 46172 2940 46452 2996
rect 46620 3108 46676 3118
rect 46172 2548 46228 2940
rect 46620 2884 46676 3052
rect 46284 2828 46676 2884
rect 46284 2770 46340 2828
rect 46284 2718 46286 2770
rect 46338 2718 46340 2770
rect 46284 2706 46340 2718
rect 46172 2492 46452 2548
rect 46060 2382 46062 2434
rect 46114 2382 46116 2434
rect 46060 2370 46116 2382
rect 45612 914 45668 924
rect 45724 2322 45780 2334
rect 45724 2270 45726 2322
rect 45778 2270 45780 2322
rect 45724 800 45780 2270
rect 45836 980 45892 1018
rect 45836 914 45892 924
rect 46396 800 46452 2492
rect 46844 1428 46900 3502
rect 46956 3444 47012 3454
rect 46956 3330 47012 3388
rect 46956 3278 46958 3330
rect 47010 3278 47012 3330
rect 46956 3266 47012 3278
rect 46844 1362 46900 1372
rect 47068 800 47124 3948
rect 47292 3388 47348 4846
rect 47404 4004 47460 8876
rect 47516 7474 47572 11564
rect 47628 11172 47684 11182
rect 47628 10388 47684 11116
rect 47852 10836 47908 10846
rect 48076 10836 48132 12572
rect 47852 10834 48132 10836
rect 47852 10782 47854 10834
rect 47906 10782 48132 10834
rect 47852 10780 48132 10782
rect 47852 10770 47908 10780
rect 48188 10722 48244 10734
rect 48188 10670 48190 10722
rect 48242 10670 48244 10722
rect 48076 10612 48132 10622
rect 47628 10322 47684 10332
rect 47964 10556 48076 10612
rect 47628 9380 47684 9390
rect 47628 7700 47684 9324
rect 47852 9268 47908 9278
rect 47964 9268 48020 10556
rect 48076 10546 48132 10556
rect 47852 9266 48020 9268
rect 47852 9214 47854 9266
rect 47906 9214 48020 9266
rect 47852 9212 48020 9214
rect 48076 9716 48132 9726
rect 47852 9202 47908 9212
rect 47740 9156 47796 9166
rect 47740 9062 47796 9100
rect 47964 8818 48020 8830
rect 47964 8766 47966 8818
rect 48018 8766 48020 8818
rect 47852 8708 47908 8718
rect 47852 8372 47908 8652
rect 47964 8596 48020 8766
rect 47964 8530 48020 8540
rect 47964 8372 48020 8382
rect 47852 8370 48020 8372
rect 47852 8318 47966 8370
rect 48018 8318 48020 8370
rect 47852 8316 48020 8318
rect 47964 8306 48020 8316
rect 47852 8148 47908 8158
rect 47628 7644 47796 7700
rect 47516 7422 47518 7474
rect 47570 7422 47572 7474
rect 47516 7410 47572 7422
rect 47628 7476 47684 7486
rect 47516 6916 47572 6926
rect 47516 6244 47572 6860
rect 47516 6178 47572 6188
rect 47628 6020 47684 7420
rect 47628 5906 47684 5964
rect 47628 5854 47630 5906
rect 47682 5854 47684 5906
rect 47628 5842 47684 5854
rect 47404 3938 47460 3948
rect 47628 5346 47684 5358
rect 47628 5294 47630 5346
rect 47682 5294 47684 5346
rect 47404 3780 47460 3790
rect 47404 3554 47460 3724
rect 47404 3502 47406 3554
rect 47458 3502 47460 3554
rect 47404 3490 47460 3502
rect 47628 3668 47684 5294
rect 47740 4676 47796 7644
rect 47852 7698 47908 8092
rect 48076 8036 48132 9660
rect 48188 9156 48244 10670
rect 48188 9090 48244 9100
rect 47852 7646 47854 7698
rect 47906 7646 47908 7698
rect 47852 7634 47908 7646
rect 47964 7980 48132 8036
rect 47852 7362 47908 7374
rect 47852 7310 47854 7362
rect 47906 7310 47908 7362
rect 47852 6916 47908 7310
rect 47852 6850 47908 6860
rect 47964 6468 48020 7980
rect 48076 7700 48132 7710
rect 48300 7700 48356 17052
rect 49512 16492 49776 16502
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49512 16426 49776 16436
rect 48524 15876 48580 15886
rect 48412 11282 48468 11294
rect 48412 11230 48414 11282
rect 48466 11230 48468 11282
rect 48412 10500 48468 11230
rect 48412 10434 48468 10444
rect 48412 9604 48468 9614
rect 48412 8372 48468 9548
rect 48412 8306 48468 8316
rect 48300 7644 48468 7700
rect 48076 7606 48132 7644
rect 48188 7474 48244 7486
rect 48188 7422 48190 7474
rect 48242 7422 48244 7474
rect 48188 7140 48244 7422
rect 48188 7074 48244 7084
rect 47740 4610 47796 4620
rect 47852 6412 48020 6468
rect 48076 6578 48132 6590
rect 48076 6526 48078 6578
rect 48130 6526 48132 6578
rect 47628 3444 47684 3612
rect 47740 3444 47796 3454
rect 47628 3442 47796 3444
rect 47628 3390 47742 3442
rect 47794 3390 47796 3442
rect 47628 3388 47796 3390
rect 47180 3332 47348 3388
rect 47740 3378 47796 3388
rect 47180 2994 47236 3332
rect 47852 3220 47908 6412
rect 47964 6244 48020 6254
rect 47964 5010 48020 6188
rect 47964 4958 47966 5010
rect 48018 4958 48020 5010
rect 47964 4946 48020 4958
rect 47964 4564 48020 4574
rect 47964 4450 48020 4508
rect 47964 4398 47966 4450
rect 48018 4398 48020 4450
rect 47964 4386 48020 4398
rect 48076 3444 48132 6526
rect 48300 6020 48356 6030
rect 48188 5794 48244 5806
rect 48188 5742 48190 5794
rect 48242 5742 48244 5794
rect 48188 5124 48244 5742
rect 48188 5058 48244 5068
rect 48300 5122 48356 5964
rect 48300 5070 48302 5122
rect 48354 5070 48356 5122
rect 48300 5058 48356 5070
rect 48188 4676 48244 4686
rect 48244 4620 48356 4676
rect 48188 4610 48244 4620
rect 48076 3378 48132 3388
rect 48300 3388 48356 4620
rect 48412 3666 48468 7644
rect 48524 4564 48580 15820
rect 51436 15540 51492 15550
rect 51436 15148 51492 15484
rect 54236 15316 54292 15326
rect 51436 15092 51716 15148
rect 49512 14924 49776 14934
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49512 14858 49776 14868
rect 49512 13356 49776 13366
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49512 13290 49776 13300
rect 48636 12738 48692 12750
rect 48636 12686 48638 12738
rect 48690 12686 48692 12738
rect 48636 11172 48692 12686
rect 48748 12290 48804 12302
rect 49308 12292 49364 12302
rect 48748 12238 48750 12290
rect 48802 12238 48804 12290
rect 48748 11844 48804 12238
rect 48972 12290 49364 12292
rect 48972 12238 49310 12290
rect 49362 12238 49364 12290
rect 48972 12236 49364 12238
rect 48748 11778 48804 11788
rect 48860 11956 48916 11966
rect 48636 11106 48692 11116
rect 48748 11284 48804 11294
rect 48748 10724 48804 11228
rect 48636 10668 48804 10724
rect 48636 9492 48692 10668
rect 48748 10498 48804 10510
rect 48748 10446 48750 10498
rect 48802 10446 48804 10498
rect 48748 10388 48804 10446
rect 48748 10322 48804 10332
rect 48860 9604 48916 11900
rect 48860 9538 48916 9548
rect 48972 9492 49028 12236
rect 49308 12226 49364 12236
rect 49868 12066 49924 12078
rect 50316 12068 50372 12078
rect 49868 12014 49870 12066
rect 49922 12014 49924 12066
rect 49512 11788 49776 11798
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49512 11722 49776 11732
rect 49868 11788 49924 12014
rect 50204 12012 50316 12068
rect 49868 11732 50036 11788
rect 49644 11508 49700 11518
rect 49868 11508 49924 11732
rect 49196 11506 49924 11508
rect 49196 11454 49646 11506
rect 49698 11454 49924 11506
rect 49196 11452 49924 11454
rect 49196 11394 49252 11452
rect 49644 11442 49700 11452
rect 49196 11342 49198 11394
rect 49250 11342 49252 11394
rect 49196 11330 49252 11342
rect 49196 10610 49252 10622
rect 49196 10558 49198 10610
rect 49250 10558 49252 10610
rect 49196 10164 49252 10558
rect 49756 10500 49812 10510
rect 49756 10406 49812 10444
rect 49196 10098 49252 10108
rect 49308 10388 49364 10398
rect 49308 9938 49364 10332
rect 49512 10220 49776 10230
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49512 10154 49776 10164
rect 49308 9886 49310 9938
rect 49362 9886 49364 9938
rect 49308 9874 49364 9886
rect 49980 9940 50036 11732
rect 49980 9826 50036 9884
rect 49980 9774 49982 9826
rect 50034 9774 50036 9826
rect 49980 9762 50036 9774
rect 50092 11508 50148 11518
rect 48636 9436 48804 9492
rect 48748 8932 48804 9436
rect 48972 9426 49028 9436
rect 49308 9492 49364 9502
rect 48860 9156 48916 9194
rect 48860 9090 48916 9100
rect 48860 8932 48916 8942
rect 48748 8930 48916 8932
rect 48748 8878 48862 8930
rect 48914 8878 48916 8930
rect 48748 8876 48916 8878
rect 48860 8866 48916 8876
rect 49084 8930 49140 8942
rect 49084 8878 49086 8930
rect 49138 8878 49140 8930
rect 48636 8596 48692 8606
rect 48972 8596 49028 8606
rect 48636 8370 48692 8540
rect 48860 8540 48972 8596
rect 48636 8318 48638 8370
rect 48690 8318 48692 8370
rect 48636 8306 48692 8318
rect 48748 8372 48804 8382
rect 48636 8036 48692 8046
rect 48636 7140 48692 7980
rect 48748 7588 48804 8316
rect 48748 7494 48804 7532
rect 48636 7074 48692 7084
rect 48636 6580 48692 6590
rect 48636 5124 48692 6524
rect 48860 6132 48916 8540
rect 48972 8530 49028 8540
rect 49084 7812 49140 8878
rect 49308 8596 49364 9436
rect 50092 9380 50148 11452
rect 49868 9324 50148 9380
rect 49420 9154 49476 9166
rect 49420 9102 49422 9154
rect 49474 9102 49476 9154
rect 49420 8820 49476 9102
rect 49420 8754 49476 8764
rect 49644 9044 49700 9054
rect 49644 8820 49700 8988
rect 49644 8754 49700 8764
rect 49512 8652 49776 8662
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49512 8586 49776 8596
rect 49308 8530 49364 8540
rect 49308 8372 49364 8382
rect 49868 8372 49924 9324
rect 50204 9268 50260 12012
rect 50316 11974 50372 12012
rect 50876 12068 50932 12078
rect 50876 12066 51044 12068
rect 50876 12014 50878 12066
rect 50930 12014 51044 12066
rect 50876 12012 51044 12014
rect 50876 12002 50932 12012
rect 50988 11788 51044 12012
rect 50988 11732 51380 11788
rect 50540 11506 50596 11518
rect 50540 11454 50542 11506
rect 50594 11454 50596 11506
rect 50540 10388 50596 11454
rect 50764 10724 50820 10734
rect 50764 10630 50820 10668
rect 50540 10322 50596 10332
rect 50876 10500 50932 10510
rect 50092 9212 50260 9268
rect 50428 10052 50484 10062
rect 50092 8930 50148 9212
rect 50092 8878 50094 8930
rect 50146 8878 50148 8930
rect 49084 7756 49252 7812
rect 48972 7700 49028 7710
rect 48972 7606 49028 7644
rect 49084 7476 49140 7486
rect 49084 7382 49140 7420
rect 49196 6802 49252 7756
rect 49196 6750 49198 6802
rect 49250 6750 49252 6802
rect 49196 6738 49252 6750
rect 49308 7474 49364 8316
rect 49532 8316 49924 8372
rect 49980 8596 50036 8606
rect 49532 7588 49588 8316
rect 49980 8260 50036 8540
rect 50092 8372 50148 8878
rect 50092 8306 50148 8316
rect 50204 9044 50260 9054
rect 49756 8204 50036 8260
rect 49644 8148 49700 8158
rect 49644 8054 49700 8092
rect 49532 7522 49588 7532
rect 49308 7422 49310 7474
rect 49362 7422 49364 7474
rect 49196 6580 49252 6590
rect 49196 6356 49252 6524
rect 49196 6290 49252 6300
rect 48860 6076 49140 6132
rect 48860 5908 48916 5918
rect 48860 5814 48916 5852
rect 48972 5684 49028 5694
rect 48972 5236 49028 5628
rect 48636 5122 48804 5124
rect 48636 5070 48638 5122
rect 48690 5070 48804 5122
rect 48636 5068 48804 5070
rect 48636 5058 48692 5068
rect 48636 4564 48692 4574
rect 48524 4562 48692 4564
rect 48524 4510 48638 4562
rect 48690 4510 48692 4562
rect 48524 4508 48692 4510
rect 48636 4498 48692 4508
rect 48412 3614 48414 3666
rect 48466 3614 48468 3666
rect 48412 3602 48468 3614
rect 48748 3556 48804 5068
rect 48972 5010 49028 5180
rect 48972 4958 48974 5010
rect 49026 4958 49028 5010
rect 48972 4946 49028 4958
rect 48748 3490 48804 3500
rect 48300 3332 48468 3388
rect 47180 2942 47182 2994
rect 47234 2942 47236 2994
rect 47180 2930 47236 2942
rect 47740 3164 47908 3220
rect 47740 800 47796 3164
rect 48412 800 48468 3332
rect 49084 800 49140 6076
rect 49196 5908 49252 5918
rect 49196 5572 49252 5852
rect 49196 5506 49252 5516
rect 49308 5794 49364 7422
rect 49756 7364 49812 8204
rect 49980 8036 50036 8046
rect 49756 7298 49812 7308
rect 49868 7588 49924 7598
rect 49512 7084 49776 7094
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49512 7018 49776 7028
rect 49868 6748 49924 7532
rect 49308 5742 49310 5794
rect 49362 5742 49364 5794
rect 49308 1540 49364 5742
rect 49756 6692 49924 6748
rect 49756 5684 49812 6692
rect 49756 5618 49812 5628
rect 49868 6466 49924 6478
rect 49868 6414 49870 6466
rect 49922 6414 49924 6466
rect 49512 5516 49776 5526
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49512 5450 49776 5460
rect 49644 5348 49700 5358
rect 49420 4898 49476 4910
rect 49420 4846 49422 4898
rect 49474 4846 49476 4898
rect 49420 4228 49476 4846
rect 49644 4788 49700 5292
rect 49868 5124 49924 6414
rect 49756 5068 49924 5124
rect 49756 5012 49812 5068
rect 49756 4946 49812 4956
rect 49868 4898 49924 4910
rect 49868 4846 49870 4898
rect 49922 4846 49924 4898
rect 49868 4788 49924 4846
rect 49644 4732 49924 4788
rect 49420 4162 49476 4172
rect 49512 3948 49776 3958
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49512 3882 49776 3892
rect 49980 3780 50036 7980
rect 50092 7476 50148 7486
rect 50092 7362 50148 7420
rect 50092 7310 50094 7362
rect 50146 7310 50148 7362
rect 50092 7298 50148 7310
rect 50204 6802 50260 8988
rect 50428 8484 50484 9996
rect 50764 9714 50820 9726
rect 50764 9662 50766 9714
rect 50818 9662 50820 9714
rect 50540 9602 50596 9614
rect 50540 9550 50542 9602
rect 50594 9550 50596 9602
rect 50540 9492 50596 9550
rect 50540 9426 50596 9436
rect 50652 9602 50708 9614
rect 50652 9550 50654 9602
rect 50706 9550 50708 9602
rect 50652 9156 50708 9550
rect 50652 9090 50708 9100
rect 50764 9044 50820 9662
rect 50764 8978 50820 8988
rect 50764 8708 50820 8718
rect 50316 8428 50484 8484
rect 50652 8652 50764 8708
rect 50316 6914 50372 8428
rect 50428 8260 50484 8270
rect 50652 8260 50708 8652
rect 50764 8642 50820 8652
rect 50428 8166 50484 8204
rect 50540 8204 50708 8260
rect 50764 8370 50820 8382
rect 50764 8318 50766 8370
rect 50818 8318 50820 8370
rect 50316 6862 50318 6914
rect 50370 6862 50372 6914
rect 50316 6850 50372 6862
rect 50204 6750 50206 6802
rect 50258 6750 50260 6802
rect 50204 6738 50260 6750
rect 49644 3724 50036 3780
rect 50092 6690 50148 6702
rect 50092 6638 50094 6690
rect 50146 6638 50148 6690
rect 49644 3442 49700 3724
rect 50092 3668 50148 6638
rect 50204 6578 50260 6590
rect 50204 6526 50206 6578
rect 50258 6526 50260 6578
rect 50204 5794 50260 6526
rect 50204 5742 50206 5794
rect 50258 5742 50260 5794
rect 50204 5730 50260 5742
rect 50316 6466 50372 6478
rect 50316 6414 50318 6466
rect 50370 6414 50372 6466
rect 50204 5572 50260 5582
rect 50204 5124 50260 5516
rect 50316 5348 50372 6414
rect 50316 5282 50372 5292
rect 50316 5124 50372 5134
rect 50204 5122 50372 5124
rect 50204 5070 50318 5122
rect 50370 5070 50372 5122
rect 50204 5068 50372 5070
rect 50316 5058 50372 5068
rect 49644 3390 49646 3442
rect 49698 3390 49700 3442
rect 49644 3378 49700 3390
rect 49756 3612 50148 3668
rect 50316 4900 50372 4910
rect 49308 1474 49364 1484
rect 49756 800 49812 3612
rect 50204 3332 50260 3342
rect 50204 3238 50260 3276
rect 50316 2884 50372 4844
rect 50540 3892 50596 8204
rect 50652 8034 50708 8046
rect 50652 7982 50654 8034
rect 50706 7982 50708 8034
rect 50652 7700 50708 7982
rect 50652 7634 50708 7644
rect 50764 7364 50820 8318
rect 50764 7298 50820 7308
rect 50540 3826 50596 3836
rect 50652 6692 50708 6702
rect 50428 3556 50484 3594
rect 50428 3490 50484 3500
rect 50652 3388 50708 6636
rect 50316 2818 50372 2828
rect 50428 3332 50708 3388
rect 50764 6692 50820 6702
rect 50876 6692 50932 10444
rect 51324 9940 51380 11732
rect 51548 11284 51604 11294
rect 51548 11190 51604 11228
rect 51548 10722 51604 10734
rect 51548 10670 51550 10722
rect 51602 10670 51604 10722
rect 51548 10052 51604 10670
rect 51548 9986 51604 9996
rect 51100 9602 51156 9614
rect 51100 9550 51102 9602
rect 51154 9550 51156 9602
rect 50764 6690 50932 6692
rect 50764 6638 50766 6690
rect 50818 6638 50932 6690
rect 50764 6636 50932 6638
rect 50988 9268 51044 9278
rect 50988 6692 51044 9212
rect 51100 8820 51156 9550
rect 51100 8754 51156 8764
rect 51100 8484 51156 8494
rect 51156 8428 51268 8484
rect 51100 8418 51156 8428
rect 50204 1764 50260 1774
rect 50204 1092 50260 1708
rect 50204 1026 50260 1036
rect 50428 800 50484 3332
rect 50764 2772 50820 6636
rect 50988 6626 51044 6636
rect 51100 6690 51156 6702
rect 51100 6638 51102 6690
rect 51154 6638 51156 6690
rect 50988 6468 51044 6478
rect 50988 6374 51044 6412
rect 50988 6244 51044 6254
rect 50764 2706 50820 2716
rect 50876 5684 50932 5694
rect 50876 2322 50932 5628
rect 50988 4450 51044 6188
rect 51100 6132 51156 6638
rect 51100 6066 51156 6076
rect 51100 5010 51156 5022
rect 51100 4958 51102 5010
rect 51154 4958 51156 5010
rect 51100 4676 51156 4958
rect 51100 4610 51156 4620
rect 50988 4398 50990 4450
rect 51042 4398 51044 4450
rect 50988 4386 51044 4398
rect 51212 3442 51268 8428
rect 51324 8036 51380 9884
rect 51548 9602 51604 9614
rect 51548 9550 51550 9602
rect 51602 9550 51604 9602
rect 51548 8932 51604 9550
rect 51548 8866 51604 8876
rect 51548 8596 51604 8606
rect 51548 8370 51604 8540
rect 51548 8318 51550 8370
rect 51602 8318 51604 8370
rect 51548 8306 51604 8318
rect 51324 7970 51380 7980
rect 51660 7700 51716 15092
rect 53228 13188 53284 13198
rect 53284 13132 53396 13188
rect 53228 13122 53284 13132
rect 52332 11060 52388 11070
rect 52388 11004 52500 11060
rect 52332 10994 52388 11004
rect 51996 10724 52052 10734
rect 51548 7644 51716 7700
rect 51772 10722 52052 10724
rect 51772 10670 51998 10722
rect 52050 10670 52052 10722
rect 51772 10668 52052 10670
rect 51324 7364 51380 7374
rect 51380 7308 51492 7364
rect 51324 7298 51380 7308
rect 51436 6690 51492 7308
rect 51436 6638 51438 6690
rect 51490 6638 51492 6690
rect 51436 6626 51492 6638
rect 51548 6692 51604 7644
rect 51772 7588 51828 10668
rect 51996 10658 52052 10668
rect 51996 10164 52052 10174
rect 51884 10108 51996 10164
rect 51884 8484 51940 10108
rect 51996 10098 52052 10108
rect 51996 9716 52052 9726
rect 51996 9602 52052 9660
rect 51996 9550 51998 9602
rect 52050 9550 52052 9602
rect 51996 9538 52052 9550
rect 52220 8932 52276 8942
rect 52220 8838 52276 8876
rect 52220 8484 52276 8494
rect 51884 8428 52052 8484
rect 51996 8372 52052 8428
rect 51996 8316 52164 8372
rect 51884 8260 51940 8270
rect 51884 8166 51940 8204
rect 51996 8146 52052 8158
rect 51996 8094 51998 8146
rect 52050 8094 52052 8146
rect 51548 6626 51604 6636
rect 51660 7532 51828 7588
rect 51884 8036 51940 8046
rect 51548 6466 51604 6478
rect 51548 6414 51550 6466
rect 51602 6414 51604 6466
rect 51324 6020 51380 6030
rect 51548 6020 51604 6414
rect 51324 6018 51604 6020
rect 51324 5966 51326 6018
rect 51378 5966 51604 6018
rect 51324 5964 51604 5966
rect 51324 5954 51380 5964
rect 51660 5796 51716 7532
rect 51772 7364 51828 7374
rect 51772 6802 51828 7308
rect 51772 6750 51774 6802
rect 51826 6750 51828 6802
rect 51772 6738 51828 6750
rect 51212 3390 51214 3442
rect 51266 3390 51268 3442
rect 51212 3378 51268 3390
rect 51324 5740 51716 5796
rect 51772 6468 51828 6478
rect 50876 2270 50878 2322
rect 50930 2270 50932 2322
rect 50876 2258 50932 2270
rect 51324 1764 51380 5740
rect 51660 5572 51716 5582
rect 51660 4564 51716 5516
rect 51436 4562 51716 4564
rect 51436 4510 51662 4562
rect 51714 4510 51716 4562
rect 51436 4508 51716 4510
rect 51436 1876 51492 4508
rect 51660 4498 51716 4508
rect 51772 5236 51828 6412
rect 51884 6244 51940 7980
rect 51996 7700 52052 8094
rect 51996 7634 52052 7644
rect 52108 7476 52164 8316
rect 51884 6178 51940 6188
rect 51996 7420 52164 7476
rect 51884 5796 51940 5806
rect 51884 5702 51940 5740
rect 51996 5572 52052 7420
rect 52108 6804 52164 6814
rect 52108 6710 52164 6748
rect 51996 5506 52052 5516
rect 52108 5682 52164 5694
rect 52108 5630 52110 5682
rect 52162 5630 52164 5682
rect 51772 4562 51828 5180
rect 51772 4510 51774 4562
rect 51826 4510 51828 4562
rect 51772 4498 51828 4510
rect 51996 5348 52052 5358
rect 51548 3892 51604 3902
rect 51604 3836 51828 3892
rect 51548 3826 51604 3836
rect 51548 3332 51604 3342
rect 51548 3238 51604 3276
rect 51436 1810 51492 1820
rect 51100 1708 51380 1764
rect 51100 800 51156 1708
rect 51772 800 51828 3836
rect 51884 3666 51940 3678
rect 51884 3614 51886 3666
rect 51938 3614 51940 3666
rect 51884 2436 51940 3614
rect 51996 3442 52052 5292
rect 52108 5234 52164 5630
rect 52220 5348 52276 8428
rect 52332 8372 52388 8382
rect 52332 7586 52388 8316
rect 52332 7534 52334 7586
rect 52386 7534 52388 7586
rect 52332 7522 52388 7534
rect 52444 7028 52500 11004
rect 52556 10500 52612 10510
rect 52556 10406 52612 10444
rect 53004 10498 53060 10510
rect 53004 10446 53006 10498
rect 53058 10446 53060 10498
rect 52668 10386 52724 10398
rect 52668 10334 52670 10386
rect 52722 10334 52724 10386
rect 52668 10276 52724 10334
rect 52556 10220 52724 10276
rect 52556 9380 52612 10220
rect 53004 10164 53060 10446
rect 53004 10098 53060 10108
rect 53004 9828 53060 9838
rect 52668 9604 52724 9614
rect 52668 9510 52724 9548
rect 52556 8036 52612 9324
rect 52892 9492 52948 9502
rect 52556 7970 52612 7980
rect 52668 8146 52724 8158
rect 52668 8094 52670 8146
rect 52722 8094 52724 8146
rect 52444 6972 52612 7028
rect 52332 6916 52388 6926
rect 52332 6132 52388 6860
rect 52556 6914 52612 6972
rect 52556 6862 52558 6914
rect 52610 6862 52612 6914
rect 52556 6850 52612 6862
rect 52332 6130 52612 6132
rect 52332 6078 52334 6130
rect 52386 6078 52612 6130
rect 52332 6076 52612 6078
rect 52332 6066 52388 6076
rect 52556 5348 52612 6076
rect 52668 5682 52724 8094
rect 52892 8146 52948 9436
rect 53004 9044 53060 9772
rect 53116 9602 53172 9614
rect 53116 9550 53118 9602
rect 53170 9550 53172 9602
rect 53116 9268 53172 9550
rect 53116 9202 53172 9212
rect 53004 9042 53284 9044
rect 53004 8990 53006 9042
rect 53058 8990 53284 9042
rect 53004 8988 53284 8990
rect 53004 8978 53060 8988
rect 53228 8818 53284 8988
rect 53228 8766 53230 8818
rect 53282 8766 53284 8818
rect 52892 8094 52894 8146
rect 52946 8094 52948 8146
rect 52892 8082 52948 8094
rect 53004 8370 53060 8382
rect 53004 8318 53006 8370
rect 53058 8318 53060 8370
rect 53004 8148 53060 8318
rect 53004 8082 53060 8092
rect 53228 7924 53284 8766
rect 53004 7868 53284 7924
rect 53004 7474 53060 7868
rect 53340 7812 53396 13132
rect 53788 10948 53844 10958
rect 53564 10498 53620 10510
rect 53564 10446 53566 10498
rect 53618 10446 53620 10498
rect 53564 10386 53620 10446
rect 53564 10334 53566 10386
rect 53618 10334 53620 10386
rect 53564 10322 53620 10334
rect 53564 9602 53620 9614
rect 53564 9550 53566 9602
rect 53618 9550 53620 9602
rect 53452 8930 53508 8942
rect 53452 8878 53454 8930
rect 53506 8878 53508 8930
rect 53452 8818 53508 8878
rect 53452 8766 53454 8818
rect 53506 8766 53508 8818
rect 53452 8754 53508 8766
rect 53564 8708 53620 9550
rect 53564 8642 53620 8652
rect 53676 9604 53732 9614
rect 53340 7756 53620 7812
rect 53228 7700 53284 7710
rect 53004 7422 53006 7474
rect 53058 7422 53060 7474
rect 53004 7410 53060 7422
rect 53116 7644 53228 7700
rect 52780 6914 52836 6926
rect 52780 6862 52782 6914
rect 52834 6862 52836 6914
rect 52780 6804 52836 6862
rect 52892 6804 52948 6814
rect 52780 6802 52948 6804
rect 52780 6750 52894 6802
rect 52946 6750 52948 6802
rect 52780 6748 52948 6750
rect 52892 6738 52948 6748
rect 52668 5630 52670 5682
rect 52722 5630 52724 5682
rect 52668 5618 52724 5630
rect 52780 5794 52836 5806
rect 52780 5742 52782 5794
rect 52834 5742 52836 5794
rect 52780 5572 52836 5742
rect 53116 5684 53172 7644
rect 53228 7634 53284 7644
rect 53452 7586 53508 7598
rect 53452 7534 53454 7586
rect 53506 7534 53508 7586
rect 53228 5908 53284 5918
rect 53228 5814 53284 5852
rect 53452 5684 53508 7534
rect 53116 5628 53284 5684
rect 52780 5506 52836 5516
rect 52668 5348 52724 5358
rect 52556 5346 52724 5348
rect 52556 5294 52670 5346
rect 52722 5294 52724 5346
rect 52556 5292 52724 5294
rect 52220 5282 52276 5292
rect 52108 5182 52110 5234
rect 52162 5182 52164 5234
rect 52108 5170 52164 5182
rect 52220 5124 52276 5134
rect 52220 4450 52276 5068
rect 52444 4788 52500 4798
rect 52332 4676 52388 4686
rect 52332 4562 52388 4620
rect 52332 4510 52334 4562
rect 52386 4510 52388 4562
rect 52332 4498 52388 4510
rect 52220 4398 52222 4450
rect 52274 4398 52276 4450
rect 52220 4386 52276 4398
rect 51996 3390 51998 3442
rect 52050 3390 52052 3442
rect 51996 3378 52052 3390
rect 52108 4338 52164 4350
rect 52108 4286 52110 4338
rect 52162 4286 52164 4338
rect 52108 2996 52164 4286
rect 52220 3668 52276 3678
rect 52220 3574 52276 3612
rect 52108 2930 52164 2940
rect 51884 2370 51940 2380
rect 52444 800 52500 4732
rect 52668 4676 52724 5292
rect 52668 4610 52724 4620
rect 52780 5348 52836 5358
rect 52668 4340 52724 4350
rect 52556 4228 52612 4238
rect 52556 4134 52612 4172
rect 52556 3668 52612 3678
rect 52556 3574 52612 3612
rect 52668 3666 52724 4284
rect 52780 4338 52836 5292
rect 53228 5234 53284 5628
rect 53452 5618 53508 5628
rect 53228 5182 53230 5234
rect 53282 5182 53284 5234
rect 53228 5170 53284 5182
rect 53452 5236 53508 5246
rect 53452 5142 53508 5180
rect 52780 4286 52782 4338
rect 52834 4286 52836 4338
rect 52780 4274 52836 4286
rect 53004 5122 53060 5134
rect 53004 5070 53006 5122
rect 53058 5070 53060 5122
rect 53004 4340 53060 5070
rect 53004 4274 53060 4284
rect 53116 5012 53172 5022
rect 53564 5012 53620 7756
rect 52668 3614 52670 3666
rect 52722 3614 52724 3666
rect 52668 3602 52724 3614
rect 53004 4004 53060 4014
rect 52892 3556 52948 3566
rect 53004 3556 53060 3948
rect 52892 3554 53060 3556
rect 52892 3502 52894 3554
rect 52946 3502 53060 3554
rect 52892 3500 53060 3502
rect 52892 3490 52948 3500
rect 53116 800 53172 4956
rect 53228 4956 53620 5012
rect 53228 3666 53284 4956
rect 53340 4564 53396 4574
rect 53340 4338 53396 4508
rect 53340 4286 53342 4338
rect 53394 4286 53396 4338
rect 53340 4274 53396 4286
rect 53228 3614 53230 3666
rect 53282 3614 53284 3666
rect 53228 3602 53284 3614
rect 53340 4116 53396 4126
rect 53340 2660 53396 4060
rect 53564 4116 53620 4126
rect 53564 4022 53620 4060
rect 53676 4004 53732 9548
rect 53788 8820 53844 10892
rect 54012 10500 54068 10510
rect 54012 10406 54068 10444
rect 54012 9604 54068 9614
rect 54012 9602 54180 9604
rect 54012 9550 54014 9602
rect 54066 9550 54180 9602
rect 54012 9548 54180 9550
rect 54012 9538 54068 9548
rect 53900 9044 53956 9054
rect 53900 8950 53956 8988
rect 53788 8764 53956 8820
rect 53788 8372 53844 8382
rect 53788 8278 53844 8316
rect 53676 3938 53732 3948
rect 53788 8036 53844 8046
rect 53676 3668 53732 3678
rect 53676 3574 53732 3612
rect 53564 3554 53620 3566
rect 53564 3502 53566 3554
rect 53618 3502 53620 3554
rect 53564 3444 53620 3502
rect 53676 3444 53732 3454
rect 53564 3388 53676 3444
rect 53676 3378 53732 3388
rect 53340 2594 53396 2604
rect 53788 800 53844 7980
rect 53900 7698 53956 8764
rect 54124 8708 54180 9548
rect 53900 7646 53902 7698
rect 53954 7646 53956 7698
rect 53900 7634 53956 7646
rect 54012 8652 54180 8708
rect 53900 6692 53956 6702
rect 53900 6130 53956 6636
rect 53900 6078 53902 6130
rect 53954 6078 53956 6130
rect 53900 6066 53956 6078
rect 54012 4788 54068 8652
rect 54236 7476 54292 15260
rect 54572 9940 54628 18508
rect 68832 18060 69096 18070
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 68832 17994 69096 18004
rect 67116 17444 67172 17454
rect 59172 17276 59436 17286
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59172 17210 59436 17220
rect 56028 16996 56084 17006
rect 56028 15148 56084 16940
rect 59172 15708 59436 15718
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59172 15642 59436 15652
rect 57372 15428 57428 15438
rect 56028 15092 56532 15148
rect 55692 13636 55748 13646
rect 54460 9938 54628 9940
rect 54460 9886 54574 9938
rect 54626 9886 54628 9938
rect 54460 9884 54628 9886
rect 54348 8932 54404 8942
rect 54348 8838 54404 8876
rect 54348 7700 54404 7710
rect 54348 7606 54404 7644
rect 54460 7586 54516 9884
rect 54572 9874 54628 9884
rect 54684 10500 54740 10510
rect 54684 9828 54740 10444
rect 54460 7534 54462 7586
rect 54514 7534 54516 7586
rect 54460 7522 54516 7534
rect 54572 8596 54628 8606
rect 54012 4722 54068 4732
rect 54124 7420 54292 7476
rect 54124 4564 54180 7420
rect 54572 7140 54628 8540
rect 54236 7084 54628 7140
rect 54236 6018 54292 7084
rect 54236 5966 54238 6018
rect 54290 5966 54292 6018
rect 54236 5954 54292 5966
rect 54460 6916 54516 6926
rect 54124 4498 54180 4508
rect 54236 5796 54292 5806
rect 53900 4340 53956 4350
rect 53900 4246 53956 4284
rect 54236 4116 54292 5740
rect 54236 4050 54292 4060
rect 54348 5572 54404 5582
rect 54348 4562 54404 5516
rect 54348 4510 54350 4562
rect 54402 4510 54404 4562
rect 54348 2546 54404 4510
rect 54348 2494 54350 2546
rect 54402 2494 54404 2546
rect 54348 2482 54404 2494
rect 54460 800 54516 6860
rect 54572 6018 54628 6030
rect 54572 5966 54574 6018
rect 54626 5966 54628 6018
rect 54572 3668 54628 5966
rect 54684 5796 54740 9772
rect 54908 10500 54964 10510
rect 54796 8260 54852 8270
rect 54796 7700 54852 8204
rect 54796 5906 54852 7644
rect 54796 5854 54798 5906
rect 54850 5854 54852 5906
rect 54796 5842 54852 5854
rect 54684 5730 54740 5740
rect 54572 3602 54628 3612
rect 54684 5236 54740 5246
rect 54572 3332 54628 3342
rect 54684 3332 54740 5180
rect 54796 4900 54852 4910
rect 54796 4338 54852 4844
rect 54908 4788 54964 10444
rect 55020 9604 55076 9614
rect 55020 9510 55076 9548
rect 55468 9156 55524 9166
rect 55468 9062 55524 9100
rect 55356 9044 55412 9054
rect 55020 8148 55076 8158
rect 55244 8148 55300 8158
rect 55020 8146 55244 8148
rect 55020 8094 55022 8146
rect 55074 8094 55244 8146
rect 55020 8092 55244 8094
rect 55020 8082 55076 8092
rect 55244 8082 55300 8092
rect 55132 7474 55188 7486
rect 55132 7422 55134 7474
rect 55186 7422 55188 7474
rect 55132 6020 55188 7422
rect 55356 6578 55412 8988
rect 55468 8036 55524 8046
rect 55468 8034 55636 8036
rect 55468 7982 55470 8034
rect 55522 7982 55636 8034
rect 55468 7980 55636 7982
rect 55468 7970 55524 7980
rect 55468 7700 55524 7710
rect 55468 7606 55524 7644
rect 55356 6526 55358 6578
rect 55410 6526 55412 6578
rect 55356 6514 55412 6526
rect 55468 6020 55524 6030
rect 54908 4722 54964 4732
rect 55020 6018 55524 6020
rect 55020 5966 55470 6018
rect 55522 5966 55524 6018
rect 55020 5964 55524 5966
rect 54796 4286 54798 4338
rect 54850 4286 54852 4338
rect 54796 4274 54852 4286
rect 54908 4340 54964 4350
rect 55020 4340 55076 5964
rect 55468 5954 55524 5964
rect 54964 4284 55076 4340
rect 55244 5796 55300 5806
rect 55244 4338 55300 5740
rect 55580 5236 55636 7980
rect 55692 6914 55748 13580
rect 56252 13524 56308 13534
rect 56140 8932 56196 8942
rect 55804 8260 55860 8270
rect 55804 7924 55860 8204
rect 56028 8148 56084 8158
rect 55916 8036 55972 8046
rect 55916 7942 55972 7980
rect 55804 7858 55860 7868
rect 55804 7586 55860 7598
rect 55804 7534 55806 7586
rect 55858 7534 55860 7586
rect 55804 7476 55860 7534
rect 55804 7410 55860 7420
rect 55692 6862 55694 6914
rect 55746 6862 55748 6914
rect 55692 6850 55748 6862
rect 56028 7028 56084 8092
rect 56028 6580 56084 6972
rect 55804 6524 56084 6580
rect 55804 5906 55860 6524
rect 55804 5854 55806 5906
rect 55858 5854 55860 5906
rect 55804 5842 55860 5854
rect 56028 5908 56084 5918
rect 56140 5908 56196 8876
rect 56028 5906 56196 5908
rect 56028 5854 56030 5906
rect 56082 5854 56196 5906
rect 56028 5852 56196 5854
rect 55916 5796 55972 5806
rect 55916 5702 55972 5740
rect 55916 5572 55972 5582
rect 55468 5180 55636 5236
rect 55692 5348 55748 5358
rect 55468 5012 55524 5180
rect 55468 4946 55524 4956
rect 55244 4286 55246 4338
rect 55298 4286 55300 4338
rect 54908 3444 54964 4284
rect 55244 4274 55300 4286
rect 55356 4788 55412 4798
rect 55020 4116 55076 4154
rect 55020 4050 55076 4060
rect 55020 3892 55076 3902
rect 55020 3668 55076 3836
rect 55020 3612 55188 3668
rect 55020 3444 55076 3454
rect 54908 3442 55076 3444
rect 54908 3390 55022 3442
rect 55074 3390 55076 3442
rect 54908 3388 55076 3390
rect 55020 3378 55076 3388
rect 54572 3330 54740 3332
rect 54572 3278 54574 3330
rect 54626 3278 54740 3330
rect 54572 3276 54740 3278
rect 54572 2434 54628 3276
rect 54572 2382 54574 2434
rect 54626 2382 54628 2434
rect 54572 2370 54628 2382
rect 55132 800 55188 3612
rect 55356 3554 55412 4732
rect 55468 4676 55524 4686
rect 55692 4676 55748 5292
rect 55916 5010 55972 5516
rect 56028 5460 56084 5852
rect 56028 5394 56084 5404
rect 56252 5346 56308 13468
rect 56364 8034 56420 8046
rect 56364 7982 56366 8034
rect 56418 7982 56420 8034
rect 56364 6916 56420 7982
rect 56364 6850 56420 6860
rect 56252 5294 56254 5346
rect 56306 5294 56308 5346
rect 56252 5282 56308 5294
rect 56364 5796 56420 5806
rect 55916 4958 55918 5010
rect 55970 4958 55972 5010
rect 55916 4946 55972 4958
rect 56140 5124 56196 5134
rect 55524 4620 55748 4676
rect 55468 4450 55524 4620
rect 56140 4564 56196 5068
rect 56140 4498 56196 4508
rect 56252 4788 56308 4798
rect 55468 4398 55470 4450
rect 55522 4398 55524 4450
rect 55468 4386 55524 4398
rect 55804 4450 55860 4462
rect 55804 4398 55806 4450
rect 55858 4398 55860 4450
rect 55468 4116 55524 4126
rect 55468 3666 55524 4060
rect 55468 3614 55470 3666
rect 55522 3614 55524 3666
rect 55468 3602 55524 3614
rect 55356 3502 55358 3554
rect 55410 3502 55412 3554
rect 55356 3444 55412 3502
rect 55356 3378 55412 3388
rect 55692 3554 55748 3566
rect 55692 3502 55694 3554
rect 55746 3502 55748 3554
rect 55692 2772 55748 3502
rect 55692 2706 55748 2716
rect 55804 2100 55860 4398
rect 55916 3668 55972 3678
rect 55916 3574 55972 3612
rect 56252 3554 56308 4732
rect 56252 3502 56254 3554
rect 56306 3502 56308 3554
rect 56252 3490 56308 3502
rect 56364 3388 56420 5740
rect 56476 4228 56532 15092
rect 56588 8932 56644 8942
rect 56812 8932 56868 8942
rect 56644 8930 56868 8932
rect 56644 8878 56814 8930
rect 56866 8878 56868 8930
rect 56644 8876 56868 8878
rect 56588 8866 56644 8876
rect 56812 8866 56868 8876
rect 57148 8932 57204 8942
rect 57148 8838 57204 8876
rect 56700 8708 56756 8718
rect 56588 7700 56644 7710
rect 56588 7606 56644 7644
rect 56700 7588 56756 8652
rect 56588 7028 56644 7038
rect 56588 4452 56644 6972
rect 56700 6130 56756 7532
rect 56700 6078 56702 6130
rect 56754 6078 56756 6130
rect 56700 6066 56756 6078
rect 56812 8034 56868 8046
rect 57260 8036 57316 8046
rect 56812 7982 56814 8034
rect 56866 7982 56868 8034
rect 56812 4676 56868 7982
rect 57148 8034 57316 8036
rect 57148 7982 57262 8034
rect 57314 7982 57316 8034
rect 57148 7980 57316 7982
rect 56924 7588 56980 7598
rect 56924 7494 56980 7532
rect 57036 7476 57092 7486
rect 56924 6916 56980 6926
rect 56924 4900 56980 6860
rect 56924 4834 56980 4844
rect 56812 4620 56980 4676
rect 56812 4452 56868 4462
rect 56588 4450 56868 4452
rect 56588 4398 56814 4450
rect 56866 4398 56868 4450
rect 56588 4396 56868 4398
rect 56812 4386 56868 4396
rect 56700 4228 56756 4238
rect 56476 4226 56756 4228
rect 56476 4174 56702 4226
rect 56754 4174 56756 4226
rect 56476 4172 56756 4174
rect 56700 4162 56756 4172
rect 56924 3892 56980 4620
rect 56924 3826 56980 3836
rect 57036 4450 57092 7420
rect 57036 4398 57038 4450
rect 57090 4398 57092 4450
rect 55692 2044 55860 2100
rect 56028 3330 56084 3342
rect 56028 3278 56030 3330
rect 56082 3278 56084 3330
rect 55692 980 55748 2044
rect 55692 914 55748 924
rect 55804 1764 55860 1774
rect 55804 800 55860 1708
rect 56028 1316 56084 3278
rect 56140 3332 56420 3388
rect 56476 3780 56532 3790
rect 56140 1652 56196 3332
rect 56140 1586 56196 1596
rect 56028 1250 56084 1260
rect 56476 800 56532 3724
rect 56924 3668 56980 3678
rect 57036 3668 57092 4398
rect 57148 3780 57204 7980
rect 57260 7970 57316 7980
rect 57372 7812 57428 15372
rect 59172 14140 59436 14150
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59172 14074 59436 14084
rect 59172 12572 59436 12582
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59172 12506 59436 12516
rect 58828 12180 58884 12190
rect 58044 11956 58100 11966
rect 57708 11844 57764 11854
rect 57596 11788 57708 11844
rect 57260 7756 57428 7812
rect 57484 10164 57540 10174
rect 57260 7586 57316 7756
rect 57484 7700 57540 10108
rect 57260 7534 57262 7586
rect 57314 7534 57316 7586
rect 57260 7522 57316 7534
rect 57372 7644 57540 7700
rect 57260 7140 57316 7150
rect 57260 6244 57316 7084
rect 57372 6916 57428 7644
rect 57484 7476 57540 7514
rect 57484 7410 57540 7420
rect 57372 6860 57540 6916
rect 57260 6188 57428 6244
rect 57260 6020 57316 6030
rect 57260 3892 57316 5964
rect 57260 3826 57316 3836
rect 57148 3714 57204 3724
rect 57372 3668 57428 6188
rect 57484 5796 57540 6860
rect 57596 6020 57652 11788
rect 57708 11778 57764 11788
rect 57820 8932 57876 8942
rect 57708 7474 57764 7486
rect 57708 7422 57710 7474
rect 57762 7422 57764 7474
rect 57708 6468 57764 7422
rect 57820 6916 57876 8876
rect 57932 8146 57988 8158
rect 57932 8094 57934 8146
rect 57986 8094 57988 8146
rect 57932 7252 57988 8094
rect 57932 7186 57988 7196
rect 57820 6860 57988 6916
rect 57708 6412 57876 6468
rect 57596 5964 57764 6020
rect 57596 5796 57652 5806
rect 57484 5794 57652 5796
rect 57484 5742 57598 5794
rect 57650 5742 57652 5794
rect 57484 5740 57652 5742
rect 57484 4452 57540 5740
rect 57596 5730 57652 5740
rect 57708 5572 57764 5964
rect 57708 5506 57764 5516
rect 57820 5124 57876 6412
rect 57708 5068 57876 5124
rect 57708 4900 57764 5068
rect 57708 4834 57764 4844
rect 57932 4788 57988 6860
rect 58044 6356 58100 11900
rect 58268 10612 58324 10622
rect 58156 10276 58212 10286
rect 58156 6578 58212 10220
rect 58156 6526 58158 6578
rect 58210 6526 58212 6578
rect 58156 6514 58212 6526
rect 58044 6300 58212 6356
rect 57932 4722 57988 4732
rect 58044 6018 58100 6030
rect 58044 5966 58046 6018
rect 58098 5966 58100 6018
rect 57484 4386 57540 4396
rect 57932 4564 57988 4574
rect 57596 4228 57652 4238
rect 56924 3666 57036 3668
rect 56924 3614 56926 3666
rect 56978 3614 57036 3666
rect 56924 3612 57036 3614
rect 56924 3602 56980 3612
rect 57036 3574 57092 3612
rect 57260 3612 57428 3668
rect 57484 4226 57652 4228
rect 57484 4174 57598 4226
rect 57650 4174 57652 4226
rect 57484 4172 57652 4174
rect 57260 3556 57316 3612
rect 57148 3500 57316 3556
rect 56700 3442 56756 3454
rect 56700 3390 56702 3442
rect 56754 3390 56756 3442
rect 56700 2772 56756 3390
rect 56812 3330 56868 3342
rect 56812 3278 56814 3330
rect 56866 3278 56868 3330
rect 56812 3108 56868 3278
rect 56812 3042 56868 3052
rect 56700 2706 56756 2716
rect 57148 800 57204 3500
rect 57372 3442 57428 3454
rect 57372 3390 57374 3442
rect 57426 3390 57428 3442
rect 57372 2324 57428 3390
rect 57484 3220 57540 4172
rect 57596 4162 57652 4172
rect 57820 3780 57876 3790
rect 57596 3668 57652 3678
rect 57596 3574 57652 3612
rect 57484 3154 57540 3164
rect 57372 2258 57428 2268
rect 57820 800 57876 3724
rect 57932 3554 57988 4508
rect 57932 3502 57934 3554
rect 57986 3502 57988 3554
rect 57932 3490 57988 3502
rect 58044 2548 58100 5966
rect 58156 5460 58212 6300
rect 58268 6020 58324 10556
rect 58716 9604 58772 9614
rect 58604 9548 58716 9604
rect 58380 8370 58436 8382
rect 58380 8318 58382 8370
rect 58434 8318 58436 8370
rect 58380 7588 58436 8318
rect 58492 8372 58548 8382
rect 58492 8258 58548 8316
rect 58492 8206 58494 8258
rect 58546 8206 58548 8258
rect 58492 8194 58548 8206
rect 58604 7698 58660 9548
rect 58716 9538 58772 9548
rect 58828 9380 58884 12124
rect 66556 11844 66612 11854
rect 59052 11620 59108 11630
rect 58716 9324 58884 9380
rect 58940 9604 58996 9614
rect 58716 8260 58772 9324
rect 58940 9266 58996 9548
rect 58940 9214 58942 9266
rect 58994 9214 58996 9266
rect 58940 9202 58996 9214
rect 59052 8820 59108 11564
rect 59172 11004 59436 11014
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59172 10938 59436 10948
rect 60844 10948 60900 10958
rect 59500 10836 59556 10846
rect 59172 9436 59436 9446
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59172 9370 59436 9380
rect 59388 9268 59444 9278
rect 59500 9268 59556 10780
rect 59388 9266 59556 9268
rect 59388 9214 59390 9266
rect 59442 9214 59556 9266
rect 59388 9212 59556 9214
rect 59948 9602 60004 9614
rect 59948 9550 59950 9602
rect 60002 9550 60004 9602
rect 59388 9202 59444 9212
rect 59052 8754 59108 8764
rect 59724 8708 59780 8718
rect 59948 8708 60004 9550
rect 60172 9604 60228 9614
rect 60172 9268 60228 9548
rect 60844 9604 60900 10892
rect 62076 10836 62132 10846
rect 61180 9828 61236 9838
rect 60844 9602 61012 9604
rect 60844 9550 60846 9602
rect 60898 9550 61012 9602
rect 60844 9548 61012 9550
rect 60844 9538 60900 9548
rect 60172 9266 60340 9268
rect 60172 9214 60174 9266
rect 60226 9214 60340 9266
rect 60172 9212 60340 9214
rect 60172 9202 60228 9212
rect 59780 8652 60004 8708
rect 60060 8820 60116 8830
rect 59724 8260 59780 8652
rect 58716 8204 58884 8260
rect 58604 7646 58606 7698
rect 58658 7646 58660 7698
rect 58604 7634 58660 7646
rect 58380 7252 58436 7532
rect 58492 7364 58548 7374
rect 58492 7270 58548 7308
rect 58380 6804 58436 7196
rect 58828 7140 58884 8204
rect 59724 8194 59780 8204
rect 59948 8484 60004 8494
rect 59052 8034 59108 8046
rect 59052 7982 59054 8034
rect 59106 7982 59108 8034
rect 58940 7812 58996 7822
rect 59052 7812 59108 7982
rect 59500 8034 59556 8046
rect 59500 7982 59502 8034
rect 59554 7982 59556 8034
rect 59500 7924 59556 7982
rect 58996 7756 59108 7812
rect 59172 7868 59436 7878
rect 59500 7868 59892 7924
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59172 7802 59436 7812
rect 58940 7746 58996 7756
rect 59276 7588 59332 7598
rect 59276 7494 59332 7532
rect 59724 7586 59780 7598
rect 59724 7534 59726 7586
rect 59778 7534 59780 7586
rect 59164 7362 59220 7374
rect 59164 7310 59166 7362
rect 59218 7310 59220 7362
rect 59052 7252 59108 7262
rect 59052 7158 59108 7196
rect 58716 7084 58884 7140
rect 58716 7028 58772 7084
rect 58604 6972 58772 7028
rect 59164 7028 59220 7310
rect 59276 7364 59332 7374
rect 59276 7140 59332 7308
rect 59724 7140 59780 7534
rect 59276 7084 59444 7140
rect 59164 6972 59332 7028
rect 58604 6804 58660 6972
rect 58716 6804 58772 6814
rect 58380 6748 58548 6804
rect 58604 6802 58772 6804
rect 58604 6750 58718 6802
rect 58770 6750 58772 6802
rect 58604 6748 58772 6750
rect 58492 6580 58548 6748
rect 58716 6738 58772 6748
rect 59276 6804 59332 6972
rect 59276 6738 59332 6748
rect 58940 6692 58996 6702
rect 58940 6598 58996 6636
rect 58604 6580 58660 6590
rect 58492 6578 58660 6580
rect 58492 6526 58606 6578
rect 58658 6526 58660 6578
rect 58492 6524 58660 6526
rect 58604 6514 58660 6524
rect 58268 5954 58324 5964
rect 58380 6468 58436 6478
rect 59388 6468 59444 7084
rect 59724 7074 59780 7084
rect 59612 7028 59668 7038
rect 59612 6914 59668 6972
rect 59612 6862 59614 6914
rect 59666 6862 59668 6914
rect 59612 6850 59668 6862
rect 58380 5684 58436 6412
rect 59052 6412 59444 6468
rect 59500 6578 59556 6590
rect 59500 6526 59502 6578
rect 59554 6526 59556 6578
rect 58604 6132 58660 6142
rect 58380 5618 58436 5628
rect 58492 5908 58548 5918
rect 58156 5404 58436 5460
rect 58380 5010 58436 5404
rect 58380 4958 58382 5010
rect 58434 4958 58436 5010
rect 58380 4946 58436 4958
rect 58044 2482 58100 2492
rect 58492 800 58548 5852
rect 58604 4450 58660 6076
rect 58716 6018 58772 6030
rect 58716 5966 58718 6018
rect 58770 5966 58772 6018
rect 58716 5236 58772 5966
rect 58828 6020 58884 6030
rect 59052 6020 59108 6412
rect 59172 6300 59436 6310
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59172 6234 59436 6244
rect 59500 6132 59556 6526
rect 59724 6468 59780 6478
rect 59612 6466 59780 6468
rect 59612 6414 59726 6466
rect 59778 6414 59780 6466
rect 59612 6412 59780 6414
rect 59612 6356 59668 6412
rect 59724 6402 59780 6412
rect 59612 6290 59668 6300
rect 59724 6244 59780 6254
rect 59500 6076 59668 6132
rect 59052 5964 59220 6020
rect 58828 5908 58884 5964
rect 58940 5908 58996 5918
rect 58828 5906 58996 5908
rect 58828 5854 58942 5906
rect 58994 5854 58996 5906
rect 58828 5852 58996 5854
rect 58940 5842 58996 5852
rect 58716 5170 58772 5180
rect 58940 5684 58996 5694
rect 58604 4398 58606 4450
rect 58658 4398 58660 4450
rect 58604 4386 58660 4398
rect 58716 4900 58772 4910
rect 58716 3444 58772 4844
rect 58716 3378 58772 3388
rect 58940 3332 58996 5628
rect 59164 4900 59220 5964
rect 59500 5908 59556 5918
rect 59388 5682 59444 5694
rect 59388 5630 59390 5682
rect 59442 5630 59444 5682
rect 59388 5122 59444 5630
rect 59500 5684 59556 5852
rect 59500 5618 59556 5628
rect 59388 5070 59390 5122
rect 59442 5070 59444 5122
rect 59388 5058 59444 5070
rect 59500 5122 59556 5134
rect 59500 5070 59502 5122
rect 59554 5070 59556 5122
rect 59052 4844 59220 4900
rect 59388 4900 59444 4910
rect 59500 4900 59556 5070
rect 59444 4844 59556 4900
rect 59052 3780 59108 4844
rect 59388 4834 59444 4844
rect 59612 4788 59668 6076
rect 59724 5234 59780 6188
rect 59724 5182 59726 5234
rect 59778 5182 59780 5234
rect 59724 5170 59780 5182
rect 59172 4732 59436 4742
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59172 4666 59436 4676
rect 59500 4732 59668 4788
rect 59724 4898 59780 4910
rect 59724 4846 59726 4898
rect 59778 4846 59780 4898
rect 59388 4228 59444 4238
rect 59052 3714 59108 3724
rect 59164 4116 59220 4126
rect 59164 3778 59220 4060
rect 59164 3726 59166 3778
rect 59218 3726 59220 3778
rect 59164 3714 59220 3726
rect 59276 4114 59332 4126
rect 59276 4062 59278 4114
rect 59330 4062 59332 4114
rect 59276 3388 59332 4062
rect 59388 3778 59444 4172
rect 59388 3726 59390 3778
rect 59442 3726 59444 3778
rect 59388 3714 59444 3726
rect 58940 3266 58996 3276
rect 59052 3332 59332 3388
rect 59052 1204 59108 3332
rect 59500 3330 59556 4732
rect 59724 4676 59780 4846
rect 59500 3278 59502 3330
rect 59554 3278 59556 3330
rect 59500 3266 59556 3278
rect 59612 3554 59668 3566
rect 59612 3502 59614 3554
rect 59666 3502 59668 3554
rect 59172 3164 59436 3174
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59172 3098 59436 3108
rect 59612 2996 59668 3502
rect 59724 3556 59780 4620
rect 59724 3490 59780 3500
rect 59836 3388 59892 7868
rect 59948 7364 60004 8428
rect 59948 7298 60004 7308
rect 59948 7028 60004 7038
rect 59948 6692 60004 6972
rect 60060 6804 60116 8764
rect 60060 6738 60116 6748
rect 60172 7586 60228 7598
rect 60172 7534 60174 7586
rect 60226 7534 60228 7586
rect 59948 6626 60004 6636
rect 59948 6468 60004 6478
rect 59948 6466 60116 6468
rect 59948 6414 59950 6466
rect 60002 6414 60116 6466
rect 59948 6412 60116 6414
rect 59948 6402 60004 6412
rect 59948 5794 60004 5806
rect 59948 5742 59950 5794
rect 60002 5742 60004 5794
rect 59948 5460 60004 5742
rect 60060 5684 60116 6412
rect 60172 6020 60228 7534
rect 60172 5954 60228 5964
rect 60172 5796 60228 5806
rect 60284 5796 60340 9212
rect 60844 8930 60900 8942
rect 60844 8878 60846 8930
rect 60898 8878 60900 8930
rect 60508 8818 60564 8830
rect 60508 8766 60510 8818
rect 60562 8766 60564 8818
rect 60396 8708 60452 8718
rect 60396 6020 60452 8652
rect 60396 5954 60452 5964
rect 60172 5794 60340 5796
rect 60172 5742 60174 5794
rect 60226 5742 60340 5794
rect 60172 5740 60340 5742
rect 60396 5796 60452 5806
rect 60172 5730 60228 5740
rect 60396 5702 60452 5740
rect 60060 5618 60116 5628
rect 59948 5394 60004 5404
rect 60284 5460 60340 5470
rect 59948 5122 60004 5134
rect 59948 5070 59950 5122
rect 60002 5070 60004 5122
rect 59948 4788 60004 5070
rect 60284 4900 60340 5404
rect 59948 3554 60004 4732
rect 59948 3502 59950 3554
rect 60002 3502 60004 3554
rect 59948 3490 60004 3502
rect 60060 4844 60340 4900
rect 60396 5346 60452 5358
rect 60396 5294 60398 5346
rect 60450 5294 60452 5346
rect 59612 2930 59668 2940
rect 59724 3332 59892 3388
rect 59724 2772 59780 3332
rect 59052 1138 59108 1148
rect 59164 2716 59780 2772
rect 59836 3220 59892 3230
rect 59164 800 59220 2716
rect 59836 800 59892 3164
rect 60060 2884 60116 4844
rect 60172 3556 60228 3566
rect 60172 3462 60228 3500
rect 60396 3554 60452 5294
rect 60396 3502 60398 3554
rect 60450 3502 60452 3554
rect 60396 3490 60452 3502
rect 60284 3442 60340 3454
rect 60284 3390 60286 3442
rect 60338 3390 60340 3442
rect 60284 3388 60340 3390
rect 60284 3332 60452 3388
rect 60396 2996 60452 3332
rect 60396 2930 60452 2940
rect 60060 2818 60116 2828
rect 60508 800 60564 8766
rect 60732 8820 60788 8830
rect 60732 8148 60788 8764
rect 60732 8082 60788 8092
rect 60620 8034 60676 8046
rect 60620 7982 60622 8034
rect 60674 7982 60676 8034
rect 60620 5460 60676 7982
rect 60732 7924 60788 7934
rect 60732 7700 60788 7868
rect 60844 7812 60900 8878
rect 60956 7924 61012 9548
rect 61180 9266 61236 9772
rect 61180 9214 61182 9266
rect 61234 9214 61236 9266
rect 61180 8484 61236 9214
rect 61292 9716 61348 9726
rect 61292 9602 61348 9660
rect 61292 9550 61294 9602
rect 61346 9550 61348 9602
rect 61292 8708 61348 9550
rect 61964 9156 62020 9166
rect 61628 9154 62020 9156
rect 61628 9102 61966 9154
rect 62018 9102 62020 9154
rect 61628 9100 62020 9102
rect 61292 8642 61348 8652
rect 61404 9044 61460 9054
rect 61180 8418 61236 8428
rect 61068 8148 61124 8158
rect 61068 8146 61348 8148
rect 61068 8094 61070 8146
rect 61122 8094 61348 8146
rect 61068 8092 61348 8094
rect 61068 8082 61124 8092
rect 60956 7868 61124 7924
rect 60844 7746 60900 7756
rect 60732 6802 60788 7644
rect 60956 7588 61012 7598
rect 60732 6750 60734 6802
rect 60786 6750 60788 6802
rect 60732 6738 60788 6750
rect 60844 7586 61012 7588
rect 60844 7534 60958 7586
rect 61010 7534 61012 7586
rect 60844 7532 61012 7534
rect 60732 6580 60788 6590
rect 60732 5684 60788 6524
rect 60732 5618 60788 5628
rect 60620 5394 60676 5404
rect 60620 5236 60676 5246
rect 60620 5142 60676 5180
rect 60620 4004 60676 4014
rect 60620 3554 60676 3948
rect 60844 3668 60900 7532
rect 60956 7522 61012 7532
rect 60956 7252 61012 7262
rect 60956 6244 61012 7196
rect 60956 6178 61012 6188
rect 61068 7028 61124 7868
rect 61068 6466 61124 6972
rect 61068 6414 61070 6466
rect 61122 6414 61124 6466
rect 60620 3502 60622 3554
rect 60674 3502 60676 3554
rect 60620 3490 60676 3502
rect 60732 3612 60900 3668
rect 60956 5908 61012 5918
rect 60732 3220 60788 3612
rect 60956 3554 61012 5852
rect 61068 5346 61124 6414
rect 61068 5294 61070 5346
rect 61122 5294 61124 5346
rect 61068 5282 61124 5294
rect 61180 7812 61236 7822
rect 61068 5124 61124 5134
rect 61068 5030 61124 5068
rect 61068 4228 61124 4238
rect 61068 3666 61124 4172
rect 61180 4004 61236 7756
rect 61180 3938 61236 3948
rect 61068 3614 61070 3666
rect 61122 3614 61124 3666
rect 61068 3602 61124 3614
rect 61180 3780 61236 3790
rect 60956 3502 60958 3554
rect 61010 3502 61012 3554
rect 60956 3490 61012 3502
rect 61180 3554 61236 3724
rect 61180 3502 61182 3554
rect 61234 3502 61236 3554
rect 61180 3490 61236 3502
rect 61292 3388 61348 8092
rect 61404 5236 61460 8988
rect 61628 8818 61684 9100
rect 61964 9090 62020 9100
rect 61740 8932 61796 8942
rect 61740 8930 62020 8932
rect 61740 8878 61742 8930
rect 61794 8878 62020 8930
rect 61740 8876 62020 8878
rect 61740 8866 61796 8876
rect 61628 8766 61630 8818
rect 61682 8766 61684 8818
rect 61628 8754 61684 8766
rect 61740 8484 61796 8494
rect 61740 8258 61796 8428
rect 61740 8206 61742 8258
rect 61794 8206 61796 8258
rect 61516 8034 61572 8046
rect 61516 7982 61518 8034
rect 61570 7982 61572 8034
rect 61516 7588 61572 7982
rect 61516 7522 61572 7532
rect 61740 7476 61796 8206
rect 61740 7410 61796 7420
rect 61852 8260 61908 8270
rect 61516 7364 61572 7374
rect 61516 7270 61572 7308
rect 61740 7028 61796 7038
rect 61516 6916 61572 6926
rect 61516 6802 61572 6860
rect 61516 6750 61518 6802
rect 61570 6750 61572 6802
rect 61516 6738 61572 6750
rect 61740 6468 61796 6972
rect 61852 6580 61908 8204
rect 61852 6514 61908 6524
rect 61740 6402 61796 6412
rect 61964 6356 62020 8876
rect 61964 6290 62020 6300
rect 62076 6132 62132 10780
rect 63532 10500 63588 10510
rect 63532 10498 63700 10500
rect 63532 10446 63534 10498
rect 63586 10446 63700 10498
rect 63532 10444 63700 10446
rect 63532 10434 63588 10444
rect 62748 10388 62804 10398
rect 62524 9604 62580 9614
rect 62412 9602 62580 9604
rect 62412 9550 62526 9602
rect 62578 9550 62580 9602
rect 62412 9548 62580 9550
rect 62300 8932 62356 8942
rect 62300 8484 62356 8876
rect 62300 8418 62356 8428
rect 62188 8370 62244 8382
rect 62188 8318 62190 8370
rect 62242 8318 62244 8370
rect 62188 8260 62244 8318
rect 62188 8194 62244 8204
rect 62188 8036 62244 8046
rect 62188 7700 62244 7980
rect 62188 7364 62244 7644
rect 62188 7298 62244 7308
rect 62300 8034 62356 8046
rect 62300 7982 62302 8034
rect 62354 7982 62356 8034
rect 62076 6066 62132 6076
rect 62188 7140 62244 7150
rect 61740 6018 61796 6030
rect 61740 5966 61742 6018
rect 61794 5966 61796 6018
rect 61740 5908 61796 5966
rect 62188 5908 62244 7084
rect 62300 6804 62356 7982
rect 62300 6738 62356 6748
rect 62412 6580 62468 9548
rect 62524 9538 62580 9548
rect 62524 9044 62580 9054
rect 62524 8950 62580 8988
rect 62636 8484 62692 8494
rect 62524 8260 62580 8270
rect 62524 8166 62580 8204
rect 62412 6514 62468 6524
rect 62524 7588 62580 7598
rect 62524 6468 62580 7532
rect 62524 6356 62580 6412
rect 61740 5852 62244 5908
rect 62300 6300 62580 6356
rect 61740 5684 61796 5694
rect 61628 5628 61740 5684
rect 61404 5170 61460 5180
rect 61516 5572 61572 5582
rect 61516 5234 61572 5516
rect 61516 5182 61518 5234
rect 61570 5182 61572 5234
rect 61516 5170 61572 5182
rect 61628 4564 61684 5628
rect 61740 5618 61796 5628
rect 62076 5460 62132 5470
rect 62132 5404 62244 5460
rect 62076 5394 62132 5404
rect 61404 4508 61684 4564
rect 61404 3554 61460 4508
rect 61404 3502 61406 3554
rect 61458 3502 61460 3554
rect 61404 3490 61460 3502
rect 61740 4450 61796 4462
rect 61740 4398 61742 4450
rect 61794 4398 61796 4450
rect 60732 3154 60788 3164
rect 60956 3332 61012 3342
rect 60956 800 61012 3276
rect 61180 3332 61348 3388
rect 61180 800 61236 3332
rect 61740 2996 61796 4398
rect 62076 4004 62132 4014
rect 61740 2930 61796 2940
rect 61852 3332 61908 3342
rect 61404 2882 61460 2894
rect 61404 2830 61406 2882
rect 61458 2830 61460 2882
rect 61404 800 61460 2830
rect 61628 1874 61684 1886
rect 61628 1822 61630 1874
rect 61682 1822 61684 1874
rect 61628 800 61684 1822
rect 61852 800 61908 3276
rect 61964 3330 62020 3342
rect 61964 3278 61966 3330
rect 62018 3278 62020 3330
rect 61964 1764 62020 3278
rect 61964 1698 62020 1708
rect 62076 800 62132 3948
rect 62188 3332 62244 5404
rect 62300 4788 62356 6300
rect 62524 6132 62580 6142
rect 62300 4722 62356 4732
rect 62412 5794 62468 5806
rect 62412 5742 62414 5794
rect 62466 5742 62468 5794
rect 62412 4452 62468 5742
rect 62412 4386 62468 4396
rect 62524 4450 62580 6076
rect 62636 5348 62692 8428
rect 62748 7140 62804 10332
rect 63532 10164 63588 10174
rect 63084 9828 63140 9838
rect 62860 9154 62916 9166
rect 62860 9102 62862 9154
rect 62914 9102 62916 9154
rect 62860 8932 62916 9102
rect 62860 8866 62916 8876
rect 63084 8708 63140 9772
rect 63420 9604 63476 9614
rect 63308 9602 63476 9604
rect 63308 9550 63422 9602
rect 63474 9550 63476 9602
rect 63308 9548 63476 9550
rect 63196 9042 63252 9054
rect 63196 8990 63198 9042
rect 63250 8990 63252 9042
rect 63196 8820 63252 8990
rect 63196 8754 63252 8764
rect 62860 8652 63140 8708
rect 62860 7812 62916 8652
rect 63308 8484 63364 9548
rect 63420 9538 63476 9548
rect 63532 9266 63588 10108
rect 63532 9214 63534 9266
rect 63586 9214 63588 9266
rect 63532 9202 63588 9214
rect 63644 9044 63700 10444
rect 63980 10498 64036 10510
rect 63980 10446 63982 10498
rect 64034 10446 64036 10498
rect 63196 8428 63364 8484
rect 63532 8988 63700 9044
rect 63868 9042 63924 9054
rect 63868 8990 63870 9042
rect 63922 8990 63924 9042
rect 63532 8484 63588 8988
rect 62860 7756 63028 7812
rect 62860 7588 62916 7598
rect 62860 7494 62916 7532
rect 62972 7364 63028 7756
rect 62748 7074 62804 7084
rect 62860 7308 63028 7364
rect 62860 6578 62916 7308
rect 63084 6692 63140 6702
rect 62860 6526 62862 6578
rect 62914 6526 62916 6578
rect 62860 6514 62916 6526
rect 62972 6580 63028 6590
rect 62636 5282 62692 5292
rect 62748 6356 62804 6366
rect 62748 6018 62804 6300
rect 62748 5966 62750 6018
rect 62802 5966 62804 6018
rect 62524 4398 62526 4450
rect 62578 4398 62580 4450
rect 62412 4116 62468 4126
rect 62188 3266 62244 3276
rect 62300 3668 62356 3678
rect 62300 800 62356 3612
rect 62412 2996 62468 4060
rect 62524 3444 62580 4398
rect 62524 3378 62580 3388
rect 62636 5010 62692 5022
rect 62636 4958 62638 5010
rect 62690 4958 62692 5010
rect 62636 3220 62692 4958
rect 62748 3780 62804 5966
rect 62860 6020 62916 6030
rect 62860 5794 62916 5964
rect 62860 5742 62862 5794
rect 62914 5742 62916 5794
rect 62860 4228 62916 5742
rect 62860 4162 62916 4172
rect 62748 3714 62804 3724
rect 62860 4004 62916 4014
rect 62860 3442 62916 3948
rect 62860 3390 62862 3442
rect 62914 3390 62916 3442
rect 62860 3378 62916 3390
rect 62636 3154 62692 3164
rect 62412 2940 62580 2996
rect 62524 800 62580 2940
rect 62748 2770 62804 2782
rect 62748 2718 62750 2770
rect 62802 2718 62804 2770
rect 62748 800 62804 2718
rect 62972 800 63028 6524
rect 63084 5908 63140 6636
rect 63084 5814 63140 5852
rect 63196 5124 63252 8428
rect 63532 8418 63588 8428
rect 63868 8484 63924 8990
rect 63868 8418 63924 8428
rect 63644 8372 63700 8382
rect 63532 8260 63588 8270
rect 63532 8166 63588 8204
rect 63644 8258 63700 8316
rect 63644 8206 63646 8258
rect 63698 8206 63700 8258
rect 63644 8194 63700 8206
rect 63868 8260 63924 8270
rect 63868 8166 63924 8204
rect 63308 8034 63364 8046
rect 63308 7982 63310 8034
rect 63362 7982 63364 8034
rect 63308 6690 63364 7982
rect 63420 8036 63476 8046
rect 63420 8034 63924 8036
rect 63420 7982 63422 8034
rect 63474 7982 63924 8034
rect 63420 7980 63924 7982
rect 63420 7970 63476 7980
rect 63868 7812 63924 7980
rect 63980 7924 64036 10446
rect 64540 10498 64596 10510
rect 64540 10446 64542 10498
rect 64594 10446 64596 10498
rect 64204 9604 64260 9614
rect 64092 9602 64260 9604
rect 64092 9550 64206 9602
rect 64258 9550 64260 9602
rect 64092 9548 64260 9550
rect 64092 8148 64148 9548
rect 64204 9538 64260 9548
rect 64428 9492 64484 9502
rect 64316 9436 64428 9492
rect 64092 8082 64148 8092
rect 64204 9380 64260 9390
rect 63980 7858 64036 7868
rect 63868 7476 63924 7756
rect 64204 7588 64260 9324
rect 64204 7522 64260 7532
rect 63644 7420 63924 7476
rect 63532 7364 63588 7402
rect 63532 7298 63588 7308
rect 63420 7252 63476 7290
rect 63420 7186 63476 7196
rect 63644 7140 63700 7420
rect 63532 7084 63700 7140
rect 63756 7250 63812 7262
rect 63756 7198 63758 7250
rect 63810 7198 63812 7250
rect 63420 6804 63476 6814
rect 63420 6710 63476 6748
rect 63308 6638 63310 6690
rect 63362 6638 63364 6690
rect 63308 6468 63364 6638
rect 63308 6402 63364 6412
rect 63532 6466 63588 7084
rect 63756 6916 63812 7198
rect 63868 7250 63924 7262
rect 63868 7198 63870 7250
rect 63922 7198 63924 7250
rect 63868 7028 63924 7198
rect 63868 6962 63924 6972
rect 63532 6414 63534 6466
rect 63586 6414 63588 6466
rect 63196 5068 63364 5124
rect 63196 4900 63252 4910
rect 63084 4898 63252 4900
rect 63084 4846 63198 4898
rect 63250 4846 63252 4898
rect 63084 4844 63252 4846
rect 63084 1540 63140 4844
rect 63196 4834 63252 4844
rect 63308 4676 63364 5068
rect 63084 1474 63140 1484
rect 63196 4620 63364 4676
rect 63532 4676 63588 6414
rect 63644 6804 63700 6814
rect 63644 6356 63700 6748
rect 63756 6692 63812 6860
rect 64204 6916 64260 6926
rect 63756 6636 63924 6692
rect 63644 6290 63700 6300
rect 63756 6468 63812 6478
rect 63756 6132 63812 6412
rect 63868 6356 63924 6636
rect 63868 6290 63924 6300
rect 63980 6578 64036 6590
rect 63980 6526 63982 6578
rect 64034 6526 64036 6578
rect 63196 800 63252 4620
rect 63532 4610 63588 4620
rect 63644 6076 63812 6132
rect 63644 4564 63700 6076
rect 63756 5908 63812 5918
rect 63756 5814 63812 5852
rect 63980 5348 64036 6526
rect 64204 6244 64260 6860
rect 64316 6468 64372 9436
rect 64428 9426 64484 9436
rect 64428 8258 64484 8270
rect 64428 8206 64430 8258
rect 64482 8206 64484 8258
rect 64428 7364 64484 8206
rect 64540 7476 64596 10446
rect 65100 10498 65156 10510
rect 65100 10446 65102 10498
rect 65154 10446 65156 10498
rect 64764 9602 64820 9614
rect 64764 9550 64766 9602
rect 64818 9550 64820 9602
rect 64652 9268 64708 9278
rect 64652 9174 64708 9212
rect 64540 7382 64596 7420
rect 64652 8484 64708 8494
rect 64428 6804 64484 7308
rect 64428 6738 64484 6748
rect 64540 6580 64596 6590
rect 64540 6486 64596 6524
rect 64316 6402 64372 6412
rect 64652 6244 64708 8428
rect 64204 6188 64372 6244
rect 63980 5282 64036 5292
rect 64204 5460 64260 5470
rect 64092 5236 64148 5246
rect 63644 4498 63700 4508
rect 63756 4788 63812 4798
rect 63420 4452 63476 4462
rect 63420 800 63476 4396
rect 63756 3388 63812 4732
rect 63980 4676 64036 4686
rect 63868 4228 63924 4238
rect 63868 4134 63924 4172
rect 63644 3332 63812 3388
rect 63644 800 63700 3332
rect 63980 2996 64036 4620
rect 63868 2940 64036 2996
rect 63868 800 63924 2940
rect 64092 800 64148 5180
rect 64204 2772 64260 5404
rect 64204 2706 64260 2716
rect 64316 800 64372 6188
rect 64652 6178 64708 6188
rect 64540 6018 64596 6030
rect 64540 5966 64542 6018
rect 64594 5966 64596 6018
rect 64540 4676 64596 5966
rect 64540 4610 64596 4620
rect 64652 6020 64708 6030
rect 64428 4564 64484 4574
rect 64428 1874 64484 4508
rect 64540 4452 64596 4462
rect 64540 4358 64596 4396
rect 64652 4116 64708 5964
rect 64764 5236 64820 9550
rect 64876 9042 64932 9054
rect 64876 8990 64878 9042
rect 64930 8990 64932 9042
rect 64876 8484 64932 8990
rect 64876 8418 64932 8428
rect 64988 9044 65044 9054
rect 64988 8260 65044 8988
rect 64988 8166 65044 8204
rect 64988 7476 65044 7486
rect 64876 7362 64932 7374
rect 64876 7310 64878 7362
rect 64930 7310 64932 7362
rect 64876 7140 64932 7310
rect 64876 6692 64932 7084
rect 64876 6626 64932 6636
rect 64764 5170 64820 5180
rect 64652 4050 64708 4060
rect 64428 1822 64430 1874
rect 64482 1822 64484 1874
rect 64428 1810 64484 1822
rect 64540 3780 64596 3790
rect 64540 800 64596 3724
rect 64876 3556 64932 3566
rect 64876 3388 64932 3500
rect 64764 3332 64932 3388
rect 64764 800 64820 3332
rect 64988 800 65044 7420
rect 65100 6356 65156 10446
rect 65436 10498 65492 10510
rect 65436 10446 65438 10498
rect 65490 10446 65492 10498
rect 65212 9940 65268 9950
rect 65212 9268 65268 9884
rect 65324 9602 65380 9614
rect 65324 9550 65326 9602
rect 65378 9550 65380 9602
rect 65324 9492 65380 9550
rect 65324 9426 65380 9436
rect 65324 9268 65380 9278
rect 65212 9266 65380 9268
rect 65212 9214 65326 9266
rect 65378 9214 65380 9266
rect 65212 9212 65380 9214
rect 65324 9202 65380 9212
rect 65212 8820 65268 8830
rect 65212 7812 65268 8764
rect 65324 8484 65380 8494
rect 65324 8260 65380 8428
rect 65436 8372 65492 10446
rect 65548 10500 65604 10510
rect 65548 9044 65604 10444
rect 66220 10498 66276 10510
rect 66220 10446 66222 10498
rect 66274 10446 66276 10498
rect 66220 9828 66276 10446
rect 66556 10052 66612 11788
rect 67116 11508 67172 17388
rect 78492 17276 78756 17286
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78492 17210 78756 17220
rect 68832 16492 69096 16502
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 68832 16426 69096 16436
rect 78492 15708 78756 15718
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78492 15642 78756 15652
rect 69804 15204 69860 15214
rect 68832 14924 69096 14934
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 68832 14858 69096 14868
rect 68832 13356 69096 13366
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 68832 13290 69096 13300
rect 67116 11442 67172 11452
rect 67452 11956 67508 11966
rect 67004 10500 67060 10510
rect 67004 10498 67172 10500
rect 67004 10446 67006 10498
rect 67058 10446 67172 10498
rect 67004 10444 67172 10446
rect 67004 10434 67060 10444
rect 66556 9986 66612 9996
rect 66668 10276 66724 10286
rect 65772 9772 66276 9828
rect 65660 9714 65716 9726
rect 65660 9662 65662 9714
rect 65714 9662 65716 9714
rect 65660 9268 65716 9662
rect 65660 9202 65716 9212
rect 65548 8978 65604 8988
rect 65660 9042 65716 9054
rect 65660 8990 65662 9042
rect 65714 8990 65716 9042
rect 65660 8820 65716 8990
rect 65660 8754 65716 8764
rect 65436 8316 65604 8372
rect 65548 8260 65604 8316
rect 65324 8204 65492 8260
rect 65324 8036 65380 8046
rect 65436 8036 65492 8204
rect 65548 8166 65604 8204
rect 65436 7980 65716 8036
rect 65324 7942 65380 7980
rect 65548 7812 65604 7822
rect 65212 7756 65492 7812
rect 65324 7588 65380 7598
rect 65100 6290 65156 6300
rect 65212 7586 65380 7588
rect 65212 7534 65326 7586
rect 65378 7534 65380 7586
rect 65212 7532 65380 7534
rect 65100 6018 65156 6030
rect 65100 5966 65102 6018
rect 65154 5966 65156 6018
rect 65100 5236 65156 5966
rect 65100 5170 65156 5180
rect 65212 3780 65268 7532
rect 65324 7522 65380 7532
rect 65436 7028 65492 7756
rect 65212 3714 65268 3724
rect 65324 6972 65492 7028
rect 65324 3778 65380 6972
rect 65324 3726 65326 3778
rect 65378 3726 65380 3778
rect 65324 3714 65380 3726
rect 65436 6804 65492 6814
rect 65436 3556 65492 6748
rect 65548 4564 65604 7756
rect 65660 6802 65716 7980
rect 65660 6750 65662 6802
rect 65714 6750 65716 6802
rect 65660 6738 65716 6750
rect 65660 6468 65716 6478
rect 65660 5236 65716 6412
rect 65772 6356 65828 9772
rect 66220 9602 66276 9614
rect 66220 9550 66222 9602
rect 66274 9550 66276 9602
rect 66108 9268 66164 9278
rect 66220 9268 66276 9550
rect 66668 9268 66724 10220
rect 66780 9716 66836 9726
rect 66780 9622 66836 9660
rect 67004 9604 67060 9614
rect 66892 9602 67060 9604
rect 66892 9550 67006 9602
rect 67058 9550 67060 9602
rect 66892 9548 67060 9550
rect 66780 9268 66836 9278
rect 66220 9212 66500 9268
rect 66668 9266 66836 9268
rect 66668 9214 66782 9266
rect 66834 9214 66836 9266
rect 66668 9212 66836 9214
rect 65996 9154 66052 9166
rect 65996 9102 65998 9154
rect 66050 9102 66052 9154
rect 65996 9044 66052 9102
rect 65996 8978 66052 8988
rect 65996 8372 66052 8382
rect 65884 8260 65940 8270
rect 65884 7812 65940 8204
rect 65996 8146 66052 8316
rect 65996 8094 65998 8146
rect 66050 8094 66052 8146
rect 65996 8082 66052 8094
rect 65884 7746 65940 7756
rect 65884 7586 65940 7598
rect 65884 7534 65886 7586
rect 65938 7534 65940 7586
rect 65884 7364 65940 7534
rect 65884 7298 65940 7308
rect 65996 7588 66052 7598
rect 65996 6468 66052 7532
rect 66108 6580 66164 9212
rect 66220 9042 66276 9054
rect 66220 8990 66222 9042
rect 66274 8990 66276 9042
rect 66220 7252 66276 8990
rect 66332 8372 66388 8382
rect 66444 8372 66500 9212
rect 66780 9202 66836 9212
rect 66388 8316 66500 8372
rect 66668 8596 66724 8606
rect 66892 8596 66948 9548
rect 67004 9538 67060 9548
rect 67116 9268 67172 10444
rect 66332 8306 66388 8316
rect 66556 8260 66612 8270
rect 66332 8148 66388 8158
rect 66332 8146 66500 8148
rect 66332 8094 66334 8146
rect 66386 8094 66500 8146
rect 66332 8092 66500 8094
rect 66332 8082 66388 8092
rect 66220 7186 66276 7196
rect 66332 7474 66388 7486
rect 66332 7422 66334 7474
rect 66386 7422 66388 7474
rect 66332 7140 66388 7422
rect 66332 7074 66388 7084
rect 66108 6524 66388 6580
rect 65996 6412 66276 6468
rect 65772 6300 66052 6356
rect 65660 5180 65828 5236
rect 65548 4498 65604 4508
rect 65660 5010 65716 5022
rect 65660 4958 65662 5010
rect 65714 4958 65716 5010
rect 65324 3500 65492 3556
rect 65548 3892 65604 3902
rect 65324 3332 65380 3500
rect 65548 3442 65604 3836
rect 65548 3390 65550 3442
rect 65602 3390 65604 3442
rect 65548 3378 65604 3390
rect 65212 3276 65380 3332
rect 65436 3332 65492 3342
rect 65212 800 65268 3276
rect 65436 800 65492 3276
rect 65660 3332 65716 4958
rect 65772 4452 65828 5180
rect 65772 4386 65828 4396
rect 65884 5012 65940 5022
rect 65772 4228 65828 4238
rect 65772 3554 65828 4172
rect 65772 3502 65774 3554
rect 65826 3502 65828 3554
rect 65772 3490 65828 3502
rect 65660 3266 65716 3276
rect 65660 2548 65716 2558
rect 65660 800 65716 2492
rect 65884 800 65940 4956
rect 65996 2770 66052 6300
rect 66108 6244 66164 6254
rect 66108 5234 66164 6188
rect 66108 5182 66110 5234
rect 66162 5182 66164 5234
rect 66108 5170 66164 5182
rect 66220 3556 66276 6412
rect 66332 3778 66388 6524
rect 66444 5012 66500 8092
rect 66556 7588 66612 8204
rect 66668 8146 66724 8540
rect 66668 8094 66670 8146
rect 66722 8094 66724 8146
rect 66668 8082 66724 8094
rect 66780 8540 66948 8596
rect 67004 9212 67172 9268
rect 67228 9716 67284 9726
rect 66668 7700 66724 7710
rect 66668 7606 66724 7644
rect 66556 7522 66612 7532
rect 66668 7364 66724 7374
rect 66556 7028 66612 7038
rect 66556 6690 66612 6972
rect 66556 6638 66558 6690
rect 66610 6638 66612 6690
rect 66556 6626 66612 6638
rect 66668 6578 66724 7308
rect 66668 6526 66670 6578
rect 66722 6526 66724 6578
rect 66668 6514 66724 6526
rect 66780 6468 66836 8540
rect 66892 8372 66948 8382
rect 66892 8258 66948 8316
rect 66892 8206 66894 8258
rect 66946 8206 66948 8258
rect 66892 8194 66948 8206
rect 66892 7812 66948 7822
rect 66892 7474 66948 7756
rect 66892 7422 66894 7474
rect 66946 7422 66948 7474
rect 66892 7410 66948 7422
rect 66780 6402 66836 6412
rect 66892 7140 66948 7150
rect 66892 5908 66948 7084
rect 66668 5852 66948 5908
rect 66444 4956 66612 5012
rect 66556 4564 66612 4956
rect 66668 4788 66724 5852
rect 66668 4722 66724 4732
rect 66780 5124 66836 5134
rect 66556 4508 66724 4564
rect 66444 4452 66500 4462
rect 66500 4396 66612 4452
rect 66444 4386 66500 4396
rect 66332 3726 66334 3778
rect 66386 3726 66388 3778
rect 66332 3714 66388 3726
rect 66220 3500 66388 3556
rect 65996 2718 65998 2770
rect 66050 2718 66052 2770
rect 65996 2706 66052 2718
rect 66108 2658 66164 2670
rect 66108 2606 66110 2658
rect 66162 2606 66164 2658
rect 66108 800 66164 2606
rect 66332 800 66388 3500
rect 66556 800 66612 4396
rect 66668 4226 66724 4508
rect 66668 4174 66670 4226
rect 66722 4174 66724 4226
rect 66668 4162 66724 4174
rect 66780 800 66836 5068
rect 67004 4788 67060 9212
rect 67116 9042 67172 9054
rect 67116 8990 67118 9042
rect 67170 8990 67172 9042
rect 67116 7364 67172 8990
rect 67228 8260 67284 9660
rect 67452 9714 67508 11900
rect 68832 11788 69096 11798
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 68832 11722 69096 11732
rect 69020 11618 69076 11630
rect 69020 11566 69022 11618
rect 69074 11566 69076 11618
rect 68908 11508 68964 11518
rect 69020 11508 69076 11566
rect 68964 11452 69076 11508
rect 68908 11442 68964 11452
rect 69020 11394 69076 11452
rect 69020 11342 69022 11394
rect 69074 11342 69076 11394
rect 69020 11330 69076 11342
rect 68572 11170 68628 11182
rect 68572 11118 68574 11170
rect 68626 11118 68628 11170
rect 68572 10724 68628 11118
rect 69468 11172 69524 11182
rect 69468 11170 69636 11172
rect 69468 11118 69470 11170
rect 69522 11118 69636 11170
rect 69468 11116 69636 11118
rect 69468 11106 69524 11116
rect 68012 10668 68628 10724
rect 69356 10724 69412 10734
rect 67452 9662 67454 9714
rect 67506 9662 67508 9714
rect 67452 9650 67508 9662
rect 67676 10498 67732 10510
rect 67676 10446 67678 10498
rect 67730 10446 67732 10498
rect 67228 8194 67284 8204
rect 67452 9154 67508 9166
rect 67452 9102 67454 9154
rect 67506 9102 67508 9154
rect 67340 8036 67396 8046
rect 67116 7298 67172 7308
rect 67228 8034 67396 8036
rect 67228 7982 67342 8034
rect 67394 7982 67396 8034
rect 67228 7980 67396 7982
rect 66892 4732 67060 4788
rect 67116 6580 67172 6590
rect 66892 4228 66948 4732
rect 67116 4676 67172 6524
rect 67228 5460 67284 7980
rect 67340 7970 67396 7980
rect 67340 7588 67396 7598
rect 67340 7494 67396 7532
rect 67340 7252 67396 7262
rect 67340 5794 67396 7196
rect 67452 6692 67508 9102
rect 67452 6626 67508 6636
rect 67564 8258 67620 8270
rect 67564 8206 67566 8258
rect 67618 8206 67620 8258
rect 67452 6466 67508 6478
rect 67452 6414 67454 6466
rect 67506 6414 67508 6466
rect 67452 6356 67508 6414
rect 67452 6290 67508 6300
rect 67340 5742 67342 5794
rect 67394 5742 67396 5794
rect 67340 5730 67396 5742
rect 67228 5394 67284 5404
rect 66892 3556 66948 4172
rect 66892 3490 66948 3500
rect 67004 4620 67172 4676
rect 67228 5010 67284 5022
rect 67228 4958 67230 5010
rect 67282 4958 67284 5010
rect 67004 800 67060 4620
rect 67228 4564 67284 4958
rect 67228 4498 67284 4508
rect 67340 4676 67396 4686
rect 67228 4116 67284 4126
rect 67228 800 67284 4060
rect 67340 2882 67396 4620
rect 67452 4564 67508 4574
rect 67452 3444 67508 4508
rect 67564 4452 67620 8206
rect 67676 7252 67732 10446
rect 67788 9714 67844 9726
rect 67788 9662 67790 9714
rect 67842 9662 67844 9714
rect 67788 8036 67844 9662
rect 67900 9156 67956 9166
rect 67900 9062 67956 9100
rect 67788 7970 67844 7980
rect 67900 8596 67956 8606
rect 67900 7588 67956 8540
rect 68012 7924 68068 10668
rect 68124 10498 68180 10510
rect 68124 10446 68126 10498
rect 68178 10446 68180 10498
rect 68124 8148 68180 10446
rect 68348 10500 68404 10510
rect 68236 9042 68292 9054
rect 68236 8990 68238 9042
rect 68290 8990 68292 9042
rect 68236 8260 68292 8990
rect 68348 8596 68404 10444
rect 68796 10498 68852 10510
rect 68796 10446 68798 10498
rect 68850 10446 68852 10498
rect 68796 10388 68852 10446
rect 69132 10500 69188 10510
rect 69132 10406 69188 10444
rect 68348 8530 68404 8540
rect 68460 10332 68852 10388
rect 68348 8372 68404 8382
rect 68348 8278 68404 8316
rect 68236 8194 68292 8204
rect 68124 8082 68180 8092
rect 68348 8036 68404 8046
rect 68012 7868 68180 7924
rect 67900 7522 67956 7532
rect 67676 7196 68068 7252
rect 67900 7028 67956 7038
rect 67676 6972 67900 7028
rect 67676 6690 67732 6972
rect 67900 6962 67956 6972
rect 67676 6638 67678 6690
rect 67730 6638 67732 6690
rect 67676 6626 67732 6638
rect 67788 6692 67844 6702
rect 67844 6636 67956 6692
rect 67788 6626 67844 6636
rect 67788 6020 67844 6030
rect 67788 5926 67844 5964
rect 67900 5124 67956 6636
rect 67788 5068 67956 5124
rect 68012 6020 68068 7196
rect 67788 5012 67844 5068
rect 67788 4946 67844 4956
rect 67900 4900 67956 4910
rect 67788 4788 67844 4798
rect 67564 4386 67620 4396
rect 67676 4450 67732 4462
rect 67676 4398 67678 4450
rect 67730 4398 67732 4450
rect 67676 4228 67732 4398
rect 67676 4162 67732 4172
rect 67452 3378 67508 3388
rect 67788 3108 67844 4732
rect 67676 3052 67844 3108
rect 67340 2830 67342 2882
rect 67394 2830 67396 2882
rect 67340 2818 67396 2830
rect 67452 2994 67508 3006
rect 67452 2942 67454 2994
rect 67506 2942 67508 2994
rect 67452 800 67508 2942
rect 67676 800 67732 3052
rect 67900 800 67956 4844
rect 68012 2994 68068 5964
rect 68124 5012 68180 7868
rect 68236 7588 68292 7598
rect 68236 7364 68292 7532
rect 68348 7476 68404 7980
rect 68460 7700 68516 10332
rect 68832 10220 69096 10230
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 68832 10154 69096 10164
rect 69244 10052 69300 10062
rect 68572 9604 68628 9614
rect 68572 9602 68740 9604
rect 68572 9550 68574 9602
rect 68626 9550 68740 9602
rect 68572 9548 68740 9550
rect 68572 9538 68628 9548
rect 68460 7634 68516 7644
rect 68572 9154 68628 9166
rect 68572 9102 68574 9154
rect 68626 9102 68628 9154
rect 68348 7420 68516 7476
rect 68236 7308 68404 7364
rect 68348 6580 68404 7308
rect 68460 7362 68516 7420
rect 68460 7310 68462 7362
rect 68514 7310 68516 7362
rect 68460 7298 68516 7310
rect 68572 7028 68628 9102
rect 68572 6962 68628 6972
rect 68572 6580 68628 6590
rect 68348 6524 68572 6580
rect 68572 6486 68628 6524
rect 68124 4676 68180 4956
rect 68124 4610 68180 4620
rect 68236 6468 68292 6478
rect 68012 2942 68014 2994
rect 68066 2942 68068 2994
rect 68012 2930 68068 2942
rect 68124 4340 68180 4350
rect 68124 800 68180 4284
rect 68236 3108 68292 6412
rect 68572 6244 68628 6254
rect 68460 6188 68572 6244
rect 68348 6020 68404 6030
rect 68348 5926 68404 5964
rect 68460 5236 68516 6188
rect 68572 6178 68628 6188
rect 68348 5180 68516 5236
rect 68348 4788 68404 5180
rect 68460 5012 68516 5022
rect 68460 4918 68516 4956
rect 68348 4722 68404 4732
rect 68684 4676 68740 9548
rect 69020 9602 69076 9614
rect 69020 9550 69022 9602
rect 69074 9550 69076 9602
rect 68796 9156 68852 9166
rect 68796 9042 68852 9100
rect 68796 8990 68798 9042
rect 68850 8990 68852 9042
rect 68796 8978 68852 8990
rect 69020 8820 69076 9550
rect 69244 9266 69300 9996
rect 69244 9214 69246 9266
rect 69298 9214 69300 9266
rect 69244 9202 69300 9214
rect 69020 8764 69300 8820
rect 68832 8652 69096 8662
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 68832 8586 69096 8596
rect 69244 8484 69300 8764
rect 69132 8428 69300 8484
rect 68908 8148 68964 8158
rect 68908 7252 68964 8092
rect 69020 7364 69076 7374
rect 69020 7270 69076 7308
rect 69132 7252 69188 8428
rect 69356 8372 69412 10668
rect 69244 8316 69412 8372
rect 69468 9602 69524 9614
rect 69468 9550 69470 9602
rect 69522 9550 69524 9602
rect 69244 7364 69300 8316
rect 69356 8148 69412 8158
rect 69356 8054 69412 8092
rect 69244 7308 69412 7364
rect 69132 7196 69300 7252
rect 68908 7186 68964 7196
rect 68832 7084 69096 7094
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 68832 7018 69096 7028
rect 68832 5516 69096 5526
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 68832 5450 69096 5460
rect 69020 5012 69076 5022
rect 68460 4620 68740 4676
rect 68908 4956 69020 5012
rect 68460 4116 68516 4620
rect 68908 4564 68964 4956
rect 69020 4946 69076 4956
rect 69244 4900 69300 7196
rect 69244 4834 69300 4844
rect 68460 4050 68516 4060
rect 68572 4508 68964 4564
rect 68460 3442 68516 3454
rect 68460 3390 68462 3442
rect 68514 3390 68516 3442
rect 68236 3052 68404 3108
rect 68348 800 68404 3052
rect 68460 2770 68516 3390
rect 68460 2718 68462 2770
rect 68514 2718 68516 2770
rect 68460 2706 68516 2718
rect 68572 800 68628 4508
rect 68796 4116 68852 4126
rect 68684 4060 68796 4116
rect 68684 3388 68740 4060
rect 68796 4050 68852 4060
rect 68832 3948 69096 3958
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 68832 3882 69096 3892
rect 69020 3556 69076 3566
rect 68684 3332 68852 3388
rect 68796 800 68852 3332
rect 69020 800 69076 3500
rect 69244 3332 69300 3342
rect 69132 3330 69300 3332
rect 69132 3278 69246 3330
rect 69298 3278 69300 3330
rect 69132 3276 69300 3278
rect 69132 3108 69188 3276
rect 69244 3266 69300 3276
rect 69356 3108 69412 7308
rect 69468 5012 69524 9550
rect 69580 9268 69636 11116
rect 69804 10498 69860 15148
rect 78492 14140 78756 14150
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78492 14074 78756 14084
rect 78492 12572 78756 12582
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78492 12506 78756 12516
rect 70476 11618 70532 11630
rect 70476 11566 70478 11618
rect 70530 11566 70532 11618
rect 69804 10446 69806 10498
rect 69858 10446 69860 10498
rect 69804 9828 69860 10446
rect 69804 9762 69860 9772
rect 69916 11170 69972 11182
rect 69916 11118 69918 11170
rect 69970 11118 69972 11170
rect 69916 9268 69972 11118
rect 70364 11170 70420 11182
rect 70364 11118 70366 11170
rect 70418 11118 70420 11170
rect 70252 10724 70308 10734
rect 70252 10630 70308 10668
rect 70140 10612 70196 10622
rect 70140 10050 70196 10556
rect 70140 9998 70142 10050
rect 70194 9998 70196 10050
rect 70140 9986 70196 9998
rect 69580 9212 69748 9268
rect 69580 9044 69636 9054
rect 69580 8950 69636 8988
rect 69580 8596 69636 8606
rect 69580 6132 69636 8540
rect 69692 6580 69748 9212
rect 69804 9212 69972 9268
rect 69804 9154 69860 9212
rect 69804 9102 69806 9154
rect 69858 9102 69860 9154
rect 69804 9090 69860 9102
rect 69804 8818 69860 8830
rect 69804 8766 69806 8818
rect 69858 8766 69860 8818
rect 69804 8708 69860 8766
rect 70140 8818 70196 8830
rect 70140 8766 70142 8818
rect 70194 8766 70196 8818
rect 69804 8652 69972 8708
rect 69916 7140 69972 8652
rect 70140 8596 70196 8766
rect 70140 8530 70196 8540
rect 70252 8708 70308 8718
rect 70140 8370 70196 8382
rect 70140 8318 70142 8370
rect 70194 8318 70196 8370
rect 70140 8260 70196 8318
rect 70140 8194 70196 8204
rect 70028 7586 70084 7598
rect 70028 7534 70030 7586
rect 70082 7534 70084 7586
rect 70028 7476 70084 7534
rect 70028 7410 70084 7420
rect 69916 7074 69972 7084
rect 69804 7028 69860 7038
rect 69804 6802 69860 6972
rect 69804 6750 69806 6802
rect 69858 6750 69860 6802
rect 69804 6738 69860 6750
rect 70028 6916 70084 6926
rect 69692 6524 69860 6580
rect 69580 6066 69636 6076
rect 69692 5796 69748 5806
rect 69468 4946 69524 4956
rect 69580 5236 69636 5246
rect 69468 4452 69524 4462
rect 69468 4226 69524 4396
rect 69468 4174 69470 4226
rect 69522 4174 69524 4226
rect 69468 4162 69524 4174
rect 69468 3556 69524 3566
rect 69580 3556 69636 5180
rect 69468 3554 69636 3556
rect 69468 3502 69470 3554
rect 69522 3502 69636 3554
rect 69468 3500 69636 3502
rect 69468 3490 69524 3500
rect 69692 3444 69748 5740
rect 69804 4900 69860 6524
rect 69804 4834 69860 4844
rect 69580 3388 69748 3444
rect 69804 4452 69860 4462
rect 69580 3332 69636 3388
rect 69804 3332 69860 4396
rect 69132 3042 69188 3052
rect 69244 3052 69412 3108
rect 69468 3276 69636 3332
rect 69692 3276 69860 3332
rect 69244 800 69300 3052
rect 69468 800 69524 3276
rect 69692 800 69748 3276
rect 70028 3108 70084 6860
rect 69916 3052 70084 3108
rect 70140 6020 70196 6030
rect 69916 800 69972 3052
rect 70140 800 70196 5964
rect 70252 4226 70308 8652
rect 70364 6578 70420 11118
rect 70476 10050 70532 11566
rect 70700 11172 70756 11182
rect 71260 11172 71316 11182
rect 71708 11172 71764 11182
rect 70700 11170 70868 11172
rect 70700 11118 70702 11170
rect 70754 11118 70868 11170
rect 70700 11116 70868 11118
rect 70700 11106 70756 11116
rect 70700 10722 70756 10734
rect 70700 10670 70702 10722
rect 70754 10670 70756 10722
rect 70700 10388 70756 10670
rect 70700 10322 70756 10332
rect 70476 9998 70478 10050
rect 70530 9998 70532 10050
rect 70476 9986 70532 9998
rect 70476 9828 70532 9838
rect 70476 9042 70532 9772
rect 70476 8990 70478 9042
rect 70530 8990 70532 9042
rect 70476 8978 70532 8990
rect 70588 9044 70644 9054
rect 70364 6526 70366 6578
rect 70418 6526 70420 6578
rect 70364 5124 70420 6526
rect 70476 6132 70532 6142
rect 70476 5684 70532 6076
rect 70588 5794 70644 8988
rect 70812 7924 70868 11116
rect 71260 11170 71652 11172
rect 71260 11118 71262 11170
rect 71314 11118 71652 11170
rect 71260 11116 71652 11118
rect 71260 11106 71316 11116
rect 71372 10722 71428 10734
rect 71372 10670 71374 10722
rect 71426 10670 71428 10722
rect 70924 10610 70980 10622
rect 70924 10558 70926 10610
rect 70978 10558 70980 10610
rect 70924 8484 70980 10558
rect 71260 9828 71316 9838
rect 71260 9734 71316 9772
rect 71036 9714 71092 9726
rect 71036 9662 71038 9714
rect 71090 9662 71092 9714
rect 71036 8708 71092 9662
rect 71372 9492 71428 10670
rect 71372 9426 71428 9436
rect 71484 9268 71540 9278
rect 71372 9212 71484 9268
rect 71260 9156 71316 9166
rect 71260 9062 71316 9100
rect 71148 9044 71204 9054
rect 71148 8950 71204 8988
rect 71036 8642 71092 8652
rect 71036 8484 71092 8494
rect 70924 8428 71036 8484
rect 71036 8418 71092 8428
rect 71260 8146 71316 8158
rect 71260 8094 71262 8146
rect 71314 8094 71316 8146
rect 70812 7868 70980 7924
rect 70924 7812 70980 7868
rect 70924 7756 71092 7812
rect 70588 5742 70590 5794
rect 70642 5742 70644 5794
rect 70588 5730 70644 5742
rect 70700 7700 70756 7710
rect 70476 5618 70532 5628
rect 70588 5236 70644 5246
rect 70588 5142 70644 5180
rect 70364 5058 70420 5068
rect 70476 5012 70532 5022
rect 70700 5012 70756 7644
rect 70812 7642 70868 7654
rect 70812 7590 70814 7642
rect 70866 7590 70868 7642
rect 70812 5908 70868 7590
rect 71036 6356 71092 7756
rect 71148 7476 71204 7486
rect 71148 7382 71204 7420
rect 70812 5842 70868 5852
rect 70924 6300 71092 6356
rect 71148 7252 71204 7262
rect 70924 5796 70980 6300
rect 71036 6132 71092 6142
rect 71036 6018 71092 6076
rect 71036 5966 71038 6018
rect 71090 5966 71092 6018
rect 71036 5954 71092 5966
rect 70924 5740 71092 5796
rect 70252 4174 70254 4226
rect 70306 4174 70308 4226
rect 70252 4162 70308 4174
rect 70364 4900 70420 4910
rect 70364 3444 70420 4844
rect 70252 3442 70420 3444
rect 70252 3390 70366 3442
rect 70418 3390 70420 3442
rect 70252 3388 70420 3390
rect 70252 2658 70308 3388
rect 70364 3378 70420 3388
rect 70476 3220 70532 4956
rect 70252 2606 70254 2658
rect 70306 2606 70308 2658
rect 70252 2594 70308 2606
rect 70364 3164 70532 3220
rect 70588 4956 70756 5012
rect 70812 5684 70868 5694
rect 70364 800 70420 3164
rect 70588 800 70644 4956
rect 70812 800 70868 5628
rect 70924 5572 70980 5582
rect 70924 4452 70980 5516
rect 70924 4386 70980 4396
rect 71036 4450 71092 5740
rect 71036 4398 71038 4450
rect 71090 4398 71092 4450
rect 71036 3780 71092 4398
rect 71036 3714 71092 3724
rect 71148 3388 71204 7196
rect 71260 7140 71316 8094
rect 71260 7074 71316 7084
rect 71260 5906 71316 5918
rect 71260 5854 71262 5906
rect 71314 5854 71316 5906
rect 71260 5234 71316 5854
rect 71260 5182 71262 5234
rect 71314 5182 71316 5234
rect 71260 5170 71316 5182
rect 71372 3388 71428 9212
rect 71484 9202 71540 9212
rect 71484 7586 71540 7598
rect 71484 7534 71486 7586
rect 71538 7534 71540 7586
rect 71484 6804 71540 7534
rect 71484 6738 71540 6748
rect 71036 3332 71204 3388
rect 71260 3332 71428 3388
rect 71484 4452 71540 4462
rect 71036 800 71092 3332
rect 71260 800 71316 3332
rect 71484 800 71540 4396
rect 71596 4340 71652 11116
rect 71708 11170 71876 11172
rect 71708 11118 71710 11170
rect 71762 11118 71876 11170
rect 71708 11116 71876 11118
rect 71708 11106 71764 11116
rect 71708 9602 71764 9614
rect 71708 9550 71710 9602
rect 71762 9550 71764 9602
rect 71708 9380 71764 9550
rect 71708 9314 71764 9324
rect 71708 8596 71764 8606
rect 71708 8036 71764 8540
rect 71820 8148 71876 11116
rect 72156 11170 72212 11182
rect 72156 11118 72158 11170
rect 72210 11118 72212 11170
rect 71932 10612 71988 10622
rect 71932 8596 71988 10556
rect 71932 8530 71988 8540
rect 72044 9714 72100 9726
rect 72044 9662 72046 9714
rect 72098 9662 72100 9714
rect 72044 8372 72100 9662
rect 72044 8306 72100 8316
rect 72044 8148 72100 8158
rect 71820 8146 72100 8148
rect 71820 8094 72046 8146
rect 72098 8094 72100 8146
rect 71820 8092 72100 8094
rect 71708 7980 71876 8036
rect 71596 4274 71652 4284
rect 71708 5460 71764 5470
rect 71708 2548 71764 5404
rect 71596 2492 71764 2548
rect 71820 2548 71876 7980
rect 71932 7364 71988 7374
rect 71932 4004 71988 7308
rect 72044 5012 72100 8092
rect 72156 7588 72212 11118
rect 72492 11172 72548 11182
rect 72492 11170 72772 11172
rect 72492 11118 72494 11170
rect 72546 11118 72772 11170
rect 72492 11116 72772 11118
rect 72492 11106 72548 11116
rect 72268 10722 72324 10734
rect 72268 10670 72270 10722
rect 72322 10670 72324 10722
rect 72268 9268 72324 10670
rect 72604 9828 72660 9838
rect 72492 9826 72660 9828
rect 72492 9774 72606 9826
rect 72658 9774 72660 9826
rect 72492 9772 72660 9774
rect 72380 9604 72436 9614
rect 72380 9510 72436 9548
rect 72268 9202 72324 9212
rect 72268 8932 72324 8942
rect 72268 8838 72324 8876
rect 72380 7588 72436 7598
rect 72156 7586 72436 7588
rect 72156 7534 72382 7586
rect 72434 7534 72436 7586
rect 72156 7532 72436 7534
rect 72380 7252 72436 7532
rect 72380 7186 72436 7196
rect 72492 6916 72548 9772
rect 72604 9762 72660 9772
rect 72604 9492 72660 9502
rect 72604 7700 72660 9436
rect 72604 7634 72660 7644
rect 72268 6860 72548 6916
rect 72604 7476 72660 7486
rect 72268 6692 72324 6860
rect 72044 4946 72100 4956
rect 72156 6636 72324 6692
rect 72380 6692 72436 6702
rect 72156 4562 72212 6636
rect 72380 6020 72436 6636
rect 72380 5926 72436 5964
rect 72156 4510 72158 4562
rect 72210 4510 72212 4562
rect 72156 4498 72212 4510
rect 72380 5236 72436 5246
rect 71932 3948 72100 4004
rect 71596 2324 71652 2492
rect 71820 2482 71876 2492
rect 71932 3780 71988 3790
rect 71596 2268 71764 2324
rect 71708 800 71764 2268
rect 71932 800 71988 3724
rect 72044 3332 72100 3948
rect 72044 3266 72100 3276
rect 72156 3444 72212 3454
rect 72156 800 72212 3388
rect 72380 800 72436 5180
rect 72492 4676 72548 4686
rect 72492 3388 72548 4620
rect 72604 3666 72660 7420
rect 72716 6692 72772 11116
rect 72940 11170 72996 11182
rect 73836 11172 73892 11182
rect 72940 11118 72942 11170
rect 72994 11118 72996 11170
rect 72828 10612 72884 10622
rect 72828 10518 72884 10556
rect 72940 9716 72996 11118
rect 73724 11170 73892 11172
rect 73724 11118 73838 11170
rect 73890 11118 73892 11170
rect 73724 11116 73892 11118
rect 73276 10498 73332 10510
rect 73276 10446 73278 10498
rect 73330 10446 73332 10498
rect 72828 9660 72996 9716
rect 73052 9714 73108 9726
rect 73052 9662 73054 9714
rect 73106 9662 73108 9714
rect 72828 7140 72884 9660
rect 73052 9604 73108 9662
rect 72940 9548 73108 9604
rect 72940 8932 72996 9548
rect 73276 9380 73332 10446
rect 73724 9828 73780 11116
rect 73836 11106 73892 11116
rect 76748 11004 77028 11060
rect 73836 10498 73892 10510
rect 73836 10446 73838 10498
rect 73890 10446 73892 10498
rect 73836 9940 73892 10446
rect 74172 10498 74228 10510
rect 74172 10446 74174 10498
rect 74226 10446 74228 10498
rect 74172 10386 74228 10446
rect 74172 10334 74174 10386
rect 74226 10334 74228 10386
rect 74172 10322 74228 10334
rect 74620 10498 74676 10510
rect 75180 10500 75236 10510
rect 75964 10500 76020 10510
rect 74620 10446 74622 10498
rect 74674 10446 74676 10498
rect 73836 9884 74228 9940
rect 73724 9772 73892 9828
rect 72940 8866 72996 8876
rect 73052 9324 73332 9380
rect 73388 9602 73444 9614
rect 73724 9604 73780 9614
rect 73388 9550 73390 9602
rect 73442 9550 73444 9602
rect 72828 7074 72884 7084
rect 72828 6804 72884 6814
rect 72828 6710 72884 6748
rect 73052 6692 73108 9324
rect 73276 9154 73332 9166
rect 73276 9102 73278 9154
rect 73330 9102 73332 9154
rect 73276 8596 73332 9102
rect 73388 8820 73444 9550
rect 73388 8754 73444 8764
rect 73500 9602 73780 9604
rect 73500 9550 73726 9602
rect 73778 9550 73780 9602
rect 73500 9548 73780 9550
rect 73276 8530 73332 8540
rect 73164 8372 73220 8382
rect 73500 8372 73556 9548
rect 73724 9538 73780 9548
rect 73836 9156 73892 9772
rect 73724 9100 73892 9156
rect 74060 9714 74116 9726
rect 74060 9662 74062 9714
rect 74114 9662 74116 9714
rect 73724 8932 73780 9100
rect 73724 8876 74004 8932
rect 73164 8278 73220 8316
rect 73276 8316 73556 8372
rect 73724 8484 73780 8494
rect 73724 8370 73780 8428
rect 73724 8318 73726 8370
rect 73778 8318 73780 8370
rect 73276 7364 73332 8316
rect 73724 8306 73780 8318
rect 73276 7298 73332 7308
rect 73388 8036 73444 8046
rect 73164 6692 73220 6702
rect 73052 6636 73164 6692
rect 72716 6626 72772 6636
rect 73164 6626 73220 6636
rect 73276 6132 73332 6142
rect 73052 6076 73276 6132
rect 72828 5908 72884 5918
rect 72828 5684 72884 5852
rect 72828 5618 72884 5628
rect 72604 3614 72606 3666
rect 72658 3614 72660 3666
rect 72604 3602 72660 3614
rect 72828 5012 72884 5022
rect 72492 3332 72660 3388
rect 72604 800 72660 3332
rect 72828 800 72884 4956
rect 73052 800 73108 6076
rect 73276 6066 73332 6076
rect 73276 5124 73332 5134
rect 73164 5010 73220 5022
rect 73164 4958 73166 5010
rect 73218 4958 73220 5010
rect 73164 4340 73220 4958
rect 73164 4274 73220 4284
rect 73164 3330 73220 3342
rect 73164 3278 73166 3330
rect 73218 3278 73220 3330
rect 73164 2884 73220 3278
rect 73164 2818 73220 2828
rect 73276 800 73332 5068
rect 73388 3220 73444 7980
rect 73724 7364 73780 7374
rect 73724 7270 73780 7308
rect 73724 7140 73780 7150
rect 73612 6692 73668 6702
rect 73500 6580 73556 6590
rect 73612 6580 73668 6636
rect 73500 6578 73668 6580
rect 73500 6526 73502 6578
rect 73554 6526 73668 6578
rect 73500 6524 73668 6526
rect 73500 6514 73556 6524
rect 73612 5908 73668 6524
rect 73612 5842 73668 5852
rect 73724 5572 73780 7084
rect 73612 5516 73780 5572
rect 73612 4116 73668 5516
rect 73836 4564 73892 4574
rect 73948 4564 74004 8876
rect 74060 5234 74116 9662
rect 74172 9154 74228 9884
rect 74396 9604 74452 9614
rect 74172 9102 74174 9154
rect 74226 9102 74228 9154
rect 74172 6580 74228 9102
rect 74172 6514 74228 6524
rect 74284 9602 74452 9604
rect 74284 9550 74398 9602
rect 74450 9550 74452 9602
rect 74284 9548 74452 9550
rect 74060 5182 74062 5234
rect 74114 5182 74116 5234
rect 74060 5170 74116 5182
rect 74284 4676 74340 9548
rect 74396 9538 74452 9548
rect 74508 9604 74564 9614
rect 74508 9044 74564 9548
rect 74396 8988 74564 9044
rect 74396 7586 74452 8988
rect 74396 7534 74398 7586
rect 74450 7534 74452 7586
rect 74396 5012 74452 7534
rect 74508 8820 74564 8830
rect 74508 5794 74564 8764
rect 74508 5742 74510 5794
rect 74562 5742 74564 5794
rect 74508 5730 74564 5742
rect 74620 5012 74676 10446
rect 75068 10498 75236 10500
rect 75068 10446 75182 10498
rect 75234 10446 75236 10498
rect 75068 10444 75236 10446
rect 74732 10386 74788 10398
rect 74732 10334 74734 10386
rect 74786 10334 74788 10386
rect 74732 8146 74788 10334
rect 74956 9604 75012 9614
rect 74956 9510 75012 9548
rect 74732 8094 74734 8146
rect 74786 8094 74788 8146
rect 74732 5572 74788 8094
rect 74732 5506 74788 5516
rect 74956 5012 75012 5022
rect 74620 5010 75012 5012
rect 74620 4958 74958 5010
rect 75010 4958 75012 5010
rect 74620 4956 75012 4958
rect 74396 4946 74452 4956
rect 74284 4610 74340 4620
rect 73892 4508 74004 4564
rect 73836 4498 73892 4508
rect 73612 4050 73668 4060
rect 74284 4450 74340 4462
rect 74284 4398 74286 4450
rect 74338 4398 74340 4450
rect 74284 4116 74340 4398
rect 74284 4050 74340 4060
rect 74956 3556 75012 4956
rect 75068 4452 75124 10444
rect 75180 10434 75236 10444
rect 75740 10498 76020 10500
rect 75740 10446 75966 10498
rect 76018 10446 76020 10498
rect 75740 10444 76020 10446
rect 75628 9716 75684 9726
rect 75404 9602 75460 9614
rect 75404 9550 75406 9602
rect 75458 9550 75460 9602
rect 75404 8428 75460 9550
rect 75516 8932 75572 8942
rect 75628 8932 75684 9660
rect 75516 8930 75684 8932
rect 75516 8878 75518 8930
rect 75570 8878 75684 8930
rect 75516 8876 75684 8878
rect 75516 8866 75572 8876
rect 75180 8372 75460 8428
rect 75180 6018 75236 8372
rect 75516 8034 75572 8046
rect 75516 7982 75518 8034
rect 75570 7982 75572 8034
rect 75516 6916 75572 7982
rect 75516 6850 75572 6860
rect 75628 7476 75684 7486
rect 75628 6914 75684 7420
rect 75628 6862 75630 6914
rect 75682 6862 75684 6914
rect 75628 6850 75684 6862
rect 75740 6580 75796 10444
rect 75964 10434 76020 10444
rect 76636 10498 76692 10510
rect 76636 10446 76638 10498
rect 76690 10446 76692 10498
rect 75852 9828 75908 9838
rect 75852 9266 75908 9772
rect 76188 9604 76244 9614
rect 75852 9214 75854 9266
rect 75906 9214 75908 9266
rect 75852 9202 75908 9214
rect 75964 9602 76244 9604
rect 75964 9550 76190 9602
rect 76242 9550 76244 9602
rect 75964 9548 76244 9550
rect 75740 6514 75796 6524
rect 75180 5966 75182 6018
rect 75234 5966 75236 6018
rect 75180 5684 75236 5966
rect 75180 5618 75236 5628
rect 75628 6020 75684 6030
rect 75180 4452 75236 4462
rect 75068 4396 75180 4452
rect 75180 4358 75236 4396
rect 74956 3490 75012 3500
rect 73500 3444 73556 3454
rect 73948 3444 74004 3454
rect 73500 3442 74004 3444
rect 73500 3390 73502 3442
rect 73554 3390 73950 3442
rect 74002 3390 74004 3442
rect 73500 3388 74004 3390
rect 73500 3378 73556 3388
rect 73948 3378 74004 3388
rect 75628 3220 75684 5964
rect 75964 5124 76020 9548
rect 76188 9538 76244 9548
rect 76636 9268 76692 10446
rect 76636 9202 76692 9212
rect 76188 9044 76244 9054
rect 76188 9042 76580 9044
rect 76188 8990 76190 9042
rect 76242 8990 76580 9042
rect 76188 8988 76580 8990
rect 76188 8978 76244 8988
rect 76188 8708 76244 8718
rect 76188 8370 76244 8652
rect 76188 8318 76190 8370
rect 76242 8318 76244 8370
rect 76188 8306 76244 8318
rect 76188 8148 76244 8158
rect 76188 5234 76244 8092
rect 76524 7362 76580 8988
rect 76524 7310 76526 7362
rect 76578 7310 76580 7362
rect 76524 7298 76580 7310
rect 76188 5182 76190 5234
rect 76242 5182 76244 5234
rect 76188 5170 76244 5182
rect 76300 6580 76356 6590
rect 76300 5236 76356 6524
rect 76748 5908 76804 11004
rect 76860 10836 76916 10846
rect 76860 9714 76916 10780
rect 76972 10834 77028 11004
rect 78492 11004 78756 11014
rect 77308 10948 77364 10958
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 77364 10892 77476 10948
rect 78492 10938 78756 10948
rect 77308 10882 77364 10892
rect 76972 10782 76974 10834
rect 77026 10782 77028 10834
rect 76972 10770 77028 10782
rect 77196 9716 77252 9726
rect 76860 9662 76862 9714
rect 76914 9662 76916 9714
rect 76860 9650 76916 9662
rect 76972 9714 77252 9716
rect 76972 9662 77198 9714
rect 77250 9662 77252 9714
rect 76972 9660 77252 9662
rect 77420 9716 77476 10892
rect 77868 10724 77924 10734
rect 77532 10722 77924 10724
rect 77532 10670 77870 10722
rect 77922 10670 77924 10722
rect 77532 10668 77924 10670
rect 77532 9940 77588 10668
rect 77868 10658 77924 10668
rect 78204 10612 78260 10622
rect 78204 10610 78484 10612
rect 78204 10558 78206 10610
rect 78258 10558 78484 10610
rect 78204 10556 78484 10558
rect 78204 10546 78260 10556
rect 77644 10500 77700 10510
rect 77644 10498 78148 10500
rect 77644 10446 77646 10498
rect 77698 10446 78148 10498
rect 77644 10444 78148 10446
rect 77644 10434 77700 10444
rect 78092 10052 78148 10444
rect 78092 9996 78372 10052
rect 77532 9874 77588 9884
rect 78092 9828 78148 9838
rect 77980 9826 78148 9828
rect 77980 9774 78094 9826
rect 78146 9774 78148 9826
rect 77980 9772 78148 9774
rect 77868 9716 77924 9726
rect 77420 9714 77924 9716
rect 77420 9662 77870 9714
rect 77922 9662 77924 9714
rect 77420 9660 77924 9662
rect 76860 9156 76916 9166
rect 76860 9062 76916 9100
rect 76748 5842 76804 5852
rect 76860 7588 76916 7598
rect 76300 5170 76356 5180
rect 75964 5058 76020 5068
rect 76076 4564 76132 4574
rect 76076 3442 76132 4508
rect 76076 3390 76078 3442
rect 76130 3390 76132 3442
rect 76076 3378 76132 3390
rect 76860 3442 76916 7532
rect 76972 7028 77028 9660
rect 77196 9650 77252 9660
rect 77868 9650 77924 9660
rect 77084 9268 77140 9278
rect 77084 9042 77140 9212
rect 77532 9154 77588 9166
rect 77532 9102 77534 9154
rect 77586 9102 77588 9154
rect 77084 8990 77086 9042
rect 77138 8990 77140 9042
rect 77084 8428 77140 8990
rect 77420 9044 77476 9054
rect 77084 8372 77252 8428
rect 77084 7924 77140 7934
rect 77084 7698 77140 7868
rect 77084 7646 77086 7698
rect 77138 7646 77140 7698
rect 77084 7634 77140 7646
rect 76972 6962 77028 6972
rect 77084 6804 77140 6814
rect 77084 3554 77140 6748
rect 77196 5460 77252 8372
rect 77196 5394 77252 5404
rect 77308 7474 77364 7486
rect 77308 7422 77310 7474
rect 77362 7422 77364 7474
rect 77308 4226 77364 7422
rect 77308 4174 77310 4226
rect 77362 4174 77364 4226
rect 77308 4162 77364 4174
rect 77420 4228 77476 8988
rect 77532 8146 77588 9102
rect 77756 9042 77812 9054
rect 77756 8990 77758 9042
rect 77810 8990 77812 9042
rect 77756 8428 77812 8990
rect 77980 8428 78036 9772
rect 78092 9762 78148 9772
rect 77532 8094 77534 8146
rect 77586 8094 77588 8146
rect 77532 8082 77588 8094
rect 77644 8372 77812 8428
rect 77868 8372 78036 8428
rect 78092 8372 78148 8382
rect 77532 7140 77588 7150
rect 77532 5348 77588 7084
rect 77644 6802 77700 8372
rect 77756 7586 77812 7598
rect 77756 7534 77758 7586
rect 77810 7534 77812 7586
rect 77756 7252 77812 7534
rect 77756 7186 77812 7196
rect 77868 7028 77924 8372
rect 78148 8316 78260 8372
rect 78092 8306 78148 8316
rect 77980 8036 78036 8046
rect 77980 7942 78036 7980
rect 77980 7476 78036 7486
rect 77980 7382 78036 7420
rect 77644 6750 77646 6802
rect 77698 6750 77700 6802
rect 77644 6738 77700 6750
rect 77756 6972 77924 7028
rect 78092 7364 78148 7374
rect 77644 6132 77700 6142
rect 77756 6132 77812 6972
rect 77980 6468 78036 6478
rect 77980 6374 78036 6412
rect 77644 6130 77812 6132
rect 77644 6078 77646 6130
rect 77698 6078 77812 6130
rect 77644 6076 77812 6078
rect 77644 6066 77700 6076
rect 77868 6020 77924 6030
rect 77868 5926 77924 5964
rect 77532 5282 77588 5292
rect 77644 5908 77700 5918
rect 77532 5012 77588 5022
rect 77644 5012 77700 5852
rect 78092 5906 78148 7308
rect 78092 5854 78094 5906
rect 78146 5854 78148 5906
rect 78092 5842 78148 5854
rect 77532 5010 77700 5012
rect 77532 4958 77534 5010
rect 77586 4958 77700 5010
rect 77532 4956 77700 4958
rect 77532 4946 77588 4956
rect 77980 4900 78036 4910
rect 77980 4898 78148 4900
rect 77980 4846 77982 4898
rect 78034 4846 78148 4898
rect 77980 4844 78148 4846
rect 77980 4834 78036 4844
rect 77868 4452 77924 4462
rect 77868 4450 78036 4452
rect 77868 4398 77870 4450
rect 77922 4398 78036 4450
rect 77868 4396 78036 4398
rect 77868 4386 77924 4396
rect 77420 4172 77924 4228
rect 77084 3502 77086 3554
rect 77138 3502 77140 3554
rect 77084 3490 77140 3502
rect 76860 3390 76862 3442
rect 76914 3390 76916 3442
rect 76860 3378 76916 3390
rect 77868 3442 77924 4172
rect 77868 3390 77870 3442
rect 77922 3390 77924 3442
rect 77868 3378 77924 3390
rect 73388 3164 73556 3220
rect 73500 800 73556 3164
rect 75628 3154 75684 3164
rect 77980 2996 78036 4396
rect 78092 3780 78148 4844
rect 78204 4450 78260 8316
rect 78204 4398 78206 4450
rect 78258 4398 78260 4450
rect 78204 4386 78260 4398
rect 78092 3714 78148 3724
rect 78092 3556 78148 3566
rect 78316 3556 78372 9996
rect 78428 9716 78484 10556
rect 78428 9650 78484 9660
rect 78492 9436 78756 9446
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78492 9370 78756 9380
rect 78492 7868 78756 7878
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78492 7802 78756 7812
rect 78492 6300 78756 6310
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78492 6234 78756 6244
rect 78492 4732 78756 4742
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78492 4666 78756 4676
rect 78092 3554 78372 3556
rect 78092 3502 78094 3554
rect 78146 3502 78372 3554
rect 78092 3500 78372 3502
rect 78092 3444 78148 3500
rect 78092 3378 78148 3388
rect 78492 3164 78756 3174
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78492 3098 78756 3108
rect 77980 2930 78036 2940
rect 6272 0 6384 800
rect 6496 0 6608 800
rect 6720 0 6832 800
rect 6944 0 7056 800
rect 7168 0 7280 800
rect 7392 0 7504 800
rect 7616 0 7728 800
rect 7840 0 7952 800
rect 8064 0 8176 800
rect 8288 0 8400 800
rect 8512 0 8624 800
rect 8736 0 8848 800
rect 8960 0 9072 800
rect 9184 0 9296 800
rect 9408 0 9520 800
rect 9632 0 9744 800
rect 9856 0 9968 800
rect 10080 0 10192 800
rect 10304 0 10416 800
rect 10528 0 10640 800
rect 10752 0 10864 800
rect 10976 0 11088 800
rect 11200 0 11312 800
rect 11424 0 11536 800
rect 11648 0 11760 800
rect 11872 0 11984 800
rect 12096 0 12208 800
rect 12320 0 12432 800
rect 12544 0 12656 800
rect 12768 0 12880 800
rect 12992 0 13104 800
rect 13216 0 13328 800
rect 13440 0 13552 800
rect 13664 0 13776 800
rect 13888 0 14000 800
rect 14112 0 14224 800
rect 14336 0 14448 800
rect 14560 0 14672 800
rect 14784 0 14896 800
rect 15008 0 15120 800
rect 15232 0 15344 800
rect 15456 0 15568 800
rect 15680 0 15792 800
rect 15904 0 16016 800
rect 16128 0 16240 800
rect 16352 0 16464 800
rect 16576 0 16688 800
rect 16800 0 16912 800
rect 17024 0 17136 800
rect 17248 0 17360 800
rect 17472 0 17584 800
rect 17696 0 17808 800
rect 17920 0 18032 800
rect 18144 0 18256 800
rect 18368 0 18480 800
rect 18592 0 18704 800
rect 18816 0 18928 800
rect 19040 0 19152 800
rect 19264 0 19376 800
rect 19488 0 19600 800
rect 19712 0 19824 800
rect 19936 0 20048 800
rect 20160 0 20272 800
rect 20384 0 20496 800
rect 20608 0 20720 800
rect 20832 0 20944 800
rect 21056 0 21168 800
rect 21280 0 21392 800
rect 21504 0 21616 800
rect 21728 0 21840 800
rect 21952 0 22064 800
rect 22176 0 22288 800
rect 22400 0 22512 800
rect 22624 0 22736 800
rect 22848 0 22960 800
rect 23072 0 23184 800
rect 23296 0 23408 800
rect 23520 0 23632 800
rect 23744 0 23856 800
rect 23968 0 24080 800
rect 24192 0 24304 800
rect 24416 0 24528 800
rect 24640 0 24752 800
rect 24864 0 24976 800
rect 25088 0 25200 800
rect 25312 0 25424 800
rect 25536 0 25648 800
rect 25760 0 25872 800
rect 25984 0 26096 800
rect 26208 0 26320 800
rect 26432 0 26544 800
rect 26656 0 26768 800
rect 26880 0 26992 800
rect 27104 0 27216 800
rect 27328 0 27440 800
rect 27552 0 27664 800
rect 27776 0 27888 800
rect 28000 0 28112 800
rect 28224 0 28336 800
rect 28448 0 28560 800
rect 28672 0 28784 800
rect 28896 0 29008 800
rect 29120 0 29232 800
rect 29344 0 29456 800
rect 29568 0 29680 800
rect 29792 0 29904 800
rect 30016 0 30128 800
rect 30240 0 30352 800
rect 30464 0 30576 800
rect 30688 0 30800 800
rect 30912 0 31024 800
rect 31136 0 31248 800
rect 31360 0 31472 800
rect 31584 0 31696 800
rect 31808 0 31920 800
rect 32032 0 32144 800
rect 32256 0 32368 800
rect 32480 0 32592 800
rect 32704 0 32816 800
rect 32928 0 33040 800
rect 33152 0 33264 800
rect 33376 0 33488 800
rect 33600 0 33712 800
rect 33824 0 33936 800
rect 34048 0 34160 800
rect 34272 0 34384 800
rect 34496 0 34608 800
rect 34720 0 34832 800
rect 34944 0 35056 800
rect 35168 0 35280 800
rect 35392 0 35504 800
rect 35616 0 35728 800
rect 35840 0 35952 800
rect 36064 0 36176 800
rect 36288 0 36400 800
rect 36512 0 36624 800
rect 36736 0 36848 800
rect 36960 0 37072 800
rect 37184 0 37296 800
rect 37408 0 37520 800
rect 37632 0 37744 800
rect 37856 0 37968 800
rect 38080 0 38192 800
rect 38304 0 38416 800
rect 38528 0 38640 800
rect 38752 0 38864 800
rect 38976 0 39088 800
rect 39200 0 39312 800
rect 39424 0 39536 800
rect 39648 0 39760 800
rect 39872 0 39984 800
rect 40096 0 40208 800
rect 40320 0 40432 800
rect 40544 0 40656 800
rect 40768 0 40880 800
rect 40992 0 41104 800
rect 41216 0 41328 800
rect 41440 0 41552 800
rect 41664 0 41776 800
rect 41888 0 42000 800
rect 42112 0 42224 800
rect 42336 0 42448 800
rect 42560 0 42672 800
rect 42784 0 42896 800
rect 43008 0 43120 800
rect 43232 0 43344 800
rect 43456 0 43568 800
rect 43680 0 43792 800
rect 43904 0 44016 800
rect 44128 0 44240 800
rect 44352 0 44464 800
rect 44576 0 44688 800
rect 44800 0 44912 800
rect 45024 0 45136 800
rect 45248 0 45360 800
rect 45472 0 45584 800
rect 45696 0 45808 800
rect 45920 0 46032 800
rect 46144 0 46256 800
rect 46368 0 46480 800
rect 46592 0 46704 800
rect 46816 0 46928 800
rect 47040 0 47152 800
rect 47264 0 47376 800
rect 47488 0 47600 800
rect 47712 0 47824 800
rect 47936 0 48048 800
rect 48160 0 48272 800
rect 48384 0 48496 800
rect 48608 0 48720 800
rect 48832 0 48944 800
rect 49056 0 49168 800
rect 49280 0 49392 800
rect 49504 0 49616 800
rect 49728 0 49840 800
rect 49952 0 50064 800
rect 50176 0 50288 800
rect 50400 0 50512 800
rect 50624 0 50736 800
rect 50848 0 50960 800
rect 51072 0 51184 800
rect 51296 0 51408 800
rect 51520 0 51632 800
rect 51744 0 51856 800
rect 51968 0 52080 800
rect 52192 0 52304 800
rect 52416 0 52528 800
rect 52640 0 52752 800
rect 52864 0 52976 800
rect 53088 0 53200 800
rect 53312 0 53424 800
rect 53536 0 53648 800
rect 53760 0 53872 800
rect 53984 0 54096 800
rect 54208 0 54320 800
rect 54432 0 54544 800
rect 54656 0 54768 800
rect 54880 0 54992 800
rect 55104 0 55216 800
rect 55328 0 55440 800
rect 55552 0 55664 800
rect 55776 0 55888 800
rect 56000 0 56112 800
rect 56224 0 56336 800
rect 56448 0 56560 800
rect 56672 0 56784 800
rect 56896 0 57008 800
rect 57120 0 57232 800
rect 57344 0 57456 800
rect 57568 0 57680 800
rect 57792 0 57904 800
rect 58016 0 58128 800
rect 58240 0 58352 800
rect 58464 0 58576 800
rect 58688 0 58800 800
rect 58912 0 59024 800
rect 59136 0 59248 800
rect 59360 0 59472 800
rect 59584 0 59696 800
rect 59808 0 59920 800
rect 60032 0 60144 800
rect 60256 0 60368 800
rect 60480 0 60592 800
rect 60704 0 60816 800
rect 60928 0 61040 800
rect 61152 0 61264 800
rect 61376 0 61488 800
rect 61600 0 61712 800
rect 61824 0 61936 800
rect 62048 0 62160 800
rect 62272 0 62384 800
rect 62496 0 62608 800
rect 62720 0 62832 800
rect 62944 0 63056 800
rect 63168 0 63280 800
rect 63392 0 63504 800
rect 63616 0 63728 800
rect 63840 0 63952 800
rect 64064 0 64176 800
rect 64288 0 64400 800
rect 64512 0 64624 800
rect 64736 0 64848 800
rect 64960 0 65072 800
rect 65184 0 65296 800
rect 65408 0 65520 800
rect 65632 0 65744 800
rect 65856 0 65968 800
rect 66080 0 66192 800
rect 66304 0 66416 800
rect 66528 0 66640 800
rect 66752 0 66864 800
rect 66976 0 67088 800
rect 67200 0 67312 800
rect 67424 0 67536 800
rect 67648 0 67760 800
rect 67872 0 67984 800
rect 68096 0 68208 800
rect 68320 0 68432 800
rect 68544 0 68656 800
rect 68768 0 68880 800
rect 68992 0 69104 800
rect 69216 0 69328 800
rect 69440 0 69552 800
rect 69664 0 69776 800
rect 69888 0 70000 800
rect 70112 0 70224 800
rect 70336 0 70448 800
rect 70560 0 70672 800
rect 70784 0 70896 800
rect 71008 0 71120 800
rect 71232 0 71344 800
rect 71456 0 71568 800
rect 71680 0 71792 800
rect 71904 0 72016 800
rect 72128 0 72240 800
rect 72352 0 72464 800
rect 72576 0 72688 800
rect 72800 0 72912 800
rect 73024 0 73136 800
rect 73248 0 73360 800
rect 73472 0 73584 800
<< via2 >>
rect 10872 36874 10928 36876
rect 10872 36822 10874 36874
rect 10874 36822 10926 36874
rect 10926 36822 10928 36874
rect 10872 36820 10928 36822
rect 10976 36874 11032 36876
rect 10976 36822 10978 36874
rect 10978 36822 11030 36874
rect 11030 36822 11032 36874
rect 10976 36820 11032 36822
rect 11080 36874 11136 36876
rect 11080 36822 11082 36874
rect 11082 36822 11134 36874
rect 11134 36822 11136 36874
rect 11080 36820 11136 36822
rect 30192 36874 30248 36876
rect 30192 36822 30194 36874
rect 30194 36822 30246 36874
rect 30246 36822 30248 36874
rect 30192 36820 30248 36822
rect 30296 36874 30352 36876
rect 30296 36822 30298 36874
rect 30298 36822 30350 36874
rect 30350 36822 30352 36874
rect 30296 36820 30352 36822
rect 30400 36874 30456 36876
rect 30400 36822 30402 36874
rect 30402 36822 30454 36874
rect 30454 36822 30456 36874
rect 30400 36820 30456 36822
rect 49512 36874 49568 36876
rect 49512 36822 49514 36874
rect 49514 36822 49566 36874
rect 49566 36822 49568 36874
rect 49512 36820 49568 36822
rect 49616 36874 49672 36876
rect 49616 36822 49618 36874
rect 49618 36822 49670 36874
rect 49670 36822 49672 36874
rect 49616 36820 49672 36822
rect 49720 36874 49776 36876
rect 49720 36822 49722 36874
rect 49722 36822 49774 36874
rect 49774 36822 49776 36874
rect 49720 36820 49776 36822
rect 68832 36874 68888 36876
rect 68832 36822 68834 36874
rect 68834 36822 68886 36874
rect 68886 36822 68888 36874
rect 68832 36820 68888 36822
rect 68936 36874 68992 36876
rect 68936 36822 68938 36874
rect 68938 36822 68990 36874
rect 68990 36822 68992 36874
rect 68936 36820 68992 36822
rect 69040 36874 69096 36876
rect 69040 36822 69042 36874
rect 69042 36822 69094 36874
rect 69094 36822 69096 36874
rect 69040 36820 69096 36822
rect 20532 36090 20588 36092
rect 20532 36038 20534 36090
rect 20534 36038 20586 36090
rect 20586 36038 20588 36090
rect 20532 36036 20588 36038
rect 20636 36090 20692 36092
rect 20636 36038 20638 36090
rect 20638 36038 20690 36090
rect 20690 36038 20692 36090
rect 20636 36036 20692 36038
rect 20740 36090 20796 36092
rect 20740 36038 20742 36090
rect 20742 36038 20794 36090
rect 20794 36038 20796 36090
rect 20740 36036 20796 36038
rect 39852 36090 39908 36092
rect 39852 36038 39854 36090
rect 39854 36038 39906 36090
rect 39906 36038 39908 36090
rect 39852 36036 39908 36038
rect 39956 36090 40012 36092
rect 39956 36038 39958 36090
rect 39958 36038 40010 36090
rect 40010 36038 40012 36090
rect 39956 36036 40012 36038
rect 40060 36090 40116 36092
rect 40060 36038 40062 36090
rect 40062 36038 40114 36090
rect 40114 36038 40116 36090
rect 40060 36036 40116 36038
rect 59172 36090 59228 36092
rect 59172 36038 59174 36090
rect 59174 36038 59226 36090
rect 59226 36038 59228 36090
rect 59172 36036 59228 36038
rect 59276 36090 59332 36092
rect 59276 36038 59278 36090
rect 59278 36038 59330 36090
rect 59330 36038 59332 36090
rect 59276 36036 59332 36038
rect 59380 36090 59436 36092
rect 59380 36038 59382 36090
rect 59382 36038 59434 36090
rect 59434 36038 59436 36090
rect 59380 36036 59436 36038
rect 78492 36090 78548 36092
rect 78492 36038 78494 36090
rect 78494 36038 78546 36090
rect 78546 36038 78548 36090
rect 78492 36036 78548 36038
rect 78596 36090 78652 36092
rect 78596 36038 78598 36090
rect 78598 36038 78650 36090
rect 78650 36038 78652 36090
rect 78596 36036 78652 36038
rect 78700 36090 78756 36092
rect 78700 36038 78702 36090
rect 78702 36038 78754 36090
rect 78754 36038 78756 36090
rect 78700 36036 78756 36038
rect 10872 35306 10928 35308
rect 10872 35254 10874 35306
rect 10874 35254 10926 35306
rect 10926 35254 10928 35306
rect 10872 35252 10928 35254
rect 10976 35306 11032 35308
rect 10976 35254 10978 35306
rect 10978 35254 11030 35306
rect 11030 35254 11032 35306
rect 10976 35252 11032 35254
rect 11080 35306 11136 35308
rect 11080 35254 11082 35306
rect 11082 35254 11134 35306
rect 11134 35254 11136 35306
rect 11080 35252 11136 35254
rect 30192 35306 30248 35308
rect 30192 35254 30194 35306
rect 30194 35254 30246 35306
rect 30246 35254 30248 35306
rect 30192 35252 30248 35254
rect 30296 35306 30352 35308
rect 30296 35254 30298 35306
rect 30298 35254 30350 35306
rect 30350 35254 30352 35306
rect 30296 35252 30352 35254
rect 30400 35306 30456 35308
rect 30400 35254 30402 35306
rect 30402 35254 30454 35306
rect 30454 35254 30456 35306
rect 30400 35252 30456 35254
rect 49512 35306 49568 35308
rect 49512 35254 49514 35306
rect 49514 35254 49566 35306
rect 49566 35254 49568 35306
rect 49512 35252 49568 35254
rect 49616 35306 49672 35308
rect 49616 35254 49618 35306
rect 49618 35254 49670 35306
rect 49670 35254 49672 35306
rect 49616 35252 49672 35254
rect 49720 35306 49776 35308
rect 49720 35254 49722 35306
rect 49722 35254 49774 35306
rect 49774 35254 49776 35306
rect 49720 35252 49776 35254
rect 68832 35306 68888 35308
rect 68832 35254 68834 35306
rect 68834 35254 68886 35306
rect 68886 35254 68888 35306
rect 68832 35252 68888 35254
rect 68936 35306 68992 35308
rect 68936 35254 68938 35306
rect 68938 35254 68990 35306
rect 68990 35254 68992 35306
rect 68936 35252 68992 35254
rect 69040 35306 69096 35308
rect 69040 35254 69042 35306
rect 69042 35254 69094 35306
rect 69094 35254 69096 35306
rect 69040 35252 69096 35254
rect 20532 34522 20588 34524
rect 20532 34470 20534 34522
rect 20534 34470 20586 34522
rect 20586 34470 20588 34522
rect 20532 34468 20588 34470
rect 20636 34522 20692 34524
rect 20636 34470 20638 34522
rect 20638 34470 20690 34522
rect 20690 34470 20692 34522
rect 20636 34468 20692 34470
rect 20740 34522 20796 34524
rect 20740 34470 20742 34522
rect 20742 34470 20794 34522
rect 20794 34470 20796 34522
rect 20740 34468 20796 34470
rect 39852 34522 39908 34524
rect 39852 34470 39854 34522
rect 39854 34470 39906 34522
rect 39906 34470 39908 34522
rect 39852 34468 39908 34470
rect 39956 34522 40012 34524
rect 39956 34470 39958 34522
rect 39958 34470 40010 34522
rect 40010 34470 40012 34522
rect 39956 34468 40012 34470
rect 40060 34522 40116 34524
rect 40060 34470 40062 34522
rect 40062 34470 40114 34522
rect 40114 34470 40116 34522
rect 40060 34468 40116 34470
rect 59172 34522 59228 34524
rect 59172 34470 59174 34522
rect 59174 34470 59226 34522
rect 59226 34470 59228 34522
rect 59172 34468 59228 34470
rect 59276 34522 59332 34524
rect 59276 34470 59278 34522
rect 59278 34470 59330 34522
rect 59330 34470 59332 34522
rect 59276 34468 59332 34470
rect 59380 34522 59436 34524
rect 59380 34470 59382 34522
rect 59382 34470 59434 34522
rect 59434 34470 59436 34522
rect 59380 34468 59436 34470
rect 78492 34522 78548 34524
rect 78492 34470 78494 34522
rect 78494 34470 78546 34522
rect 78546 34470 78548 34522
rect 78492 34468 78548 34470
rect 78596 34522 78652 34524
rect 78596 34470 78598 34522
rect 78598 34470 78650 34522
rect 78650 34470 78652 34522
rect 78596 34468 78652 34470
rect 78700 34522 78756 34524
rect 78700 34470 78702 34522
rect 78702 34470 78754 34522
rect 78754 34470 78756 34522
rect 78700 34468 78756 34470
rect 10872 33738 10928 33740
rect 10872 33686 10874 33738
rect 10874 33686 10926 33738
rect 10926 33686 10928 33738
rect 10872 33684 10928 33686
rect 10976 33738 11032 33740
rect 10976 33686 10978 33738
rect 10978 33686 11030 33738
rect 11030 33686 11032 33738
rect 10976 33684 11032 33686
rect 11080 33738 11136 33740
rect 11080 33686 11082 33738
rect 11082 33686 11134 33738
rect 11134 33686 11136 33738
rect 11080 33684 11136 33686
rect 30192 33738 30248 33740
rect 30192 33686 30194 33738
rect 30194 33686 30246 33738
rect 30246 33686 30248 33738
rect 30192 33684 30248 33686
rect 30296 33738 30352 33740
rect 30296 33686 30298 33738
rect 30298 33686 30350 33738
rect 30350 33686 30352 33738
rect 30296 33684 30352 33686
rect 30400 33738 30456 33740
rect 30400 33686 30402 33738
rect 30402 33686 30454 33738
rect 30454 33686 30456 33738
rect 30400 33684 30456 33686
rect 49512 33738 49568 33740
rect 49512 33686 49514 33738
rect 49514 33686 49566 33738
rect 49566 33686 49568 33738
rect 49512 33684 49568 33686
rect 49616 33738 49672 33740
rect 49616 33686 49618 33738
rect 49618 33686 49670 33738
rect 49670 33686 49672 33738
rect 49616 33684 49672 33686
rect 49720 33738 49776 33740
rect 49720 33686 49722 33738
rect 49722 33686 49774 33738
rect 49774 33686 49776 33738
rect 49720 33684 49776 33686
rect 68832 33738 68888 33740
rect 68832 33686 68834 33738
rect 68834 33686 68886 33738
rect 68886 33686 68888 33738
rect 68832 33684 68888 33686
rect 68936 33738 68992 33740
rect 68936 33686 68938 33738
rect 68938 33686 68990 33738
rect 68990 33686 68992 33738
rect 68936 33684 68992 33686
rect 69040 33738 69096 33740
rect 69040 33686 69042 33738
rect 69042 33686 69094 33738
rect 69094 33686 69096 33738
rect 69040 33684 69096 33686
rect 20532 32954 20588 32956
rect 20532 32902 20534 32954
rect 20534 32902 20586 32954
rect 20586 32902 20588 32954
rect 20532 32900 20588 32902
rect 20636 32954 20692 32956
rect 20636 32902 20638 32954
rect 20638 32902 20690 32954
rect 20690 32902 20692 32954
rect 20636 32900 20692 32902
rect 20740 32954 20796 32956
rect 20740 32902 20742 32954
rect 20742 32902 20794 32954
rect 20794 32902 20796 32954
rect 20740 32900 20796 32902
rect 39852 32954 39908 32956
rect 39852 32902 39854 32954
rect 39854 32902 39906 32954
rect 39906 32902 39908 32954
rect 39852 32900 39908 32902
rect 39956 32954 40012 32956
rect 39956 32902 39958 32954
rect 39958 32902 40010 32954
rect 40010 32902 40012 32954
rect 39956 32900 40012 32902
rect 40060 32954 40116 32956
rect 40060 32902 40062 32954
rect 40062 32902 40114 32954
rect 40114 32902 40116 32954
rect 40060 32900 40116 32902
rect 59172 32954 59228 32956
rect 59172 32902 59174 32954
rect 59174 32902 59226 32954
rect 59226 32902 59228 32954
rect 59172 32900 59228 32902
rect 59276 32954 59332 32956
rect 59276 32902 59278 32954
rect 59278 32902 59330 32954
rect 59330 32902 59332 32954
rect 59276 32900 59332 32902
rect 59380 32954 59436 32956
rect 59380 32902 59382 32954
rect 59382 32902 59434 32954
rect 59434 32902 59436 32954
rect 59380 32900 59436 32902
rect 78492 32954 78548 32956
rect 78492 32902 78494 32954
rect 78494 32902 78546 32954
rect 78546 32902 78548 32954
rect 78492 32900 78548 32902
rect 78596 32954 78652 32956
rect 78596 32902 78598 32954
rect 78598 32902 78650 32954
rect 78650 32902 78652 32954
rect 78596 32900 78652 32902
rect 78700 32954 78756 32956
rect 78700 32902 78702 32954
rect 78702 32902 78754 32954
rect 78754 32902 78756 32954
rect 78700 32900 78756 32902
rect 10872 32170 10928 32172
rect 10872 32118 10874 32170
rect 10874 32118 10926 32170
rect 10926 32118 10928 32170
rect 10872 32116 10928 32118
rect 10976 32170 11032 32172
rect 10976 32118 10978 32170
rect 10978 32118 11030 32170
rect 11030 32118 11032 32170
rect 10976 32116 11032 32118
rect 11080 32170 11136 32172
rect 11080 32118 11082 32170
rect 11082 32118 11134 32170
rect 11134 32118 11136 32170
rect 11080 32116 11136 32118
rect 30192 32170 30248 32172
rect 30192 32118 30194 32170
rect 30194 32118 30246 32170
rect 30246 32118 30248 32170
rect 30192 32116 30248 32118
rect 30296 32170 30352 32172
rect 30296 32118 30298 32170
rect 30298 32118 30350 32170
rect 30350 32118 30352 32170
rect 30296 32116 30352 32118
rect 30400 32170 30456 32172
rect 30400 32118 30402 32170
rect 30402 32118 30454 32170
rect 30454 32118 30456 32170
rect 30400 32116 30456 32118
rect 49512 32170 49568 32172
rect 49512 32118 49514 32170
rect 49514 32118 49566 32170
rect 49566 32118 49568 32170
rect 49512 32116 49568 32118
rect 49616 32170 49672 32172
rect 49616 32118 49618 32170
rect 49618 32118 49670 32170
rect 49670 32118 49672 32170
rect 49616 32116 49672 32118
rect 49720 32170 49776 32172
rect 49720 32118 49722 32170
rect 49722 32118 49774 32170
rect 49774 32118 49776 32170
rect 49720 32116 49776 32118
rect 68832 32170 68888 32172
rect 68832 32118 68834 32170
rect 68834 32118 68886 32170
rect 68886 32118 68888 32170
rect 68832 32116 68888 32118
rect 68936 32170 68992 32172
rect 68936 32118 68938 32170
rect 68938 32118 68990 32170
rect 68990 32118 68992 32170
rect 68936 32116 68992 32118
rect 69040 32170 69096 32172
rect 69040 32118 69042 32170
rect 69042 32118 69094 32170
rect 69094 32118 69096 32170
rect 69040 32116 69096 32118
rect 20532 31386 20588 31388
rect 20532 31334 20534 31386
rect 20534 31334 20586 31386
rect 20586 31334 20588 31386
rect 20532 31332 20588 31334
rect 20636 31386 20692 31388
rect 20636 31334 20638 31386
rect 20638 31334 20690 31386
rect 20690 31334 20692 31386
rect 20636 31332 20692 31334
rect 20740 31386 20796 31388
rect 20740 31334 20742 31386
rect 20742 31334 20794 31386
rect 20794 31334 20796 31386
rect 20740 31332 20796 31334
rect 39852 31386 39908 31388
rect 39852 31334 39854 31386
rect 39854 31334 39906 31386
rect 39906 31334 39908 31386
rect 39852 31332 39908 31334
rect 39956 31386 40012 31388
rect 39956 31334 39958 31386
rect 39958 31334 40010 31386
rect 40010 31334 40012 31386
rect 39956 31332 40012 31334
rect 40060 31386 40116 31388
rect 40060 31334 40062 31386
rect 40062 31334 40114 31386
rect 40114 31334 40116 31386
rect 40060 31332 40116 31334
rect 59172 31386 59228 31388
rect 59172 31334 59174 31386
rect 59174 31334 59226 31386
rect 59226 31334 59228 31386
rect 59172 31332 59228 31334
rect 59276 31386 59332 31388
rect 59276 31334 59278 31386
rect 59278 31334 59330 31386
rect 59330 31334 59332 31386
rect 59276 31332 59332 31334
rect 59380 31386 59436 31388
rect 59380 31334 59382 31386
rect 59382 31334 59434 31386
rect 59434 31334 59436 31386
rect 59380 31332 59436 31334
rect 78492 31386 78548 31388
rect 78492 31334 78494 31386
rect 78494 31334 78546 31386
rect 78546 31334 78548 31386
rect 78492 31332 78548 31334
rect 78596 31386 78652 31388
rect 78596 31334 78598 31386
rect 78598 31334 78650 31386
rect 78650 31334 78652 31386
rect 78596 31332 78652 31334
rect 78700 31386 78756 31388
rect 78700 31334 78702 31386
rect 78702 31334 78754 31386
rect 78754 31334 78756 31386
rect 78700 31332 78756 31334
rect 10872 30602 10928 30604
rect 10872 30550 10874 30602
rect 10874 30550 10926 30602
rect 10926 30550 10928 30602
rect 10872 30548 10928 30550
rect 10976 30602 11032 30604
rect 10976 30550 10978 30602
rect 10978 30550 11030 30602
rect 11030 30550 11032 30602
rect 10976 30548 11032 30550
rect 11080 30602 11136 30604
rect 11080 30550 11082 30602
rect 11082 30550 11134 30602
rect 11134 30550 11136 30602
rect 11080 30548 11136 30550
rect 30192 30602 30248 30604
rect 30192 30550 30194 30602
rect 30194 30550 30246 30602
rect 30246 30550 30248 30602
rect 30192 30548 30248 30550
rect 30296 30602 30352 30604
rect 30296 30550 30298 30602
rect 30298 30550 30350 30602
rect 30350 30550 30352 30602
rect 30296 30548 30352 30550
rect 30400 30602 30456 30604
rect 30400 30550 30402 30602
rect 30402 30550 30454 30602
rect 30454 30550 30456 30602
rect 30400 30548 30456 30550
rect 49512 30602 49568 30604
rect 49512 30550 49514 30602
rect 49514 30550 49566 30602
rect 49566 30550 49568 30602
rect 49512 30548 49568 30550
rect 49616 30602 49672 30604
rect 49616 30550 49618 30602
rect 49618 30550 49670 30602
rect 49670 30550 49672 30602
rect 49616 30548 49672 30550
rect 49720 30602 49776 30604
rect 49720 30550 49722 30602
rect 49722 30550 49774 30602
rect 49774 30550 49776 30602
rect 49720 30548 49776 30550
rect 68832 30602 68888 30604
rect 68832 30550 68834 30602
rect 68834 30550 68886 30602
rect 68886 30550 68888 30602
rect 68832 30548 68888 30550
rect 68936 30602 68992 30604
rect 68936 30550 68938 30602
rect 68938 30550 68990 30602
rect 68990 30550 68992 30602
rect 68936 30548 68992 30550
rect 69040 30602 69096 30604
rect 69040 30550 69042 30602
rect 69042 30550 69094 30602
rect 69094 30550 69096 30602
rect 69040 30548 69096 30550
rect 20532 29818 20588 29820
rect 20532 29766 20534 29818
rect 20534 29766 20586 29818
rect 20586 29766 20588 29818
rect 20532 29764 20588 29766
rect 20636 29818 20692 29820
rect 20636 29766 20638 29818
rect 20638 29766 20690 29818
rect 20690 29766 20692 29818
rect 20636 29764 20692 29766
rect 20740 29818 20796 29820
rect 20740 29766 20742 29818
rect 20742 29766 20794 29818
rect 20794 29766 20796 29818
rect 20740 29764 20796 29766
rect 39852 29818 39908 29820
rect 39852 29766 39854 29818
rect 39854 29766 39906 29818
rect 39906 29766 39908 29818
rect 39852 29764 39908 29766
rect 39956 29818 40012 29820
rect 39956 29766 39958 29818
rect 39958 29766 40010 29818
rect 40010 29766 40012 29818
rect 39956 29764 40012 29766
rect 40060 29818 40116 29820
rect 40060 29766 40062 29818
rect 40062 29766 40114 29818
rect 40114 29766 40116 29818
rect 40060 29764 40116 29766
rect 59172 29818 59228 29820
rect 59172 29766 59174 29818
rect 59174 29766 59226 29818
rect 59226 29766 59228 29818
rect 59172 29764 59228 29766
rect 59276 29818 59332 29820
rect 59276 29766 59278 29818
rect 59278 29766 59330 29818
rect 59330 29766 59332 29818
rect 59276 29764 59332 29766
rect 59380 29818 59436 29820
rect 59380 29766 59382 29818
rect 59382 29766 59434 29818
rect 59434 29766 59436 29818
rect 59380 29764 59436 29766
rect 78492 29818 78548 29820
rect 78492 29766 78494 29818
rect 78494 29766 78546 29818
rect 78546 29766 78548 29818
rect 78492 29764 78548 29766
rect 78596 29818 78652 29820
rect 78596 29766 78598 29818
rect 78598 29766 78650 29818
rect 78650 29766 78652 29818
rect 78596 29764 78652 29766
rect 78700 29818 78756 29820
rect 78700 29766 78702 29818
rect 78702 29766 78754 29818
rect 78754 29766 78756 29818
rect 78700 29764 78756 29766
rect 10872 29034 10928 29036
rect 10872 28982 10874 29034
rect 10874 28982 10926 29034
rect 10926 28982 10928 29034
rect 10872 28980 10928 28982
rect 10976 29034 11032 29036
rect 10976 28982 10978 29034
rect 10978 28982 11030 29034
rect 11030 28982 11032 29034
rect 10976 28980 11032 28982
rect 11080 29034 11136 29036
rect 11080 28982 11082 29034
rect 11082 28982 11134 29034
rect 11134 28982 11136 29034
rect 11080 28980 11136 28982
rect 30192 29034 30248 29036
rect 30192 28982 30194 29034
rect 30194 28982 30246 29034
rect 30246 28982 30248 29034
rect 30192 28980 30248 28982
rect 30296 29034 30352 29036
rect 30296 28982 30298 29034
rect 30298 28982 30350 29034
rect 30350 28982 30352 29034
rect 30296 28980 30352 28982
rect 30400 29034 30456 29036
rect 30400 28982 30402 29034
rect 30402 28982 30454 29034
rect 30454 28982 30456 29034
rect 30400 28980 30456 28982
rect 49512 29034 49568 29036
rect 49512 28982 49514 29034
rect 49514 28982 49566 29034
rect 49566 28982 49568 29034
rect 49512 28980 49568 28982
rect 49616 29034 49672 29036
rect 49616 28982 49618 29034
rect 49618 28982 49670 29034
rect 49670 28982 49672 29034
rect 49616 28980 49672 28982
rect 49720 29034 49776 29036
rect 49720 28982 49722 29034
rect 49722 28982 49774 29034
rect 49774 28982 49776 29034
rect 49720 28980 49776 28982
rect 68832 29034 68888 29036
rect 68832 28982 68834 29034
rect 68834 28982 68886 29034
rect 68886 28982 68888 29034
rect 68832 28980 68888 28982
rect 68936 29034 68992 29036
rect 68936 28982 68938 29034
rect 68938 28982 68990 29034
rect 68990 28982 68992 29034
rect 68936 28980 68992 28982
rect 69040 29034 69096 29036
rect 69040 28982 69042 29034
rect 69042 28982 69094 29034
rect 69094 28982 69096 29034
rect 69040 28980 69096 28982
rect 20532 28250 20588 28252
rect 20532 28198 20534 28250
rect 20534 28198 20586 28250
rect 20586 28198 20588 28250
rect 20532 28196 20588 28198
rect 20636 28250 20692 28252
rect 20636 28198 20638 28250
rect 20638 28198 20690 28250
rect 20690 28198 20692 28250
rect 20636 28196 20692 28198
rect 20740 28250 20796 28252
rect 20740 28198 20742 28250
rect 20742 28198 20794 28250
rect 20794 28198 20796 28250
rect 20740 28196 20796 28198
rect 39852 28250 39908 28252
rect 39852 28198 39854 28250
rect 39854 28198 39906 28250
rect 39906 28198 39908 28250
rect 39852 28196 39908 28198
rect 39956 28250 40012 28252
rect 39956 28198 39958 28250
rect 39958 28198 40010 28250
rect 40010 28198 40012 28250
rect 39956 28196 40012 28198
rect 40060 28250 40116 28252
rect 40060 28198 40062 28250
rect 40062 28198 40114 28250
rect 40114 28198 40116 28250
rect 40060 28196 40116 28198
rect 59172 28250 59228 28252
rect 59172 28198 59174 28250
rect 59174 28198 59226 28250
rect 59226 28198 59228 28250
rect 59172 28196 59228 28198
rect 59276 28250 59332 28252
rect 59276 28198 59278 28250
rect 59278 28198 59330 28250
rect 59330 28198 59332 28250
rect 59276 28196 59332 28198
rect 59380 28250 59436 28252
rect 59380 28198 59382 28250
rect 59382 28198 59434 28250
rect 59434 28198 59436 28250
rect 59380 28196 59436 28198
rect 78492 28250 78548 28252
rect 78492 28198 78494 28250
rect 78494 28198 78546 28250
rect 78546 28198 78548 28250
rect 78492 28196 78548 28198
rect 78596 28250 78652 28252
rect 78596 28198 78598 28250
rect 78598 28198 78650 28250
rect 78650 28198 78652 28250
rect 78596 28196 78652 28198
rect 78700 28250 78756 28252
rect 78700 28198 78702 28250
rect 78702 28198 78754 28250
rect 78754 28198 78756 28250
rect 78700 28196 78756 28198
rect 10872 27466 10928 27468
rect 10872 27414 10874 27466
rect 10874 27414 10926 27466
rect 10926 27414 10928 27466
rect 10872 27412 10928 27414
rect 10976 27466 11032 27468
rect 10976 27414 10978 27466
rect 10978 27414 11030 27466
rect 11030 27414 11032 27466
rect 10976 27412 11032 27414
rect 11080 27466 11136 27468
rect 11080 27414 11082 27466
rect 11082 27414 11134 27466
rect 11134 27414 11136 27466
rect 11080 27412 11136 27414
rect 30192 27466 30248 27468
rect 30192 27414 30194 27466
rect 30194 27414 30246 27466
rect 30246 27414 30248 27466
rect 30192 27412 30248 27414
rect 30296 27466 30352 27468
rect 30296 27414 30298 27466
rect 30298 27414 30350 27466
rect 30350 27414 30352 27466
rect 30296 27412 30352 27414
rect 30400 27466 30456 27468
rect 30400 27414 30402 27466
rect 30402 27414 30454 27466
rect 30454 27414 30456 27466
rect 30400 27412 30456 27414
rect 49512 27466 49568 27468
rect 49512 27414 49514 27466
rect 49514 27414 49566 27466
rect 49566 27414 49568 27466
rect 49512 27412 49568 27414
rect 49616 27466 49672 27468
rect 49616 27414 49618 27466
rect 49618 27414 49670 27466
rect 49670 27414 49672 27466
rect 49616 27412 49672 27414
rect 49720 27466 49776 27468
rect 49720 27414 49722 27466
rect 49722 27414 49774 27466
rect 49774 27414 49776 27466
rect 49720 27412 49776 27414
rect 68832 27466 68888 27468
rect 68832 27414 68834 27466
rect 68834 27414 68886 27466
rect 68886 27414 68888 27466
rect 68832 27412 68888 27414
rect 68936 27466 68992 27468
rect 68936 27414 68938 27466
rect 68938 27414 68990 27466
rect 68990 27414 68992 27466
rect 68936 27412 68992 27414
rect 69040 27466 69096 27468
rect 69040 27414 69042 27466
rect 69042 27414 69094 27466
rect 69094 27414 69096 27466
rect 69040 27412 69096 27414
rect 20532 26682 20588 26684
rect 20532 26630 20534 26682
rect 20534 26630 20586 26682
rect 20586 26630 20588 26682
rect 20532 26628 20588 26630
rect 20636 26682 20692 26684
rect 20636 26630 20638 26682
rect 20638 26630 20690 26682
rect 20690 26630 20692 26682
rect 20636 26628 20692 26630
rect 20740 26682 20796 26684
rect 20740 26630 20742 26682
rect 20742 26630 20794 26682
rect 20794 26630 20796 26682
rect 20740 26628 20796 26630
rect 39852 26682 39908 26684
rect 39852 26630 39854 26682
rect 39854 26630 39906 26682
rect 39906 26630 39908 26682
rect 39852 26628 39908 26630
rect 39956 26682 40012 26684
rect 39956 26630 39958 26682
rect 39958 26630 40010 26682
rect 40010 26630 40012 26682
rect 39956 26628 40012 26630
rect 40060 26682 40116 26684
rect 40060 26630 40062 26682
rect 40062 26630 40114 26682
rect 40114 26630 40116 26682
rect 40060 26628 40116 26630
rect 59172 26682 59228 26684
rect 59172 26630 59174 26682
rect 59174 26630 59226 26682
rect 59226 26630 59228 26682
rect 59172 26628 59228 26630
rect 59276 26682 59332 26684
rect 59276 26630 59278 26682
rect 59278 26630 59330 26682
rect 59330 26630 59332 26682
rect 59276 26628 59332 26630
rect 59380 26682 59436 26684
rect 59380 26630 59382 26682
rect 59382 26630 59434 26682
rect 59434 26630 59436 26682
rect 59380 26628 59436 26630
rect 78492 26682 78548 26684
rect 78492 26630 78494 26682
rect 78494 26630 78546 26682
rect 78546 26630 78548 26682
rect 78492 26628 78548 26630
rect 78596 26682 78652 26684
rect 78596 26630 78598 26682
rect 78598 26630 78650 26682
rect 78650 26630 78652 26682
rect 78596 26628 78652 26630
rect 78700 26682 78756 26684
rect 78700 26630 78702 26682
rect 78702 26630 78754 26682
rect 78754 26630 78756 26682
rect 78700 26628 78756 26630
rect 10872 25898 10928 25900
rect 10872 25846 10874 25898
rect 10874 25846 10926 25898
rect 10926 25846 10928 25898
rect 10872 25844 10928 25846
rect 10976 25898 11032 25900
rect 10976 25846 10978 25898
rect 10978 25846 11030 25898
rect 11030 25846 11032 25898
rect 10976 25844 11032 25846
rect 11080 25898 11136 25900
rect 11080 25846 11082 25898
rect 11082 25846 11134 25898
rect 11134 25846 11136 25898
rect 11080 25844 11136 25846
rect 30192 25898 30248 25900
rect 30192 25846 30194 25898
rect 30194 25846 30246 25898
rect 30246 25846 30248 25898
rect 30192 25844 30248 25846
rect 30296 25898 30352 25900
rect 30296 25846 30298 25898
rect 30298 25846 30350 25898
rect 30350 25846 30352 25898
rect 30296 25844 30352 25846
rect 30400 25898 30456 25900
rect 30400 25846 30402 25898
rect 30402 25846 30454 25898
rect 30454 25846 30456 25898
rect 30400 25844 30456 25846
rect 49512 25898 49568 25900
rect 49512 25846 49514 25898
rect 49514 25846 49566 25898
rect 49566 25846 49568 25898
rect 49512 25844 49568 25846
rect 49616 25898 49672 25900
rect 49616 25846 49618 25898
rect 49618 25846 49670 25898
rect 49670 25846 49672 25898
rect 49616 25844 49672 25846
rect 49720 25898 49776 25900
rect 49720 25846 49722 25898
rect 49722 25846 49774 25898
rect 49774 25846 49776 25898
rect 49720 25844 49776 25846
rect 68832 25898 68888 25900
rect 68832 25846 68834 25898
rect 68834 25846 68886 25898
rect 68886 25846 68888 25898
rect 68832 25844 68888 25846
rect 68936 25898 68992 25900
rect 68936 25846 68938 25898
rect 68938 25846 68990 25898
rect 68990 25846 68992 25898
rect 68936 25844 68992 25846
rect 69040 25898 69096 25900
rect 69040 25846 69042 25898
rect 69042 25846 69094 25898
rect 69094 25846 69096 25898
rect 69040 25844 69096 25846
rect 20532 25114 20588 25116
rect 20532 25062 20534 25114
rect 20534 25062 20586 25114
rect 20586 25062 20588 25114
rect 20532 25060 20588 25062
rect 20636 25114 20692 25116
rect 20636 25062 20638 25114
rect 20638 25062 20690 25114
rect 20690 25062 20692 25114
rect 20636 25060 20692 25062
rect 20740 25114 20796 25116
rect 20740 25062 20742 25114
rect 20742 25062 20794 25114
rect 20794 25062 20796 25114
rect 20740 25060 20796 25062
rect 39852 25114 39908 25116
rect 39852 25062 39854 25114
rect 39854 25062 39906 25114
rect 39906 25062 39908 25114
rect 39852 25060 39908 25062
rect 39956 25114 40012 25116
rect 39956 25062 39958 25114
rect 39958 25062 40010 25114
rect 40010 25062 40012 25114
rect 39956 25060 40012 25062
rect 40060 25114 40116 25116
rect 40060 25062 40062 25114
rect 40062 25062 40114 25114
rect 40114 25062 40116 25114
rect 40060 25060 40116 25062
rect 59172 25114 59228 25116
rect 59172 25062 59174 25114
rect 59174 25062 59226 25114
rect 59226 25062 59228 25114
rect 59172 25060 59228 25062
rect 59276 25114 59332 25116
rect 59276 25062 59278 25114
rect 59278 25062 59330 25114
rect 59330 25062 59332 25114
rect 59276 25060 59332 25062
rect 59380 25114 59436 25116
rect 59380 25062 59382 25114
rect 59382 25062 59434 25114
rect 59434 25062 59436 25114
rect 59380 25060 59436 25062
rect 78492 25114 78548 25116
rect 78492 25062 78494 25114
rect 78494 25062 78546 25114
rect 78546 25062 78548 25114
rect 78492 25060 78548 25062
rect 78596 25114 78652 25116
rect 78596 25062 78598 25114
rect 78598 25062 78650 25114
rect 78650 25062 78652 25114
rect 78596 25060 78652 25062
rect 78700 25114 78756 25116
rect 78700 25062 78702 25114
rect 78702 25062 78754 25114
rect 78754 25062 78756 25114
rect 78700 25060 78756 25062
rect 10872 24330 10928 24332
rect 10872 24278 10874 24330
rect 10874 24278 10926 24330
rect 10926 24278 10928 24330
rect 10872 24276 10928 24278
rect 10976 24330 11032 24332
rect 10976 24278 10978 24330
rect 10978 24278 11030 24330
rect 11030 24278 11032 24330
rect 10976 24276 11032 24278
rect 11080 24330 11136 24332
rect 11080 24278 11082 24330
rect 11082 24278 11134 24330
rect 11134 24278 11136 24330
rect 11080 24276 11136 24278
rect 30192 24330 30248 24332
rect 30192 24278 30194 24330
rect 30194 24278 30246 24330
rect 30246 24278 30248 24330
rect 30192 24276 30248 24278
rect 30296 24330 30352 24332
rect 30296 24278 30298 24330
rect 30298 24278 30350 24330
rect 30350 24278 30352 24330
rect 30296 24276 30352 24278
rect 30400 24330 30456 24332
rect 30400 24278 30402 24330
rect 30402 24278 30454 24330
rect 30454 24278 30456 24330
rect 30400 24276 30456 24278
rect 49512 24330 49568 24332
rect 49512 24278 49514 24330
rect 49514 24278 49566 24330
rect 49566 24278 49568 24330
rect 49512 24276 49568 24278
rect 49616 24330 49672 24332
rect 49616 24278 49618 24330
rect 49618 24278 49670 24330
rect 49670 24278 49672 24330
rect 49616 24276 49672 24278
rect 49720 24330 49776 24332
rect 49720 24278 49722 24330
rect 49722 24278 49774 24330
rect 49774 24278 49776 24330
rect 49720 24276 49776 24278
rect 68832 24330 68888 24332
rect 68832 24278 68834 24330
rect 68834 24278 68886 24330
rect 68886 24278 68888 24330
rect 68832 24276 68888 24278
rect 68936 24330 68992 24332
rect 68936 24278 68938 24330
rect 68938 24278 68990 24330
rect 68990 24278 68992 24330
rect 68936 24276 68992 24278
rect 69040 24330 69096 24332
rect 69040 24278 69042 24330
rect 69042 24278 69094 24330
rect 69094 24278 69096 24330
rect 69040 24276 69096 24278
rect 20532 23546 20588 23548
rect 20532 23494 20534 23546
rect 20534 23494 20586 23546
rect 20586 23494 20588 23546
rect 20532 23492 20588 23494
rect 20636 23546 20692 23548
rect 20636 23494 20638 23546
rect 20638 23494 20690 23546
rect 20690 23494 20692 23546
rect 20636 23492 20692 23494
rect 20740 23546 20796 23548
rect 20740 23494 20742 23546
rect 20742 23494 20794 23546
rect 20794 23494 20796 23546
rect 20740 23492 20796 23494
rect 39852 23546 39908 23548
rect 39852 23494 39854 23546
rect 39854 23494 39906 23546
rect 39906 23494 39908 23546
rect 39852 23492 39908 23494
rect 39956 23546 40012 23548
rect 39956 23494 39958 23546
rect 39958 23494 40010 23546
rect 40010 23494 40012 23546
rect 39956 23492 40012 23494
rect 40060 23546 40116 23548
rect 40060 23494 40062 23546
rect 40062 23494 40114 23546
rect 40114 23494 40116 23546
rect 40060 23492 40116 23494
rect 59172 23546 59228 23548
rect 59172 23494 59174 23546
rect 59174 23494 59226 23546
rect 59226 23494 59228 23546
rect 59172 23492 59228 23494
rect 59276 23546 59332 23548
rect 59276 23494 59278 23546
rect 59278 23494 59330 23546
rect 59330 23494 59332 23546
rect 59276 23492 59332 23494
rect 59380 23546 59436 23548
rect 59380 23494 59382 23546
rect 59382 23494 59434 23546
rect 59434 23494 59436 23546
rect 59380 23492 59436 23494
rect 78492 23546 78548 23548
rect 78492 23494 78494 23546
rect 78494 23494 78546 23546
rect 78546 23494 78548 23546
rect 78492 23492 78548 23494
rect 78596 23546 78652 23548
rect 78596 23494 78598 23546
rect 78598 23494 78650 23546
rect 78650 23494 78652 23546
rect 78596 23492 78652 23494
rect 78700 23546 78756 23548
rect 78700 23494 78702 23546
rect 78702 23494 78754 23546
rect 78754 23494 78756 23546
rect 78700 23492 78756 23494
rect 10872 22762 10928 22764
rect 10872 22710 10874 22762
rect 10874 22710 10926 22762
rect 10926 22710 10928 22762
rect 10872 22708 10928 22710
rect 10976 22762 11032 22764
rect 10976 22710 10978 22762
rect 10978 22710 11030 22762
rect 11030 22710 11032 22762
rect 10976 22708 11032 22710
rect 11080 22762 11136 22764
rect 11080 22710 11082 22762
rect 11082 22710 11134 22762
rect 11134 22710 11136 22762
rect 11080 22708 11136 22710
rect 30192 22762 30248 22764
rect 30192 22710 30194 22762
rect 30194 22710 30246 22762
rect 30246 22710 30248 22762
rect 30192 22708 30248 22710
rect 30296 22762 30352 22764
rect 30296 22710 30298 22762
rect 30298 22710 30350 22762
rect 30350 22710 30352 22762
rect 30296 22708 30352 22710
rect 30400 22762 30456 22764
rect 30400 22710 30402 22762
rect 30402 22710 30454 22762
rect 30454 22710 30456 22762
rect 30400 22708 30456 22710
rect 49512 22762 49568 22764
rect 49512 22710 49514 22762
rect 49514 22710 49566 22762
rect 49566 22710 49568 22762
rect 49512 22708 49568 22710
rect 49616 22762 49672 22764
rect 49616 22710 49618 22762
rect 49618 22710 49670 22762
rect 49670 22710 49672 22762
rect 49616 22708 49672 22710
rect 49720 22762 49776 22764
rect 49720 22710 49722 22762
rect 49722 22710 49774 22762
rect 49774 22710 49776 22762
rect 49720 22708 49776 22710
rect 68832 22762 68888 22764
rect 68832 22710 68834 22762
rect 68834 22710 68886 22762
rect 68886 22710 68888 22762
rect 68832 22708 68888 22710
rect 68936 22762 68992 22764
rect 68936 22710 68938 22762
rect 68938 22710 68990 22762
rect 68990 22710 68992 22762
rect 68936 22708 68992 22710
rect 69040 22762 69096 22764
rect 69040 22710 69042 22762
rect 69042 22710 69094 22762
rect 69094 22710 69096 22762
rect 69040 22708 69096 22710
rect 20532 21978 20588 21980
rect 20532 21926 20534 21978
rect 20534 21926 20586 21978
rect 20586 21926 20588 21978
rect 20532 21924 20588 21926
rect 20636 21978 20692 21980
rect 20636 21926 20638 21978
rect 20638 21926 20690 21978
rect 20690 21926 20692 21978
rect 20636 21924 20692 21926
rect 20740 21978 20796 21980
rect 20740 21926 20742 21978
rect 20742 21926 20794 21978
rect 20794 21926 20796 21978
rect 20740 21924 20796 21926
rect 39852 21978 39908 21980
rect 39852 21926 39854 21978
rect 39854 21926 39906 21978
rect 39906 21926 39908 21978
rect 39852 21924 39908 21926
rect 39956 21978 40012 21980
rect 39956 21926 39958 21978
rect 39958 21926 40010 21978
rect 40010 21926 40012 21978
rect 39956 21924 40012 21926
rect 40060 21978 40116 21980
rect 40060 21926 40062 21978
rect 40062 21926 40114 21978
rect 40114 21926 40116 21978
rect 40060 21924 40116 21926
rect 59172 21978 59228 21980
rect 59172 21926 59174 21978
rect 59174 21926 59226 21978
rect 59226 21926 59228 21978
rect 59172 21924 59228 21926
rect 59276 21978 59332 21980
rect 59276 21926 59278 21978
rect 59278 21926 59330 21978
rect 59330 21926 59332 21978
rect 59276 21924 59332 21926
rect 59380 21978 59436 21980
rect 59380 21926 59382 21978
rect 59382 21926 59434 21978
rect 59434 21926 59436 21978
rect 59380 21924 59436 21926
rect 78492 21978 78548 21980
rect 78492 21926 78494 21978
rect 78494 21926 78546 21978
rect 78546 21926 78548 21978
rect 78492 21924 78548 21926
rect 78596 21978 78652 21980
rect 78596 21926 78598 21978
rect 78598 21926 78650 21978
rect 78650 21926 78652 21978
rect 78596 21924 78652 21926
rect 78700 21978 78756 21980
rect 78700 21926 78702 21978
rect 78702 21926 78754 21978
rect 78754 21926 78756 21978
rect 78700 21924 78756 21926
rect 10872 21194 10928 21196
rect 10872 21142 10874 21194
rect 10874 21142 10926 21194
rect 10926 21142 10928 21194
rect 10872 21140 10928 21142
rect 10976 21194 11032 21196
rect 10976 21142 10978 21194
rect 10978 21142 11030 21194
rect 11030 21142 11032 21194
rect 10976 21140 11032 21142
rect 11080 21194 11136 21196
rect 11080 21142 11082 21194
rect 11082 21142 11134 21194
rect 11134 21142 11136 21194
rect 11080 21140 11136 21142
rect 30192 21194 30248 21196
rect 30192 21142 30194 21194
rect 30194 21142 30246 21194
rect 30246 21142 30248 21194
rect 30192 21140 30248 21142
rect 30296 21194 30352 21196
rect 30296 21142 30298 21194
rect 30298 21142 30350 21194
rect 30350 21142 30352 21194
rect 30296 21140 30352 21142
rect 30400 21194 30456 21196
rect 30400 21142 30402 21194
rect 30402 21142 30454 21194
rect 30454 21142 30456 21194
rect 30400 21140 30456 21142
rect 49512 21194 49568 21196
rect 49512 21142 49514 21194
rect 49514 21142 49566 21194
rect 49566 21142 49568 21194
rect 49512 21140 49568 21142
rect 49616 21194 49672 21196
rect 49616 21142 49618 21194
rect 49618 21142 49670 21194
rect 49670 21142 49672 21194
rect 49616 21140 49672 21142
rect 49720 21194 49776 21196
rect 49720 21142 49722 21194
rect 49722 21142 49774 21194
rect 49774 21142 49776 21194
rect 49720 21140 49776 21142
rect 68832 21194 68888 21196
rect 68832 21142 68834 21194
rect 68834 21142 68886 21194
rect 68886 21142 68888 21194
rect 68832 21140 68888 21142
rect 68936 21194 68992 21196
rect 68936 21142 68938 21194
rect 68938 21142 68990 21194
rect 68990 21142 68992 21194
rect 68936 21140 68992 21142
rect 69040 21194 69096 21196
rect 69040 21142 69042 21194
rect 69042 21142 69094 21194
rect 69094 21142 69096 21194
rect 69040 21140 69096 21142
rect 20532 20410 20588 20412
rect 20532 20358 20534 20410
rect 20534 20358 20586 20410
rect 20586 20358 20588 20410
rect 20532 20356 20588 20358
rect 20636 20410 20692 20412
rect 20636 20358 20638 20410
rect 20638 20358 20690 20410
rect 20690 20358 20692 20410
rect 20636 20356 20692 20358
rect 20740 20410 20796 20412
rect 20740 20358 20742 20410
rect 20742 20358 20794 20410
rect 20794 20358 20796 20410
rect 20740 20356 20796 20358
rect 39852 20410 39908 20412
rect 39852 20358 39854 20410
rect 39854 20358 39906 20410
rect 39906 20358 39908 20410
rect 39852 20356 39908 20358
rect 39956 20410 40012 20412
rect 39956 20358 39958 20410
rect 39958 20358 40010 20410
rect 40010 20358 40012 20410
rect 39956 20356 40012 20358
rect 40060 20410 40116 20412
rect 40060 20358 40062 20410
rect 40062 20358 40114 20410
rect 40114 20358 40116 20410
rect 40060 20356 40116 20358
rect 59172 20410 59228 20412
rect 59172 20358 59174 20410
rect 59174 20358 59226 20410
rect 59226 20358 59228 20410
rect 59172 20356 59228 20358
rect 59276 20410 59332 20412
rect 59276 20358 59278 20410
rect 59278 20358 59330 20410
rect 59330 20358 59332 20410
rect 59276 20356 59332 20358
rect 59380 20410 59436 20412
rect 59380 20358 59382 20410
rect 59382 20358 59434 20410
rect 59434 20358 59436 20410
rect 59380 20356 59436 20358
rect 78492 20410 78548 20412
rect 78492 20358 78494 20410
rect 78494 20358 78546 20410
rect 78546 20358 78548 20410
rect 78492 20356 78548 20358
rect 78596 20410 78652 20412
rect 78596 20358 78598 20410
rect 78598 20358 78650 20410
rect 78650 20358 78652 20410
rect 78596 20356 78652 20358
rect 78700 20410 78756 20412
rect 78700 20358 78702 20410
rect 78702 20358 78754 20410
rect 78754 20358 78756 20410
rect 78700 20356 78756 20358
rect 10872 19626 10928 19628
rect 10872 19574 10874 19626
rect 10874 19574 10926 19626
rect 10926 19574 10928 19626
rect 10872 19572 10928 19574
rect 10976 19626 11032 19628
rect 10976 19574 10978 19626
rect 10978 19574 11030 19626
rect 11030 19574 11032 19626
rect 10976 19572 11032 19574
rect 11080 19626 11136 19628
rect 11080 19574 11082 19626
rect 11082 19574 11134 19626
rect 11134 19574 11136 19626
rect 11080 19572 11136 19574
rect 30192 19626 30248 19628
rect 30192 19574 30194 19626
rect 30194 19574 30246 19626
rect 30246 19574 30248 19626
rect 30192 19572 30248 19574
rect 30296 19626 30352 19628
rect 30296 19574 30298 19626
rect 30298 19574 30350 19626
rect 30350 19574 30352 19626
rect 30296 19572 30352 19574
rect 30400 19626 30456 19628
rect 30400 19574 30402 19626
rect 30402 19574 30454 19626
rect 30454 19574 30456 19626
rect 30400 19572 30456 19574
rect 49512 19626 49568 19628
rect 49512 19574 49514 19626
rect 49514 19574 49566 19626
rect 49566 19574 49568 19626
rect 49512 19572 49568 19574
rect 49616 19626 49672 19628
rect 49616 19574 49618 19626
rect 49618 19574 49670 19626
rect 49670 19574 49672 19626
rect 49616 19572 49672 19574
rect 49720 19626 49776 19628
rect 49720 19574 49722 19626
rect 49722 19574 49774 19626
rect 49774 19574 49776 19626
rect 49720 19572 49776 19574
rect 68832 19626 68888 19628
rect 68832 19574 68834 19626
rect 68834 19574 68886 19626
rect 68886 19574 68888 19626
rect 68832 19572 68888 19574
rect 68936 19626 68992 19628
rect 68936 19574 68938 19626
rect 68938 19574 68990 19626
rect 68990 19574 68992 19626
rect 68936 19572 68992 19574
rect 69040 19626 69096 19628
rect 69040 19574 69042 19626
rect 69042 19574 69094 19626
rect 69094 19574 69096 19626
rect 69040 19572 69096 19574
rect 20532 18842 20588 18844
rect 20532 18790 20534 18842
rect 20534 18790 20586 18842
rect 20586 18790 20588 18842
rect 20532 18788 20588 18790
rect 20636 18842 20692 18844
rect 20636 18790 20638 18842
rect 20638 18790 20690 18842
rect 20690 18790 20692 18842
rect 20636 18788 20692 18790
rect 20740 18842 20796 18844
rect 20740 18790 20742 18842
rect 20742 18790 20794 18842
rect 20794 18790 20796 18842
rect 20740 18788 20796 18790
rect 39852 18842 39908 18844
rect 39852 18790 39854 18842
rect 39854 18790 39906 18842
rect 39906 18790 39908 18842
rect 39852 18788 39908 18790
rect 39956 18842 40012 18844
rect 39956 18790 39958 18842
rect 39958 18790 40010 18842
rect 40010 18790 40012 18842
rect 39956 18788 40012 18790
rect 40060 18842 40116 18844
rect 40060 18790 40062 18842
rect 40062 18790 40114 18842
rect 40114 18790 40116 18842
rect 40060 18788 40116 18790
rect 59172 18842 59228 18844
rect 59172 18790 59174 18842
rect 59174 18790 59226 18842
rect 59226 18790 59228 18842
rect 59172 18788 59228 18790
rect 59276 18842 59332 18844
rect 59276 18790 59278 18842
rect 59278 18790 59330 18842
rect 59330 18790 59332 18842
rect 59276 18788 59332 18790
rect 59380 18842 59436 18844
rect 59380 18790 59382 18842
rect 59382 18790 59434 18842
rect 59434 18790 59436 18842
rect 59380 18788 59436 18790
rect 78492 18842 78548 18844
rect 78492 18790 78494 18842
rect 78494 18790 78546 18842
rect 78546 18790 78548 18842
rect 78492 18788 78548 18790
rect 78596 18842 78652 18844
rect 78596 18790 78598 18842
rect 78598 18790 78650 18842
rect 78650 18790 78652 18842
rect 78596 18788 78652 18790
rect 78700 18842 78756 18844
rect 78700 18790 78702 18842
rect 78702 18790 78754 18842
rect 78754 18790 78756 18842
rect 78700 18788 78756 18790
rect 16716 18508 16772 18564
rect 10872 18058 10928 18060
rect 10872 18006 10874 18058
rect 10874 18006 10926 18058
rect 10926 18006 10928 18058
rect 10872 18004 10928 18006
rect 10976 18058 11032 18060
rect 10976 18006 10978 18058
rect 10978 18006 11030 18058
rect 11030 18006 11032 18058
rect 10976 18004 11032 18006
rect 11080 18058 11136 18060
rect 11080 18006 11082 18058
rect 11082 18006 11134 18058
rect 11134 18006 11136 18058
rect 11080 18004 11136 18006
rect 4844 17388 4900 17444
rect 3836 5516 3892 5572
rect 2604 5068 2660 5124
rect 2268 4338 2324 4340
rect 2268 4286 2270 4338
rect 2270 4286 2322 4338
rect 2322 4286 2324 4338
rect 2268 4284 2324 4286
rect 2492 3724 2548 3780
rect 2268 3554 2324 3556
rect 2268 3502 2270 3554
rect 2270 3502 2322 3554
rect 2322 3502 2324 3554
rect 2268 3500 2324 3502
rect 1932 3442 1988 3444
rect 1932 3390 1934 3442
rect 1934 3390 1986 3442
rect 1986 3390 1988 3442
rect 1932 3388 1988 3390
rect 4732 5404 4788 5460
rect 3388 4844 3444 4900
rect 10872 16490 10928 16492
rect 10872 16438 10874 16490
rect 10874 16438 10926 16490
rect 10926 16438 10928 16490
rect 10872 16436 10928 16438
rect 10976 16490 11032 16492
rect 10976 16438 10978 16490
rect 10978 16438 11030 16490
rect 11030 16438 11032 16490
rect 10976 16436 11032 16438
rect 11080 16490 11136 16492
rect 11080 16438 11082 16490
rect 11082 16438 11134 16490
rect 11134 16438 11136 16490
rect 11080 16436 11136 16438
rect 4956 15260 5012 15316
rect 6412 15148 6468 15204
rect 54572 18508 54628 18564
rect 30192 18058 30248 18060
rect 30192 18006 30194 18058
rect 30194 18006 30246 18058
rect 30246 18006 30248 18058
rect 30192 18004 30248 18006
rect 30296 18058 30352 18060
rect 30296 18006 30298 18058
rect 30298 18006 30350 18058
rect 30350 18006 30352 18058
rect 30296 18004 30352 18006
rect 30400 18058 30456 18060
rect 30400 18006 30402 18058
rect 30402 18006 30454 18058
rect 30454 18006 30456 18058
rect 30400 18004 30456 18006
rect 49512 18058 49568 18060
rect 49512 18006 49514 18058
rect 49514 18006 49566 18058
rect 49566 18006 49568 18058
rect 49512 18004 49568 18006
rect 49616 18058 49672 18060
rect 49616 18006 49618 18058
rect 49618 18006 49670 18058
rect 49670 18006 49672 18058
rect 49616 18004 49672 18006
rect 49720 18058 49776 18060
rect 49720 18006 49722 18058
rect 49722 18006 49774 18058
rect 49774 18006 49776 18058
rect 49720 18004 49776 18006
rect 20532 17274 20588 17276
rect 20532 17222 20534 17274
rect 20534 17222 20586 17274
rect 20586 17222 20588 17274
rect 20532 17220 20588 17222
rect 20636 17274 20692 17276
rect 20636 17222 20638 17274
rect 20638 17222 20690 17274
rect 20690 17222 20692 17274
rect 20636 17220 20692 17222
rect 20740 17274 20796 17276
rect 20740 17222 20742 17274
rect 20742 17222 20794 17274
rect 20794 17222 20796 17274
rect 39852 17274 39908 17276
rect 20740 17220 20796 17222
rect 37772 17164 37828 17220
rect 39852 17222 39854 17274
rect 39854 17222 39906 17274
rect 39906 17222 39908 17274
rect 39852 17220 39908 17222
rect 39956 17274 40012 17276
rect 39956 17222 39958 17274
rect 39958 17222 40010 17274
rect 40010 17222 40012 17274
rect 39956 17220 40012 17222
rect 40060 17274 40116 17276
rect 40060 17222 40062 17274
rect 40062 17222 40114 17274
rect 40114 17222 40116 17274
rect 40060 17220 40116 17222
rect 6076 7586 6132 7588
rect 6076 7534 6078 7586
rect 6078 7534 6130 7586
rect 6130 7534 6132 7586
rect 6076 7532 6132 7534
rect 5068 6860 5124 6916
rect 5852 7308 5908 7364
rect 5068 5682 5124 5684
rect 5068 5630 5070 5682
rect 5070 5630 5122 5682
rect 5122 5630 5124 5682
rect 5068 5628 5124 5630
rect 4620 4844 4676 4900
rect 5628 5292 5684 5348
rect 4284 4396 4340 4452
rect 4844 4060 4900 4116
rect 3276 3836 3332 3892
rect 3500 3836 3556 3892
rect 2940 3612 2996 3668
rect 6076 6188 6132 6244
rect 5964 6076 6020 6132
rect 5852 5180 5908 5236
rect 6300 6690 6356 6692
rect 6300 6638 6302 6690
rect 6302 6638 6354 6690
rect 6354 6638 6356 6690
rect 6300 6636 6356 6638
rect 20188 17052 20244 17108
rect 10872 14922 10928 14924
rect 10872 14870 10874 14922
rect 10874 14870 10926 14922
rect 10926 14870 10928 14922
rect 10872 14868 10928 14870
rect 10976 14922 11032 14924
rect 10976 14870 10978 14922
rect 10978 14870 11030 14922
rect 11030 14870 11032 14922
rect 10976 14868 11032 14870
rect 11080 14922 11136 14924
rect 11080 14870 11082 14922
rect 11082 14870 11134 14922
rect 11134 14870 11136 14922
rect 11080 14868 11136 14870
rect 10444 13692 10500 13748
rect 9548 12908 9604 12964
rect 10108 12962 10164 12964
rect 10108 12910 10110 12962
rect 10110 12910 10162 12962
rect 10162 12910 10164 12962
rect 10108 12908 10164 12910
rect 9772 12348 9828 12404
rect 9548 9996 9604 10052
rect 6748 9436 6804 9492
rect 6524 7362 6580 7364
rect 6524 7310 6526 7362
rect 6526 7310 6578 7362
rect 6578 7310 6580 7362
rect 6524 7308 6580 7310
rect 6524 6748 6580 6804
rect 6636 6636 6692 6692
rect 6188 6076 6244 6132
rect 6188 5234 6244 5236
rect 6188 5182 6190 5234
rect 6190 5182 6242 5234
rect 6242 5182 6244 5234
rect 6188 5180 6244 5182
rect 5740 4956 5796 5012
rect 5628 3948 5684 4004
rect 5628 3612 5684 3668
rect 3388 3500 3444 3556
rect 3612 3554 3668 3556
rect 3612 3502 3614 3554
rect 3614 3502 3666 3554
rect 3666 3502 3668 3554
rect 3612 3500 3668 3502
rect 2940 2492 2996 2548
rect 4508 3388 4564 3444
rect 4060 2604 4116 2660
rect 3164 2380 3220 2436
rect 5852 1036 5908 1092
rect 8540 8316 8596 8372
rect 7084 6524 7140 6580
rect 7084 6300 7140 6356
rect 7196 6188 7252 6244
rect 6860 5628 6916 5684
rect 6412 5122 6468 5124
rect 6412 5070 6414 5122
rect 6414 5070 6466 5122
rect 6466 5070 6468 5122
rect 6412 5068 6468 5070
rect 6524 4844 6580 4900
rect 7084 5628 7140 5684
rect 7084 5292 7140 5348
rect 7756 6690 7812 6692
rect 7756 6638 7758 6690
rect 7758 6638 7810 6690
rect 7810 6638 7812 6690
rect 7756 6636 7812 6638
rect 7644 6188 7700 6244
rect 8652 6300 8708 6356
rect 7756 5404 7812 5460
rect 7308 4508 7364 4564
rect 7420 4956 7476 5012
rect 6972 3500 7028 3556
rect 7196 3388 7252 3444
rect 7868 4226 7924 4228
rect 7868 4174 7870 4226
rect 7870 4174 7922 4226
rect 7922 4174 7924 4226
rect 7868 4172 7924 4174
rect 7756 3388 7812 3444
rect 8316 4284 8372 4340
rect 8876 5964 8932 6020
rect 8988 5906 9044 5908
rect 8988 5854 8990 5906
rect 8990 5854 9042 5906
rect 9042 5854 9044 5906
rect 8988 5852 9044 5854
rect 8764 5628 8820 5684
rect 8988 5628 9044 5684
rect 8764 4844 8820 4900
rect 9996 8764 10052 8820
rect 9884 8258 9940 8260
rect 9884 8206 9886 8258
rect 9886 8206 9938 8258
rect 9938 8206 9940 8258
rect 9884 8204 9940 8206
rect 10872 13354 10928 13356
rect 10872 13302 10874 13354
rect 10874 13302 10926 13354
rect 10926 13302 10928 13354
rect 10872 13300 10928 13302
rect 10976 13354 11032 13356
rect 10976 13302 10978 13354
rect 10978 13302 11030 13354
rect 11030 13302 11032 13354
rect 10976 13300 11032 13302
rect 11080 13354 11136 13356
rect 11080 13302 11082 13354
rect 11082 13302 11134 13354
rect 11134 13302 11136 13354
rect 11080 13300 11136 13302
rect 10872 11786 10928 11788
rect 10872 11734 10874 11786
rect 10874 11734 10926 11786
rect 10926 11734 10928 11786
rect 10872 11732 10928 11734
rect 10976 11786 11032 11788
rect 10976 11734 10978 11786
rect 10978 11734 11030 11786
rect 11030 11734 11032 11786
rect 10976 11732 11032 11734
rect 11080 11786 11136 11788
rect 11080 11734 11082 11786
rect 11082 11734 11134 11786
rect 11134 11734 11136 11786
rect 11080 11732 11136 11734
rect 11676 11788 11732 11844
rect 10872 10218 10928 10220
rect 10872 10166 10874 10218
rect 10874 10166 10926 10218
rect 10926 10166 10928 10218
rect 10872 10164 10928 10166
rect 10976 10218 11032 10220
rect 10976 10166 10978 10218
rect 10978 10166 11030 10218
rect 11030 10166 11032 10218
rect 10976 10164 11032 10166
rect 11080 10218 11136 10220
rect 11080 10166 11082 10218
rect 11082 10166 11134 10218
rect 11134 10166 11136 10218
rect 11080 10164 11136 10166
rect 11452 9660 11508 9716
rect 11564 9548 11620 9604
rect 9212 6524 9268 6580
rect 9436 6748 9492 6804
rect 9324 5516 9380 5572
rect 8876 4172 8932 4228
rect 9324 3948 9380 4004
rect 9212 3836 9268 3892
rect 9548 6300 9604 6356
rect 9660 6412 9716 6468
rect 9772 5628 9828 5684
rect 9884 6524 9940 6580
rect 9548 5180 9604 5236
rect 9996 6188 10052 6244
rect 9884 5122 9940 5124
rect 9884 5070 9886 5122
rect 9886 5070 9938 5122
rect 9938 5070 9940 5122
rect 9884 5068 9940 5070
rect 9772 3724 9828 3780
rect 9884 4060 9940 4116
rect 9660 2940 9716 2996
rect 10332 8204 10388 8260
rect 10444 7644 10500 7700
rect 10872 8650 10928 8652
rect 10872 8598 10874 8650
rect 10874 8598 10926 8650
rect 10926 8598 10928 8650
rect 10872 8596 10928 8598
rect 10976 8650 11032 8652
rect 10976 8598 10978 8650
rect 10978 8598 11030 8650
rect 11030 8598 11032 8650
rect 10976 8596 11032 8598
rect 11080 8650 11136 8652
rect 11080 8598 11082 8650
rect 11082 8598 11134 8650
rect 11134 8598 11136 8650
rect 11080 8596 11136 8598
rect 10872 7082 10928 7084
rect 10872 7030 10874 7082
rect 10874 7030 10926 7082
rect 10926 7030 10928 7082
rect 10872 7028 10928 7030
rect 10976 7082 11032 7084
rect 10976 7030 10978 7082
rect 10978 7030 11030 7082
rect 11030 7030 11032 7082
rect 10976 7028 11032 7030
rect 11080 7082 11136 7084
rect 11080 7030 11082 7082
rect 11082 7030 11134 7082
rect 11134 7030 11136 7082
rect 11080 7028 11136 7030
rect 10332 6018 10388 6020
rect 10332 5966 10334 6018
rect 10334 5966 10386 6018
rect 10386 5966 10388 6018
rect 10332 5964 10388 5966
rect 10556 5628 10612 5684
rect 10872 5514 10928 5516
rect 10872 5462 10874 5514
rect 10874 5462 10926 5514
rect 10926 5462 10928 5514
rect 10872 5460 10928 5462
rect 10976 5514 11032 5516
rect 10976 5462 10978 5514
rect 10978 5462 11030 5514
rect 11030 5462 11032 5514
rect 10976 5460 11032 5462
rect 11080 5514 11136 5516
rect 11080 5462 11082 5514
rect 11082 5462 11134 5514
rect 11134 5462 11136 5514
rect 11080 5460 11136 5462
rect 10892 5292 10948 5348
rect 10668 4562 10724 4564
rect 10668 4510 10670 4562
rect 10670 4510 10722 4562
rect 10722 4510 10724 4562
rect 10668 4508 10724 4510
rect 10872 3946 10928 3948
rect 10872 3894 10874 3946
rect 10874 3894 10926 3946
rect 10926 3894 10928 3946
rect 10872 3892 10928 3894
rect 10976 3946 11032 3948
rect 10976 3894 10978 3946
rect 10978 3894 11030 3946
rect 11030 3894 11032 3946
rect 10976 3892 11032 3894
rect 11080 3946 11136 3948
rect 11080 3894 11082 3946
rect 11082 3894 11134 3946
rect 11134 3894 11136 3946
rect 11080 3892 11136 3894
rect 12124 11228 12180 11284
rect 14924 13468 14980 13524
rect 13244 12908 13300 12964
rect 12908 11788 12964 11844
rect 13132 11228 13188 11284
rect 12348 11116 12404 11172
rect 12236 10444 12292 10500
rect 13692 12178 13748 12180
rect 13692 12126 13694 12178
rect 13694 12126 13746 12178
rect 13746 12126 13748 12178
rect 13692 12124 13748 12126
rect 13580 11170 13636 11172
rect 13580 11118 13582 11170
rect 13582 11118 13634 11170
rect 13634 11118 13636 11170
rect 13580 11116 13636 11118
rect 13244 10108 13300 10164
rect 14700 11282 14756 11284
rect 14700 11230 14702 11282
rect 14702 11230 14754 11282
rect 14754 11230 14756 11282
rect 14700 11228 14756 11230
rect 14476 10668 14532 10724
rect 14028 10498 14084 10500
rect 14028 10446 14030 10498
rect 14030 10446 14082 10498
rect 14082 10446 14084 10498
rect 14028 10444 14084 10446
rect 13580 10220 13636 10276
rect 12124 9042 12180 9044
rect 12124 8990 12126 9042
rect 12126 8990 12178 9042
rect 12178 8990 12180 9042
rect 12124 8988 12180 8990
rect 11788 7644 11844 7700
rect 11452 6300 11508 6356
rect 10108 1148 10164 1204
rect 11564 3666 11620 3668
rect 11564 3614 11566 3666
rect 11566 3614 11618 3666
rect 11618 3614 11620 3666
rect 11564 3612 11620 3614
rect 12460 6860 12516 6916
rect 13356 9660 13412 9716
rect 12908 9602 12964 9604
rect 12908 9550 12910 9602
rect 12910 9550 12962 9602
rect 12962 9550 12964 9602
rect 12908 9548 12964 9550
rect 12908 8876 12964 8932
rect 12684 5740 12740 5796
rect 15260 12124 15316 12180
rect 15148 11282 15204 11284
rect 15148 11230 15150 11282
rect 15150 11230 15202 11282
rect 15202 11230 15204 11282
rect 15148 11228 15204 11230
rect 14028 8988 14084 9044
rect 13580 8428 13636 8484
rect 13804 8146 13860 8148
rect 13804 8094 13806 8146
rect 13806 8094 13858 8146
rect 13858 8094 13860 8146
rect 13804 8092 13860 8094
rect 13468 7644 13524 7700
rect 13132 6524 13188 6580
rect 13692 6578 13748 6580
rect 13692 6526 13694 6578
rect 13694 6526 13746 6578
rect 13746 6526 13748 6578
rect 13692 6524 13748 6526
rect 13132 4396 13188 4452
rect 13132 3554 13188 3556
rect 13132 3502 13134 3554
rect 13134 3502 13186 3554
rect 13186 3502 13188 3554
rect 13132 3500 13188 3502
rect 12796 2492 12852 2548
rect 13468 3330 13524 3332
rect 13468 3278 13470 3330
rect 13470 3278 13522 3330
rect 13522 3278 13524 3330
rect 13468 3276 13524 3278
rect 13916 5964 13972 6020
rect 13916 5740 13972 5796
rect 13692 5292 13748 5348
rect 13692 5122 13748 5124
rect 13692 5070 13694 5122
rect 13694 5070 13746 5122
rect 13746 5070 13748 5122
rect 13692 5068 13748 5070
rect 13804 3276 13860 3332
rect 14588 8034 14644 8036
rect 14588 7982 14590 8034
rect 14590 7982 14642 8034
rect 14642 7982 14644 8034
rect 14588 7980 14644 7982
rect 14364 6972 14420 7028
rect 15820 10668 15876 10724
rect 15260 9996 15316 10052
rect 19292 13916 19348 13972
rect 17948 13132 18004 13188
rect 17500 12178 17556 12180
rect 17500 12126 17502 12178
rect 17502 12126 17554 12178
rect 17554 12126 17556 12178
rect 17500 12124 17556 12126
rect 16492 11228 16548 11284
rect 16380 10498 16436 10500
rect 16380 10446 16382 10498
rect 16382 10446 16434 10498
rect 16434 10446 16436 10498
rect 16380 10444 16436 10446
rect 16268 10108 16324 10164
rect 16156 9714 16212 9716
rect 16156 9662 16158 9714
rect 16158 9662 16210 9714
rect 16210 9662 16212 9714
rect 16156 9660 16212 9662
rect 15372 8204 15428 8260
rect 15260 7980 15316 8036
rect 15036 6972 15092 7028
rect 15260 7420 15316 7476
rect 14700 6690 14756 6692
rect 14700 6638 14702 6690
rect 14702 6638 14754 6690
rect 14754 6638 14756 6690
rect 14700 6636 14756 6638
rect 14476 6412 14532 6468
rect 15820 6188 15876 6244
rect 15932 8146 15988 8148
rect 15932 8094 15934 8146
rect 15934 8094 15986 8146
rect 15986 8094 15988 8146
rect 15932 8092 15988 8094
rect 15708 5964 15764 6020
rect 14924 4396 14980 4452
rect 13804 1372 13860 1428
rect 14364 3388 14420 3444
rect 14812 3442 14868 3444
rect 14812 3390 14814 3442
rect 14814 3390 14866 3442
rect 14866 3390 14868 3442
rect 14812 3388 14868 3390
rect 15708 5292 15764 5348
rect 15484 3724 15540 3780
rect 16044 5852 16100 5908
rect 16156 6300 16212 6356
rect 16380 8092 16436 8148
rect 16940 11564 16996 11620
rect 16828 10444 16884 10500
rect 16604 8146 16660 8148
rect 16604 8094 16606 8146
rect 16606 8094 16658 8146
rect 16658 8094 16660 8146
rect 16604 8092 16660 8094
rect 16604 6748 16660 6804
rect 16828 7308 16884 7364
rect 16716 6412 16772 6468
rect 16828 6300 16884 6356
rect 16716 6076 16772 6132
rect 16156 5628 16212 5684
rect 16044 5068 16100 5124
rect 16604 5234 16660 5236
rect 16604 5182 16606 5234
rect 16606 5182 16658 5234
rect 16658 5182 16660 5234
rect 16604 5180 16660 5182
rect 16156 4956 16212 5012
rect 16044 2828 16100 2884
rect 16380 3612 16436 3668
rect 18284 12684 18340 12740
rect 17500 10498 17556 10500
rect 17500 10446 17502 10498
rect 17502 10446 17554 10498
rect 17554 10446 17556 10498
rect 17500 10444 17556 10446
rect 17500 9660 17556 9716
rect 18172 11228 18228 11284
rect 18844 11170 18900 11172
rect 18844 11118 18846 11170
rect 18846 11118 18898 11170
rect 18898 11118 18900 11170
rect 18844 11116 18900 11118
rect 18284 10444 18340 10500
rect 18172 10108 18228 10164
rect 17500 8258 17556 8260
rect 17500 8206 17502 8258
rect 17502 8206 17554 8258
rect 17554 8206 17556 8258
rect 17500 8204 17556 8206
rect 17388 8092 17444 8148
rect 17724 7698 17780 7700
rect 17724 7646 17726 7698
rect 17726 7646 17778 7698
rect 17778 7646 17780 7698
rect 17724 7644 17780 7646
rect 17164 5404 17220 5460
rect 17276 6748 17332 6804
rect 17388 6300 17444 6356
rect 17500 6188 17556 6244
rect 18172 7420 18228 7476
rect 18732 9996 18788 10052
rect 18844 9266 18900 9268
rect 18844 9214 18846 9266
rect 18846 9214 18898 9266
rect 18898 9214 18900 9266
rect 18844 9212 18900 9214
rect 17388 5906 17444 5908
rect 17388 5854 17390 5906
rect 17390 5854 17442 5906
rect 17442 5854 17444 5906
rect 17388 5852 17444 5854
rect 17724 5628 17780 5684
rect 17612 5516 17668 5572
rect 16940 5122 16996 5124
rect 16940 5070 16942 5122
rect 16942 5070 16994 5122
rect 16994 5070 16996 5122
rect 16940 5068 16996 5070
rect 18060 5068 18116 5124
rect 17836 3836 17892 3892
rect 18844 7362 18900 7364
rect 18844 7310 18846 7362
rect 18846 7310 18898 7362
rect 18898 7310 18900 7362
rect 18844 7308 18900 7310
rect 18508 4956 18564 5012
rect 19628 12236 19684 12292
rect 19852 11394 19908 11396
rect 19852 11342 19854 11394
rect 19854 11342 19906 11394
rect 19906 11342 19908 11394
rect 19852 11340 19908 11342
rect 19852 9436 19908 9492
rect 19516 8146 19572 8148
rect 19516 8094 19518 8146
rect 19518 8094 19570 8146
rect 19570 8094 19572 8146
rect 19516 8092 19572 8094
rect 19516 7420 19572 7476
rect 19292 6748 19348 6804
rect 19180 6076 19236 6132
rect 19292 6300 19348 6356
rect 27580 17052 27636 17108
rect 23772 16828 23828 16884
rect 20532 15706 20588 15708
rect 20532 15654 20534 15706
rect 20534 15654 20586 15706
rect 20586 15654 20588 15706
rect 20532 15652 20588 15654
rect 20636 15706 20692 15708
rect 20636 15654 20638 15706
rect 20638 15654 20690 15706
rect 20690 15654 20692 15706
rect 20636 15652 20692 15654
rect 20740 15706 20796 15708
rect 20740 15654 20742 15706
rect 20742 15654 20794 15706
rect 20794 15654 20796 15706
rect 20740 15652 20796 15654
rect 27356 15820 27412 15876
rect 20532 14138 20588 14140
rect 20532 14086 20534 14138
rect 20534 14086 20586 14138
rect 20586 14086 20588 14138
rect 20532 14084 20588 14086
rect 20636 14138 20692 14140
rect 20636 14086 20638 14138
rect 20638 14086 20690 14138
rect 20690 14086 20692 14138
rect 20636 14084 20692 14086
rect 20740 14138 20796 14140
rect 20740 14086 20742 14138
rect 20742 14086 20794 14138
rect 20794 14086 20796 14138
rect 20740 14084 20796 14086
rect 20860 12738 20916 12740
rect 20860 12686 20862 12738
rect 20862 12686 20914 12738
rect 20914 12686 20916 12738
rect 20860 12684 20916 12686
rect 20532 12570 20588 12572
rect 20532 12518 20534 12570
rect 20534 12518 20586 12570
rect 20586 12518 20588 12570
rect 20532 12516 20588 12518
rect 20636 12570 20692 12572
rect 20636 12518 20638 12570
rect 20638 12518 20690 12570
rect 20690 12518 20692 12570
rect 20636 12516 20692 12518
rect 20740 12570 20796 12572
rect 20740 12518 20742 12570
rect 20742 12518 20794 12570
rect 20794 12518 20796 12570
rect 20740 12516 20796 12518
rect 20300 12290 20356 12292
rect 20300 12238 20302 12290
rect 20302 12238 20354 12290
rect 20354 12238 20356 12290
rect 20300 12236 20356 12238
rect 20412 11282 20468 11284
rect 20412 11230 20414 11282
rect 20414 11230 20466 11282
rect 20466 11230 20468 11282
rect 20412 11228 20468 11230
rect 20532 11002 20588 11004
rect 20532 10950 20534 11002
rect 20534 10950 20586 11002
rect 20586 10950 20588 11002
rect 20532 10948 20588 10950
rect 20636 11002 20692 11004
rect 20636 10950 20638 11002
rect 20638 10950 20690 11002
rect 20690 10950 20692 11002
rect 20636 10948 20692 10950
rect 20740 11002 20796 11004
rect 20740 10950 20742 11002
rect 20742 10950 20794 11002
rect 20794 10950 20796 11002
rect 20740 10948 20796 10950
rect 20300 9996 20356 10052
rect 22540 12684 22596 12740
rect 22652 11788 22708 11844
rect 21756 11452 21812 11508
rect 21420 11340 21476 11396
rect 21308 10108 21364 10164
rect 20972 9996 21028 10052
rect 21420 9996 21476 10052
rect 20860 9602 20916 9604
rect 20860 9550 20862 9602
rect 20862 9550 20914 9602
rect 20914 9550 20916 9602
rect 20860 9548 20916 9550
rect 20532 9434 20588 9436
rect 20532 9382 20534 9434
rect 20534 9382 20586 9434
rect 20586 9382 20588 9434
rect 20532 9380 20588 9382
rect 20636 9434 20692 9436
rect 20636 9382 20638 9434
rect 20638 9382 20690 9434
rect 20690 9382 20692 9434
rect 20636 9380 20692 9382
rect 20740 9434 20796 9436
rect 20740 9382 20742 9434
rect 20742 9382 20794 9434
rect 20794 9382 20796 9434
rect 20740 9380 20796 9382
rect 20188 9212 20244 9268
rect 20076 9100 20132 9156
rect 21532 8876 21588 8932
rect 21644 8316 21700 8372
rect 19852 7644 19908 7700
rect 19628 7308 19684 7364
rect 20532 7866 20588 7868
rect 20532 7814 20534 7866
rect 20534 7814 20586 7866
rect 20586 7814 20588 7866
rect 20532 7812 20588 7814
rect 20636 7866 20692 7868
rect 20636 7814 20638 7866
rect 20638 7814 20690 7866
rect 20690 7814 20692 7866
rect 20636 7812 20692 7814
rect 20740 7866 20796 7868
rect 20740 7814 20742 7866
rect 20742 7814 20794 7866
rect 20794 7814 20796 7866
rect 20740 7812 20796 7814
rect 20076 7308 20132 7364
rect 19628 7084 19684 7140
rect 18396 4508 18452 4564
rect 18172 3724 18228 3780
rect 16940 1036 16996 1092
rect 17948 3612 18004 3668
rect 18172 3500 18228 3556
rect 18396 3388 18452 3444
rect 18620 2716 18676 2772
rect 18956 924 19012 980
rect 20412 6636 20468 6692
rect 20524 6748 20580 6804
rect 21644 7980 21700 8036
rect 21308 7868 21364 7924
rect 19964 5122 20020 5124
rect 19964 5070 19966 5122
rect 19966 5070 20018 5122
rect 20018 5070 20020 5122
rect 19964 5068 20020 5070
rect 19852 4844 19908 4900
rect 20300 1372 20356 1428
rect 20300 1036 20356 1092
rect 20532 6298 20588 6300
rect 20532 6246 20534 6298
rect 20534 6246 20586 6298
rect 20586 6246 20588 6298
rect 20532 6244 20588 6246
rect 20636 6298 20692 6300
rect 20636 6246 20638 6298
rect 20638 6246 20690 6298
rect 20690 6246 20692 6298
rect 20636 6244 20692 6246
rect 20740 6298 20796 6300
rect 20740 6246 20742 6298
rect 20742 6246 20794 6298
rect 20794 6246 20796 6298
rect 20740 6244 20796 6246
rect 20748 5852 20804 5908
rect 21532 7308 21588 7364
rect 22204 11282 22260 11284
rect 22204 11230 22206 11282
rect 22206 11230 22258 11282
rect 22258 11230 22260 11282
rect 22204 11228 22260 11230
rect 21980 10108 22036 10164
rect 21868 9996 21924 10052
rect 21756 7868 21812 7924
rect 21868 8204 21924 8260
rect 21756 7644 21812 7700
rect 21756 6690 21812 6692
rect 21756 6638 21758 6690
rect 21758 6638 21810 6690
rect 21810 6638 21812 6690
rect 21756 6636 21812 6638
rect 22316 11004 22372 11060
rect 22540 11228 22596 11284
rect 22764 11170 22820 11172
rect 22764 11118 22766 11170
rect 22766 11118 22818 11170
rect 22818 11118 22820 11170
rect 22764 11116 22820 11118
rect 22876 10220 22932 10276
rect 22092 8204 22148 8260
rect 21980 6860 22036 6916
rect 22092 6748 22148 6804
rect 21868 6300 21924 6356
rect 20860 5068 20916 5124
rect 21084 5404 21140 5460
rect 21308 5346 21364 5348
rect 21308 5294 21310 5346
rect 21310 5294 21362 5346
rect 21362 5294 21364 5346
rect 21308 5292 21364 5294
rect 20532 4730 20588 4732
rect 20532 4678 20534 4730
rect 20534 4678 20586 4730
rect 20586 4678 20588 4730
rect 20532 4676 20588 4678
rect 20636 4730 20692 4732
rect 20636 4678 20638 4730
rect 20638 4678 20690 4730
rect 20690 4678 20692 4730
rect 20636 4676 20692 4678
rect 20740 4730 20796 4732
rect 20740 4678 20742 4730
rect 20742 4678 20794 4730
rect 20794 4678 20796 4730
rect 20740 4676 20796 4678
rect 21084 4732 21140 4788
rect 20748 4508 20804 4564
rect 20532 3162 20588 3164
rect 20532 3110 20534 3162
rect 20534 3110 20586 3162
rect 20586 3110 20588 3162
rect 20532 3108 20588 3110
rect 20636 3162 20692 3164
rect 20636 3110 20638 3162
rect 20638 3110 20690 3162
rect 20690 3110 20692 3162
rect 20636 3108 20692 3110
rect 20740 3162 20796 3164
rect 20740 3110 20742 3162
rect 20742 3110 20794 3162
rect 20794 3110 20796 3162
rect 20740 3108 20796 3110
rect 21644 5180 21700 5236
rect 22316 8652 22372 8708
rect 22876 9548 22932 9604
rect 22876 8652 22932 8708
rect 22316 6300 22372 6356
rect 23100 11170 23156 11172
rect 23100 11118 23102 11170
rect 23102 11118 23154 11170
rect 23154 11118 23156 11170
rect 23100 11116 23156 11118
rect 23100 9996 23156 10052
rect 22764 8204 22820 8260
rect 22428 5180 22484 5236
rect 22316 5122 22372 5124
rect 22316 5070 22318 5122
rect 22318 5070 22370 5122
rect 22370 5070 22372 5122
rect 22316 5068 22372 5070
rect 22204 5010 22260 5012
rect 22204 4958 22206 5010
rect 22206 4958 22258 5010
rect 22258 4958 22260 5010
rect 22204 4956 22260 4958
rect 23100 9100 23156 9156
rect 22876 7532 22932 7588
rect 22988 7308 23044 7364
rect 22876 7084 22932 7140
rect 23436 11506 23492 11508
rect 23436 11454 23438 11506
rect 23438 11454 23490 11506
rect 23490 11454 23492 11506
rect 23436 11452 23492 11454
rect 23324 11228 23380 11284
rect 23436 9212 23492 9268
rect 23548 8988 23604 9044
rect 23660 8316 23716 8372
rect 23772 9660 23828 9716
rect 22764 5906 22820 5908
rect 22764 5854 22766 5906
rect 22766 5854 22818 5906
rect 22818 5854 22820 5906
rect 22764 5852 22820 5854
rect 23212 7084 23268 7140
rect 22764 5346 22820 5348
rect 22764 5294 22766 5346
rect 22766 5294 22818 5346
rect 22818 5294 22820 5346
rect 22764 5292 22820 5294
rect 22988 6578 23044 6580
rect 22988 6526 22990 6578
rect 22990 6526 23042 6578
rect 23042 6526 23044 6578
rect 22988 6524 23044 6526
rect 22988 6300 23044 6356
rect 23100 6076 23156 6132
rect 23436 6524 23492 6580
rect 23324 6466 23380 6468
rect 23324 6414 23326 6466
rect 23326 6414 23378 6466
rect 23378 6414 23380 6466
rect 23324 6412 23380 6414
rect 22876 4844 22932 4900
rect 22092 4396 22148 4452
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 22540 3500 22596 3556
rect 23324 5010 23380 5012
rect 23324 4958 23326 5010
rect 23326 4958 23378 5010
rect 23378 4958 23380 5010
rect 23324 4956 23380 4958
rect 23324 4508 23380 4564
rect 23660 5740 23716 5796
rect 23548 5516 23604 5572
rect 23884 8370 23940 8372
rect 23884 8318 23886 8370
rect 23886 8318 23938 8370
rect 23938 8318 23940 8370
rect 23884 8316 23940 8318
rect 23884 7532 23940 7588
rect 24108 12738 24164 12740
rect 24108 12686 24110 12738
rect 24110 12686 24162 12738
rect 24162 12686 24164 12738
rect 24108 12684 24164 12686
rect 24220 12348 24276 12404
rect 24220 9212 24276 9268
rect 24108 9154 24164 9156
rect 24108 9102 24110 9154
rect 24110 9102 24162 9154
rect 24162 9102 24164 9154
rect 24108 9100 24164 9102
rect 24220 8876 24276 8932
rect 24108 8092 24164 8148
rect 25004 12738 25060 12740
rect 25004 12686 25006 12738
rect 25006 12686 25058 12738
rect 25058 12686 25060 12738
rect 25004 12684 25060 12686
rect 24444 11116 24500 11172
rect 24556 10668 24612 10724
rect 24332 8258 24388 8260
rect 24332 8206 24334 8258
rect 24334 8206 24386 8258
rect 24386 8206 24388 8258
rect 24332 8204 24388 8206
rect 24444 9996 24500 10052
rect 24444 9772 24500 9828
rect 24220 7532 24276 7588
rect 24332 7868 24388 7924
rect 24108 7474 24164 7476
rect 24108 7422 24110 7474
rect 24110 7422 24162 7474
rect 24162 7422 24164 7474
rect 24108 7420 24164 7422
rect 23996 7084 24052 7140
rect 23884 5964 23940 6020
rect 24220 6860 24276 6916
rect 24108 5740 24164 5796
rect 23436 5122 23492 5124
rect 23436 5070 23438 5122
rect 23438 5070 23490 5122
rect 23490 5070 23492 5122
rect 23436 5068 23492 5070
rect 23100 4338 23156 4340
rect 23100 4286 23102 4338
rect 23102 4286 23154 4338
rect 23154 4286 23156 4338
rect 23100 4284 23156 4286
rect 23772 4844 23828 4900
rect 23884 4284 23940 4340
rect 23884 4114 23940 4116
rect 23884 4062 23886 4114
rect 23886 4062 23938 4114
rect 23938 4062 23940 4114
rect 23884 4060 23940 4062
rect 24668 8204 24724 8260
rect 24556 7196 24612 7252
rect 24556 6860 24612 6916
rect 24332 6130 24388 6132
rect 24332 6078 24334 6130
rect 24334 6078 24386 6130
rect 24386 6078 24388 6130
rect 24332 6076 24388 6078
rect 25900 12738 25956 12740
rect 25900 12686 25902 12738
rect 25902 12686 25954 12738
rect 25954 12686 25956 12738
rect 25900 12684 25956 12686
rect 25452 12402 25508 12404
rect 25452 12350 25454 12402
rect 25454 12350 25506 12402
rect 25506 12350 25508 12402
rect 25452 12348 25508 12350
rect 25340 11788 25396 11844
rect 26236 12066 26292 12068
rect 26236 12014 26238 12066
rect 26238 12014 26290 12066
rect 26290 12014 26292 12066
rect 26236 12012 26292 12014
rect 25788 11900 25844 11956
rect 25228 10722 25284 10724
rect 25228 10670 25230 10722
rect 25230 10670 25282 10722
rect 25282 10670 25284 10722
rect 25228 10668 25284 10670
rect 26124 11452 26180 11508
rect 25788 10220 25844 10276
rect 25228 10108 25284 10164
rect 24444 6748 24500 6804
rect 24220 5628 24276 5684
rect 24332 5068 24388 5124
rect 24108 4732 24164 4788
rect 24220 4562 24276 4564
rect 24220 4510 24222 4562
rect 24222 4510 24274 4562
rect 24274 4510 24276 4562
rect 24220 4508 24276 4510
rect 23996 3724 24052 3780
rect 24108 4172 24164 4228
rect 24668 6300 24724 6356
rect 24668 5906 24724 5908
rect 24668 5854 24670 5906
rect 24670 5854 24722 5906
rect 24722 5854 24724 5906
rect 24668 5852 24724 5854
rect 24668 5628 24724 5684
rect 24780 5292 24836 5348
rect 24668 4172 24724 4228
rect 25004 8428 25060 8484
rect 25116 8370 25172 8372
rect 25116 8318 25118 8370
rect 25118 8318 25170 8370
rect 25170 8318 25172 8370
rect 25116 8316 25172 8318
rect 25900 10108 25956 10164
rect 25788 9602 25844 9604
rect 25788 9550 25790 9602
rect 25790 9550 25842 9602
rect 25842 9550 25844 9602
rect 25788 9548 25844 9550
rect 26236 11116 26292 11172
rect 26236 10444 26292 10500
rect 25340 9212 25396 9268
rect 25676 9154 25732 9156
rect 25676 9102 25678 9154
rect 25678 9102 25730 9154
rect 25730 9102 25732 9154
rect 25676 9100 25732 9102
rect 25228 6748 25284 6804
rect 25116 6300 25172 6356
rect 25004 6188 25060 6244
rect 26684 11900 26740 11956
rect 26796 12012 26852 12068
rect 28812 16940 28868 16996
rect 26460 10220 26516 10276
rect 26012 9212 26068 9268
rect 25900 7586 25956 7588
rect 25900 7534 25902 7586
rect 25902 7534 25954 7586
rect 25954 7534 25956 7586
rect 25900 7532 25956 7534
rect 26012 7420 26068 7476
rect 25564 7084 25620 7140
rect 25900 7196 25956 7252
rect 25340 6300 25396 6356
rect 25676 6300 25732 6356
rect 25116 5628 25172 5684
rect 24892 4732 24948 4788
rect 24780 3948 24836 4004
rect 25228 6076 25284 6132
rect 24892 3500 24948 3556
rect 24668 3388 24724 3444
rect 25116 3612 25172 3668
rect 24892 1260 24948 1316
rect 25340 5404 25396 5460
rect 25900 6412 25956 6468
rect 26012 4956 26068 5012
rect 25788 4732 25844 4788
rect 25676 2492 25732 2548
rect 25900 4450 25956 4452
rect 25900 4398 25902 4450
rect 25902 4398 25954 4450
rect 25954 4398 25956 4450
rect 25900 4396 25956 4398
rect 25900 4172 25956 4228
rect 25900 3554 25956 3556
rect 25900 3502 25902 3554
rect 25902 3502 25954 3554
rect 25954 3502 25956 3554
rect 25900 3500 25956 3502
rect 26124 4172 26180 4228
rect 26124 3778 26180 3780
rect 26124 3726 26126 3778
rect 26126 3726 26178 3778
rect 26178 3726 26180 3778
rect 26124 3724 26180 3726
rect 26348 9154 26404 9156
rect 26348 9102 26350 9154
rect 26350 9102 26402 9154
rect 26402 9102 26404 9154
rect 26348 9100 26404 9102
rect 27244 11170 27300 11172
rect 27244 11118 27246 11170
rect 27246 11118 27298 11170
rect 27298 11118 27300 11170
rect 27244 11116 27300 11118
rect 26684 9100 26740 9156
rect 27244 10498 27300 10500
rect 27244 10446 27246 10498
rect 27246 10446 27298 10498
rect 27298 10446 27300 10498
rect 27244 10444 27300 10446
rect 26348 7644 26404 7700
rect 26572 7644 26628 7700
rect 26460 7308 26516 7364
rect 26572 6636 26628 6692
rect 26572 5516 26628 5572
rect 26348 4898 26404 4900
rect 26348 4846 26350 4898
rect 26350 4846 26402 4898
rect 26402 4846 26404 4898
rect 26348 4844 26404 4846
rect 26348 4338 26404 4340
rect 26348 4286 26350 4338
rect 26350 4286 26402 4338
rect 26402 4286 26404 4338
rect 26348 4284 26404 4286
rect 26796 8092 26852 8148
rect 26908 9884 26964 9940
rect 26796 7868 26852 7924
rect 27132 8316 27188 8372
rect 27020 8092 27076 8148
rect 27020 7644 27076 7700
rect 27244 8204 27300 8260
rect 27244 7756 27300 7812
rect 27244 7586 27300 7588
rect 27244 7534 27246 7586
rect 27246 7534 27298 7586
rect 27298 7534 27300 7586
rect 27244 7532 27300 7534
rect 28252 15596 28308 15652
rect 27804 10668 27860 10724
rect 27580 9938 27636 9940
rect 27580 9886 27582 9938
rect 27582 9886 27634 9938
rect 27634 9886 27636 9938
rect 27580 9884 27636 9886
rect 27356 7196 27412 7252
rect 27692 8204 27748 8260
rect 28252 11506 28308 11508
rect 28252 11454 28254 11506
rect 28254 11454 28306 11506
rect 28306 11454 28308 11506
rect 28252 11452 28308 11454
rect 28028 10108 28084 10164
rect 27916 9996 27972 10052
rect 28140 9826 28196 9828
rect 28140 9774 28142 9826
rect 28142 9774 28194 9826
rect 28194 9774 28196 9826
rect 28140 9772 28196 9774
rect 30192 16490 30248 16492
rect 30192 16438 30194 16490
rect 30194 16438 30246 16490
rect 30246 16438 30248 16490
rect 30192 16436 30248 16438
rect 30296 16490 30352 16492
rect 30296 16438 30298 16490
rect 30298 16438 30350 16490
rect 30350 16438 30352 16490
rect 30296 16436 30352 16438
rect 30400 16490 30456 16492
rect 30400 16438 30402 16490
rect 30402 16438 30454 16490
rect 30454 16438 30456 16490
rect 30400 16436 30456 16438
rect 31836 15820 31892 15876
rect 31276 15484 31332 15540
rect 31948 15708 32004 15764
rect 31948 15484 32004 15540
rect 32508 15596 32564 15652
rect 30192 14922 30248 14924
rect 30192 14870 30194 14922
rect 30194 14870 30246 14922
rect 30246 14870 30248 14922
rect 30192 14868 30248 14870
rect 30296 14922 30352 14924
rect 30296 14870 30298 14922
rect 30298 14870 30350 14922
rect 30350 14870 30352 14922
rect 30296 14868 30352 14870
rect 30400 14922 30456 14924
rect 30400 14870 30402 14922
rect 30402 14870 30454 14922
rect 30454 14870 30456 14922
rect 30400 14868 30456 14870
rect 28588 11170 28644 11172
rect 28588 11118 28590 11170
rect 28590 11118 28642 11170
rect 28642 11118 28644 11170
rect 28588 11116 28644 11118
rect 28700 9996 28756 10052
rect 28700 9212 28756 9268
rect 27916 8316 27972 8372
rect 27692 7980 27748 8036
rect 28140 8146 28196 8148
rect 28140 8094 28142 8146
rect 28142 8094 28194 8146
rect 28194 8094 28196 8146
rect 28140 8092 28196 8094
rect 27580 7196 27636 7252
rect 27692 7420 27748 7476
rect 26796 6636 26852 6692
rect 26908 6412 26964 6468
rect 26796 6300 26852 6356
rect 26796 5740 26852 5796
rect 26684 5180 26740 5236
rect 27356 6300 27412 6356
rect 27244 5180 27300 5236
rect 26796 4844 26852 4900
rect 26908 4620 26964 4676
rect 26684 4226 26740 4228
rect 26684 4174 26686 4226
rect 26686 4174 26738 4226
rect 26738 4174 26740 4226
rect 26684 4172 26740 4174
rect 26460 3612 26516 3668
rect 26572 3948 26628 4004
rect 27804 6636 27860 6692
rect 27916 7196 27972 7252
rect 27804 6018 27860 6020
rect 27804 5966 27806 6018
rect 27806 5966 27858 6018
rect 27858 5966 27860 6018
rect 27804 5964 27860 5966
rect 28028 6860 28084 6916
rect 28140 7084 28196 7140
rect 28028 6636 28084 6692
rect 28028 6076 28084 6132
rect 27580 5516 27636 5572
rect 27804 5292 27860 5348
rect 28364 8204 28420 8260
rect 28476 7084 28532 7140
rect 28364 6860 28420 6916
rect 28588 6860 28644 6916
rect 28588 6300 28644 6356
rect 28364 5404 28420 5460
rect 27356 4060 27412 4116
rect 27692 4562 27748 4564
rect 27692 4510 27694 4562
rect 27694 4510 27746 4562
rect 27746 4510 27748 4562
rect 27692 4508 27748 4510
rect 27580 3948 27636 4004
rect 27692 4284 27748 4340
rect 27580 3666 27636 3668
rect 27580 3614 27582 3666
rect 27582 3614 27634 3666
rect 27634 3614 27636 3666
rect 27580 3612 27636 3614
rect 27132 3554 27188 3556
rect 27132 3502 27134 3554
rect 27134 3502 27186 3554
rect 27186 3502 27188 3554
rect 27132 3500 27188 3502
rect 26684 3330 26740 3332
rect 26684 3278 26686 3330
rect 26686 3278 26738 3330
rect 26738 3278 26740 3330
rect 26684 3276 26740 3278
rect 26348 2268 26404 2324
rect 28140 4956 28196 5012
rect 27916 3164 27972 3220
rect 27132 924 27188 980
rect 28476 6188 28532 6244
rect 28252 3276 28308 3332
rect 28028 924 28084 980
rect 28700 4284 28756 4340
rect 28588 3836 28644 3892
rect 28924 13692 28980 13748
rect 30192 13354 30248 13356
rect 30192 13302 30194 13354
rect 30194 13302 30246 13354
rect 30246 13302 30248 13354
rect 30192 13300 30248 13302
rect 30296 13354 30352 13356
rect 30296 13302 30298 13354
rect 30298 13302 30350 13354
rect 30350 13302 30352 13354
rect 30296 13300 30352 13302
rect 30400 13354 30456 13356
rect 30400 13302 30402 13354
rect 30402 13302 30454 13354
rect 30454 13302 30456 13354
rect 30400 13300 30456 13302
rect 30044 12236 30100 12292
rect 29260 11170 29316 11172
rect 29260 11118 29262 11170
rect 29262 11118 29314 11170
rect 29314 11118 29316 11170
rect 29260 11116 29316 11118
rect 29148 10780 29204 10836
rect 28924 8316 28980 8372
rect 29036 8540 29092 8596
rect 28924 7756 28980 7812
rect 29260 10444 29316 10500
rect 29932 11228 29988 11284
rect 29484 8764 29540 8820
rect 29820 10556 29876 10612
rect 29820 10108 29876 10164
rect 29932 9938 29988 9940
rect 29932 9886 29934 9938
rect 29934 9886 29986 9938
rect 29986 9886 29988 9938
rect 29932 9884 29988 9886
rect 29596 9212 29652 9268
rect 29820 8930 29876 8932
rect 29820 8878 29822 8930
rect 29822 8878 29874 8930
rect 29874 8878 29876 8930
rect 29820 8876 29876 8878
rect 29596 8540 29652 8596
rect 29708 8652 29764 8708
rect 29484 7868 29540 7924
rect 29036 7084 29092 7140
rect 29372 6802 29428 6804
rect 29372 6750 29374 6802
rect 29374 6750 29426 6802
rect 29426 6750 29428 6802
rect 29372 6748 29428 6750
rect 29260 6412 29316 6468
rect 29372 6524 29428 6580
rect 29260 5180 29316 5236
rect 29148 4620 29204 4676
rect 29036 4396 29092 4452
rect 28812 3612 28868 3668
rect 29596 6972 29652 7028
rect 29820 7698 29876 7700
rect 29820 7646 29822 7698
rect 29822 7646 29874 7698
rect 29874 7646 29876 7698
rect 29820 7644 29876 7646
rect 29708 6076 29764 6132
rect 30492 12012 30548 12068
rect 30192 11786 30248 11788
rect 30192 11734 30194 11786
rect 30194 11734 30246 11786
rect 30246 11734 30248 11786
rect 30192 11732 30248 11734
rect 30296 11786 30352 11788
rect 30296 11734 30298 11786
rect 30298 11734 30350 11786
rect 30350 11734 30352 11786
rect 30296 11732 30352 11734
rect 30400 11786 30456 11788
rect 30400 11734 30402 11786
rect 30402 11734 30454 11786
rect 30454 11734 30456 11786
rect 30400 11732 30456 11734
rect 30604 10668 30660 10724
rect 30192 10218 30248 10220
rect 30192 10166 30194 10218
rect 30194 10166 30246 10218
rect 30246 10166 30248 10218
rect 30192 10164 30248 10166
rect 30296 10218 30352 10220
rect 30296 10166 30298 10218
rect 30298 10166 30350 10218
rect 30350 10166 30352 10218
rect 30296 10164 30352 10166
rect 30400 10218 30456 10220
rect 30400 10166 30402 10218
rect 30402 10166 30454 10218
rect 30454 10166 30456 10218
rect 30400 10164 30456 10166
rect 30492 9996 30548 10052
rect 30192 8650 30248 8652
rect 30192 8598 30194 8650
rect 30194 8598 30246 8650
rect 30246 8598 30248 8650
rect 30192 8596 30248 8598
rect 30296 8650 30352 8652
rect 30296 8598 30298 8650
rect 30298 8598 30350 8650
rect 30350 8598 30352 8650
rect 30296 8596 30352 8598
rect 30400 8650 30456 8652
rect 30400 8598 30402 8650
rect 30402 8598 30454 8650
rect 30454 8598 30456 8650
rect 30400 8596 30456 8598
rect 30940 14028 30996 14084
rect 30828 10444 30884 10500
rect 32172 13356 32228 13412
rect 31612 13244 31668 13300
rect 31052 11900 31108 11956
rect 31164 12124 31220 12180
rect 31164 11228 31220 11284
rect 31164 10610 31220 10612
rect 31164 10558 31166 10610
rect 31166 10558 31218 10610
rect 31218 10558 31220 10610
rect 31164 10556 31220 10558
rect 31388 12066 31444 12068
rect 31388 12014 31390 12066
rect 31390 12014 31442 12066
rect 31442 12014 31444 12066
rect 31388 12012 31444 12014
rect 30268 7980 30324 8036
rect 30044 7868 30100 7924
rect 30604 8204 30660 8260
rect 30716 7644 30772 7700
rect 30940 8764 30996 8820
rect 30192 7082 30248 7084
rect 30192 7030 30194 7082
rect 30194 7030 30246 7082
rect 30246 7030 30248 7082
rect 30192 7028 30248 7030
rect 30296 7082 30352 7084
rect 30296 7030 30298 7082
rect 30298 7030 30350 7082
rect 30350 7030 30352 7082
rect 30296 7028 30352 7030
rect 30400 7082 30456 7084
rect 30400 7030 30402 7082
rect 30402 7030 30454 7082
rect 30454 7030 30456 7082
rect 30400 7028 30456 7030
rect 30604 7084 30660 7140
rect 29932 5906 29988 5908
rect 29932 5854 29934 5906
rect 29934 5854 29986 5906
rect 29986 5854 29988 5906
rect 29932 5852 29988 5854
rect 31500 9996 31556 10052
rect 31612 12684 31668 12740
rect 30604 5740 30660 5796
rect 31388 9154 31444 9156
rect 31388 9102 31390 9154
rect 31390 9102 31442 9154
rect 31442 9102 31444 9154
rect 31388 9100 31444 9102
rect 31500 9042 31556 9044
rect 31500 8990 31502 9042
rect 31502 8990 31554 9042
rect 31554 8990 31556 9042
rect 31500 8988 31556 8990
rect 31164 8876 31220 8932
rect 31388 8876 31444 8932
rect 29820 5122 29876 5124
rect 29820 5070 29822 5122
rect 29822 5070 29874 5122
rect 29874 5070 29876 5122
rect 29820 5068 29876 5070
rect 30192 5514 30248 5516
rect 30192 5462 30194 5514
rect 30194 5462 30246 5514
rect 30246 5462 30248 5514
rect 30192 5460 30248 5462
rect 30296 5514 30352 5516
rect 30296 5462 30298 5514
rect 30298 5462 30350 5514
rect 30350 5462 30352 5514
rect 30296 5460 30352 5462
rect 30400 5514 30456 5516
rect 30400 5462 30402 5514
rect 30402 5462 30454 5514
rect 30454 5462 30456 5514
rect 30400 5460 30456 5462
rect 30492 5234 30548 5236
rect 30492 5182 30494 5234
rect 30494 5182 30546 5234
rect 30546 5182 30548 5234
rect 30492 5180 30548 5182
rect 30604 5122 30660 5124
rect 30604 5070 30606 5122
rect 30606 5070 30658 5122
rect 30658 5070 30660 5122
rect 30604 5068 30660 5070
rect 31052 5964 31108 6020
rect 30716 4844 30772 4900
rect 29372 4172 29428 4228
rect 30192 3946 30248 3948
rect 30192 3894 30194 3946
rect 30194 3894 30246 3946
rect 30246 3894 30248 3946
rect 30192 3892 30248 3894
rect 30296 3946 30352 3948
rect 30296 3894 30298 3946
rect 30298 3894 30350 3946
rect 30350 3894 30352 3946
rect 30296 3892 30352 3894
rect 30400 3946 30456 3948
rect 30400 3894 30402 3946
rect 30402 3894 30454 3946
rect 30454 3894 30456 3946
rect 30400 3892 30456 3894
rect 29148 3164 29204 3220
rect 29820 3388 29876 3444
rect 30940 4844 30996 4900
rect 31276 8764 31332 8820
rect 31276 6188 31332 6244
rect 31836 12290 31892 12292
rect 31836 12238 31838 12290
rect 31838 12238 31890 12290
rect 31890 12238 31892 12290
rect 31836 12236 31892 12238
rect 31724 12124 31780 12180
rect 31724 11900 31780 11956
rect 34748 15596 34804 15652
rect 33404 13804 33460 13860
rect 33292 13692 33348 13748
rect 32284 12124 32340 12180
rect 32396 12066 32452 12068
rect 32396 12014 32398 12066
rect 32398 12014 32450 12066
rect 32450 12014 32452 12066
rect 32396 12012 32452 12014
rect 32284 10386 32340 10388
rect 32284 10334 32286 10386
rect 32286 10334 32338 10386
rect 32338 10334 32340 10386
rect 32284 10332 32340 10334
rect 32172 9996 32228 10052
rect 31612 7980 31668 8036
rect 31948 8428 32004 8484
rect 32396 9772 32452 9828
rect 32844 11394 32900 11396
rect 32844 11342 32846 11394
rect 32846 11342 32898 11394
rect 32898 11342 32900 11394
rect 32844 11340 32900 11342
rect 32956 11004 33012 11060
rect 33292 12738 33348 12740
rect 33292 12686 33294 12738
rect 33294 12686 33346 12738
rect 33346 12686 33348 12738
rect 33292 12684 33348 12686
rect 33516 11954 33572 11956
rect 33516 11902 33518 11954
rect 33518 11902 33570 11954
rect 33570 11902 33572 11954
rect 33516 11900 33572 11902
rect 34524 13692 34580 13748
rect 33852 12012 33908 12068
rect 34636 11788 34692 11844
rect 32844 10444 32900 10500
rect 32620 8876 32676 8932
rect 33068 10332 33124 10388
rect 33628 10780 33684 10836
rect 33852 11004 33908 11060
rect 33292 9772 33348 9828
rect 32508 8092 32564 8148
rect 33068 7980 33124 8036
rect 32060 7196 32116 7252
rect 31948 4844 32004 4900
rect 31164 4508 31220 4564
rect 31052 2380 31108 2436
rect 32396 3724 32452 3780
rect 33180 7362 33236 7364
rect 33180 7310 33182 7362
rect 33182 7310 33234 7362
rect 33234 7310 33236 7362
rect 33180 7308 33236 7310
rect 32284 3500 32340 3556
rect 32732 1484 32788 1540
rect 32732 924 32788 980
rect 33516 9772 33572 9828
rect 34412 9884 34468 9940
rect 33740 9324 33796 9380
rect 33516 9212 33572 9268
rect 33404 8876 33460 8932
rect 33628 8316 33684 8372
rect 33516 8092 33572 8148
rect 33628 7644 33684 7700
rect 33180 6018 33236 6020
rect 33180 5966 33182 6018
rect 33182 5966 33234 6018
rect 33234 5966 33236 6018
rect 33180 5964 33236 5966
rect 33292 6636 33348 6692
rect 33068 4060 33124 4116
rect 33628 4284 33684 4340
rect 48300 17052 48356 17108
rect 42252 16828 42308 16884
rect 39852 15706 39908 15708
rect 39852 15654 39854 15706
rect 39854 15654 39906 15706
rect 39906 15654 39908 15706
rect 39852 15652 39908 15654
rect 39956 15706 40012 15708
rect 39956 15654 39958 15706
rect 39958 15654 40010 15706
rect 40010 15654 40012 15706
rect 39956 15652 40012 15654
rect 40060 15706 40116 15708
rect 40060 15654 40062 15706
rect 40062 15654 40114 15706
rect 40114 15654 40116 15706
rect 40060 15652 40116 15654
rect 35756 14028 35812 14084
rect 35308 13858 35364 13860
rect 35308 13806 35310 13858
rect 35310 13806 35362 13858
rect 35362 13806 35364 13858
rect 35308 13804 35364 13806
rect 37100 13692 37156 13748
rect 36316 12962 36372 12964
rect 36316 12910 36318 12962
rect 36318 12910 36370 12962
rect 36370 12910 36372 12962
rect 36316 12908 36372 12910
rect 35420 12572 35476 12628
rect 35308 11340 35364 11396
rect 35420 11004 35476 11060
rect 34972 9996 35028 10052
rect 34076 8876 34132 8932
rect 34188 9660 34244 9716
rect 34636 9266 34692 9268
rect 34636 9214 34638 9266
rect 34638 9214 34690 9266
rect 34690 9214 34692 9266
rect 34636 9212 34692 9214
rect 35196 8876 35252 8932
rect 34860 8764 34916 8820
rect 34188 8316 34244 8372
rect 34412 8428 34468 8484
rect 34412 8258 34468 8260
rect 34412 8206 34414 8258
rect 34414 8206 34466 8258
rect 34466 8206 34468 8258
rect 34412 8204 34468 8206
rect 34412 7980 34468 8036
rect 34412 7474 34468 7476
rect 34412 7422 34414 7474
rect 34414 7422 34466 7474
rect 34466 7422 34468 7474
rect 34412 7420 34468 7422
rect 33852 6748 33908 6804
rect 33964 4508 34020 4564
rect 33740 3948 33796 4004
rect 33628 3500 33684 3556
rect 33180 3388 33236 3444
rect 33068 1484 33124 1540
rect 33068 1036 33124 1092
rect 34524 4450 34580 4452
rect 34524 4398 34526 4450
rect 34526 4398 34578 4450
rect 34578 4398 34580 4450
rect 34524 4396 34580 4398
rect 34860 7868 34916 7924
rect 35084 7644 35140 7700
rect 34972 6636 35028 6692
rect 34412 3666 34468 3668
rect 34412 3614 34414 3666
rect 34414 3614 34466 3666
rect 34466 3614 34468 3666
rect 34412 3612 34468 3614
rect 35532 12124 35588 12180
rect 35980 11788 36036 11844
rect 35644 10892 35700 10948
rect 35532 10444 35588 10500
rect 35532 9100 35588 9156
rect 35756 9996 35812 10052
rect 35868 9938 35924 9940
rect 35868 9886 35870 9938
rect 35870 9886 35922 9938
rect 35922 9886 35924 9938
rect 35868 9884 35924 9886
rect 36988 12962 37044 12964
rect 36988 12910 36990 12962
rect 36990 12910 37042 12962
rect 37042 12910 37044 12962
rect 36988 12908 37044 12910
rect 37212 12460 37268 12516
rect 37324 12012 37380 12068
rect 37548 13356 37604 13412
rect 37100 11676 37156 11732
rect 36316 11394 36372 11396
rect 36316 11342 36318 11394
rect 36318 11342 36370 11394
rect 36370 11342 36372 11394
rect 36316 11340 36372 11342
rect 36092 9212 36148 9268
rect 35868 8316 35924 8372
rect 35868 7644 35924 7700
rect 35308 3276 35364 3332
rect 35308 2492 35364 2548
rect 35644 3612 35700 3668
rect 36652 10498 36708 10500
rect 36652 10446 36654 10498
rect 36654 10446 36706 10498
rect 36706 10446 36708 10498
rect 36652 10444 36708 10446
rect 36428 10050 36484 10052
rect 36428 9998 36430 10050
rect 36430 9998 36482 10050
rect 36482 9998 36484 10050
rect 36428 9996 36484 9998
rect 36316 8988 36372 9044
rect 36316 8540 36372 8596
rect 36204 7474 36260 7476
rect 36204 7422 36206 7474
rect 36206 7422 36258 7474
rect 36258 7422 36260 7474
rect 36204 7420 36260 7422
rect 36652 8988 36708 9044
rect 36316 6636 36372 6692
rect 35980 6524 36036 6580
rect 36428 6524 36484 6580
rect 35980 5180 36036 5236
rect 37772 13074 37828 13076
rect 37772 13022 37774 13074
rect 37774 13022 37826 13074
rect 37826 13022 37828 13074
rect 37772 13020 37828 13022
rect 37660 12684 37716 12740
rect 37660 11788 37716 11844
rect 37884 11676 37940 11732
rect 37548 10892 37604 10948
rect 37100 9996 37156 10052
rect 36764 7420 36820 7476
rect 36988 9826 37044 9828
rect 36988 9774 36990 9826
rect 36990 9774 37042 9826
rect 37042 9774 37044 9826
rect 36988 9772 37044 9774
rect 37212 9660 37268 9716
rect 37436 8988 37492 9044
rect 37212 8876 37268 8932
rect 37548 8930 37604 8932
rect 37548 8878 37550 8930
rect 37550 8878 37602 8930
rect 37602 8878 37604 8930
rect 37548 8876 37604 8878
rect 37100 8764 37156 8820
rect 37548 8652 37604 8708
rect 37436 8370 37492 8372
rect 37436 8318 37438 8370
rect 37438 8318 37490 8370
rect 37490 8318 37492 8370
rect 37436 8316 37492 8318
rect 37212 8146 37268 8148
rect 37212 8094 37214 8146
rect 37214 8094 37266 8146
rect 37266 8094 37268 8146
rect 37212 8092 37268 8094
rect 36652 4508 36708 4564
rect 37212 5180 37268 5236
rect 36988 3724 37044 3780
rect 36316 3276 36372 3332
rect 38108 13804 38164 13860
rect 38220 11282 38276 11284
rect 38220 11230 38222 11282
rect 38222 11230 38274 11282
rect 38274 11230 38276 11282
rect 38220 11228 38276 11230
rect 37996 10332 38052 10388
rect 38108 9100 38164 9156
rect 37996 8764 38052 8820
rect 37884 8092 37940 8148
rect 37884 7420 37940 7476
rect 38108 8540 38164 8596
rect 37772 7308 37828 7364
rect 37996 6690 38052 6692
rect 37996 6638 37998 6690
rect 37998 6638 38050 6690
rect 38050 6638 38052 6690
rect 37996 6636 38052 6638
rect 37660 5516 37716 5572
rect 37772 6524 37828 6580
rect 39852 14138 39908 14140
rect 39852 14086 39854 14138
rect 39854 14086 39906 14138
rect 39906 14086 39908 14138
rect 39852 14084 39908 14086
rect 39956 14138 40012 14140
rect 39956 14086 39958 14138
rect 39958 14086 40010 14138
rect 40010 14086 40012 14138
rect 39956 14084 40012 14086
rect 40060 14138 40116 14140
rect 40060 14086 40062 14138
rect 40062 14086 40114 14138
rect 40114 14086 40116 14138
rect 40060 14084 40116 14086
rect 39900 13858 39956 13860
rect 39900 13806 39902 13858
rect 39902 13806 39954 13858
rect 39954 13806 39956 13858
rect 39900 13804 39956 13806
rect 40572 13580 40628 13636
rect 40236 13132 40292 13188
rect 38892 13020 38948 13076
rect 38556 12460 38612 12516
rect 38892 12012 38948 12068
rect 39116 11900 39172 11956
rect 39004 10780 39060 10836
rect 38556 8988 38612 9044
rect 38556 8764 38612 8820
rect 38668 7980 38724 8036
rect 38444 7756 38500 7812
rect 38556 7698 38612 7700
rect 38556 7646 38558 7698
rect 38558 7646 38610 7698
rect 38610 7646 38612 7698
rect 38556 7644 38612 7646
rect 38892 8876 38948 8932
rect 40236 12796 40292 12852
rect 39852 12570 39908 12572
rect 39852 12518 39854 12570
rect 39854 12518 39906 12570
rect 39906 12518 39908 12570
rect 39852 12516 39908 12518
rect 39956 12570 40012 12572
rect 39956 12518 39958 12570
rect 39958 12518 40010 12570
rect 40010 12518 40012 12570
rect 39956 12516 40012 12518
rect 40060 12570 40116 12572
rect 40060 12518 40062 12570
rect 40062 12518 40114 12570
rect 40114 12518 40116 12570
rect 40060 12516 40116 12518
rect 40460 12572 40516 12628
rect 41468 13468 41524 13524
rect 40796 12348 40852 12404
rect 39452 10386 39508 10388
rect 39452 10334 39454 10386
rect 39454 10334 39506 10386
rect 39506 10334 39508 10386
rect 39452 10332 39508 10334
rect 39340 10108 39396 10164
rect 39900 11954 39956 11956
rect 39900 11902 39902 11954
rect 39902 11902 39954 11954
rect 39954 11902 39956 11954
rect 39900 11900 39956 11902
rect 39676 11116 39732 11172
rect 39852 11002 39908 11004
rect 39852 10950 39854 11002
rect 39854 10950 39906 11002
rect 39906 10950 39908 11002
rect 39852 10948 39908 10950
rect 39956 11002 40012 11004
rect 39956 10950 39958 11002
rect 39958 10950 40010 11002
rect 40010 10950 40012 11002
rect 39956 10948 40012 10950
rect 40060 11002 40116 11004
rect 40060 10950 40062 11002
rect 40062 10950 40114 11002
rect 40114 10950 40116 11002
rect 40060 10948 40116 10950
rect 40348 12178 40404 12180
rect 40348 12126 40350 12178
rect 40350 12126 40402 12178
rect 40402 12126 40404 12178
rect 40348 12124 40404 12126
rect 39564 9884 39620 9940
rect 39228 9772 39284 9828
rect 39228 8876 39284 8932
rect 39452 9548 39508 9604
rect 38892 7532 38948 7588
rect 38220 7362 38276 7364
rect 38220 7310 38222 7362
rect 38222 7310 38274 7362
rect 38274 7310 38276 7362
rect 38220 7308 38276 7310
rect 38220 6860 38276 6916
rect 37884 5292 37940 5348
rect 38444 5852 38500 5908
rect 38892 7084 38948 7140
rect 37548 4284 37604 4340
rect 38556 2828 38612 2884
rect 39452 8316 39508 8372
rect 39228 8092 39284 8148
rect 39004 3836 39060 3892
rect 39340 7980 39396 8036
rect 39452 7084 39508 7140
rect 39676 9772 39732 9828
rect 40348 10610 40404 10612
rect 40348 10558 40350 10610
rect 40350 10558 40402 10610
rect 40402 10558 40404 10610
rect 40348 10556 40404 10558
rect 40236 10108 40292 10164
rect 40124 9660 40180 9716
rect 40012 9548 40068 9604
rect 39852 9434 39908 9436
rect 39852 9382 39854 9434
rect 39854 9382 39906 9434
rect 39906 9382 39908 9434
rect 39852 9380 39908 9382
rect 39956 9434 40012 9436
rect 39956 9382 39958 9434
rect 39958 9382 40010 9434
rect 40010 9382 40012 9434
rect 39956 9380 40012 9382
rect 40060 9434 40116 9436
rect 40060 9382 40062 9434
rect 40062 9382 40114 9434
rect 40114 9382 40116 9434
rect 40060 9380 40116 9382
rect 39900 8316 39956 8372
rect 39676 7980 39732 8036
rect 39852 7866 39908 7868
rect 39852 7814 39854 7866
rect 39854 7814 39906 7866
rect 39906 7814 39908 7866
rect 39852 7812 39908 7814
rect 39956 7866 40012 7868
rect 39956 7814 39958 7866
rect 39958 7814 40010 7866
rect 40010 7814 40012 7866
rect 39956 7812 40012 7814
rect 40060 7866 40116 7868
rect 40060 7814 40062 7866
rect 40062 7814 40114 7866
rect 40114 7814 40116 7866
rect 40060 7812 40116 7814
rect 39900 7474 39956 7476
rect 39900 7422 39902 7474
rect 39902 7422 39954 7474
rect 39954 7422 39956 7474
rect 39900 7420 39956 7422
rect 40348 9100 40404 9156
rect 40348 7644 40404 7700
rect 40348 7362 40404 7364
rect 40348 7310 40350 7362
rect 40350 7310 40402 7362
rect 40402 7310 40404 7362
rect 40348 7308 40404 7310
rect 39340 6412 39396 6468
rect 40012 6802 40068 6804
rect 40012 6750 40014 6802
rect 40014 6750 40066 6802
rect 40066 6750 40068 6802
rect 40012 6748 40068 6750
rect 39788 6690 39844 6692
rect 39788 6638 39790 6690
rect 39790 6638 39842 6690
rect 39842 6638 39844 6690
rect 39788 6636 39844 6638
rect 39452 5964 39508 6020
rect 39340 5906 39396 5908
rect 39340 5854 39342 5906
rect 39342 5854 39394 5906
rect 39394 5854 39396 5906
rect 39340 5852 39396 5854
rect 39228 3276 39284 3332
rect 38780 1484 38836 1540
rect 41356 12850 41412 12852
rect 41356 12798 41358 12850
rect 41358 12798 41410 12850
rect 41410 12798 41412 12850
rect 41356 12796 41412 12798
rect 40572 12124 40628 12180
rect 41244 12066 41300 12068
rect 41244 12014 41246 12066
rect 41246 12014 41298 12066
rect 41298 12014 41300 12066
rect 41244 12012 41300 12014
rect 40908 11788 40964 11844
rect 41020 10892 41076 10948
rect 41020 9996 41076 10052
rect 41020 9772 41076 9828
rect 40908 9548 40964 9604
rect 41356 10892 41412 10948
rect 41580 12738 41636 12740
rect 41580 12686 41582 12738
rect 41582 12686 41634 12738
rect 41634 12686 41636 12738
rect 41580 12684 41636 12686
rect 42028 12348 42084 12404
rect 41580 12124 41636 12180
rect 41132 8764 41188 8820
rect 41244 10220 41300 10276
rect 41020 8316 41076 8372
rect 40908 8204 40964 8260
rect 39564 4396 39620 4452
rect 39852 6298 39908 6300
rect 39852 6246 39854 6298
rect 39854 6246 39906 6298
rect 39906 6246 39908 6298
rect 39852 6244 39908 6246
rect 39956 6298 40012 6300
rect 39956 6246 39958 6298
rect 39958 6246 40010 6298
rect 40010 6246 40012 6298
rect 39956 6244 40012 6246
rect 40060 6298 40116 6300
rect 40060 6246 40062 6298
rect 40062 6246 40114 6298
rect 40114 6246 40116 6298
rect 40060 6244 40116 6246
rect 40908 7420 40964 7476
rect 41132 7532 41188 7588
rect 41020 6748 41076 6804
rect 40236 6130 40292 6132
rect 40236 6078 40238 6130
rect 40238 6078 40290 6130
rect 40290 6078 40292 6130
rect 40236 6076 40292 6078
rect 39788 5964 39844 6020
rect 41132 7308 41188 7364
rect 41132 6188 41188 6244
rect 39852 4730 39908 4732
rect 39852 4678 39854 4730
rect 39854 4678 39906 4730
rect 39906 4678 39908 4730
rect 39852 4676 39908 4678
rect 39956 4730 40012 4732
rect 39956 4678 39958 4730
rect 39958 4678 40010 4730
rect 40010 4678 40012 4730
rect 39956 4676 40012 4678
rect 40060 4730 40116 4732
rect 40060 4678 40062 4730
rect 40062 4678 40114 4730
rect 40114 4678 40116 4730
rect 40060 4676 40116 4678
rect 40908 4396 40964 4452
rect 40348 4338 40404 4340
rect 40348 4286 40350 4338
rect 40350 4286 40402 4338
rect 40402 4286 40404 4338
rect 40348 4284 40404 4286
rect 39564 2380 39620 2436
rect 39900 4060 39956 4116
rect 39852 3162 39908 3164
rect 39852 3110 39854 3162
rect 39854 3110 39906 3162
rect 39906 3110 39908 3162
rect 39852 3108 39908 3110
rect 39956 3162 40012 3164
rect 39956 3110 39958 3162
rect 39958 3110 40010 3162
rect 40010 3110 40012 3162
rect 39956 3108 40012 3110
rect 40060 3162 40116 3164
rect 40060 3110 40062 3162
rect 40062 3110 40114 3162
rect 40114 3110 40116 3162
rect 40060 3108 40116 3110
rect 41132 4114 41188 4116
rect 41132 4062 41134 4114
rect 41134 4062 41186 4114
rect 41186 4062 41188 4114
rect 41132 4060 41188 4062
rect 40908 924 40964 980
rect 41020 3388 41076 3444
rect 41468 10444 41524 10500
rect 41916 11228 41972 11284
rect 41692 9660 41748 9716
rect 41356 8316 41412 8372
rect 41356 7868 41412 7924
rect 41804 9042 41860 9044
rect 41804 8990 41806 9042
rect 41806 8990 41858 9042
rect 41858 8990 41860 9042
rect 41804 8988 41860 8990
rect 41580 8652 41636 8708
rect 41580 7698 41636 7700
rect 41580 7646 41582 7698
rect 41582 7646 41634 7698
rect 41634 7646 41636 7698
rect 41580 7644 41636 7646
rect 41692 7420 41748 7476
rect 41356 5180 41412 5236
rect 41580 6578 41636 6580
rect 41580 6526 41582 6578
rect 41582 6526 41634 6578
rect 41634 6526 41636 6578
rect 41580 6524 41636 6526
rect 42140 11170 42196 11172
rect 42140 11118 42142 11170
rect 42142 11118 42194 11170
rect 42194 11118 42196 11170
rect 42140 11116 42196 11118
rect 42028 10108 42084 10164
rect 42028 8764 42084 8820
rect 46060 13916 46116 13972
rect 43372 13468 43428 13524
rect 42364 12572 42420 12628
rect 42812 12572 42868 12628
rect 42476 12012 42532 12068
rect 43260 12236 43316 12292
rect 43148 11788 43204 11844
rect 42812 11116 42868 11172
rect 42476 10556 42532 10612
rect 42364 9772 42420 9828
rect 41804 6690 41860 6692
rect 41804 6638 41806 6690
rect 41806 6638 41858 6690
rect 41858 6638 41860 6690
rect 41804 6636 41860 6638
rect 42140 6636 42196 6692
rect 41468 4060 41524 4116
rect 42252 7756 42308 7812
rect 42700 8988 42756 9044
rect 42476 7644 42532 7700
rect 42700 7868 42756 7924
rect 42812 7532 42868 7588
rect 42364 7308 42420 7364
rect 42476 7084 42532 7140
rect 42588 6972 42644 7028
rect 42028 6466 42084 6468
rect 42028 6414 42030 6466
rect 42030 6414 42082 6466
rect 42082 6414 42084 6466
rect 42028 6412 42084 6414
rect 42252 6076 42308 6132
rect 42140 5628 42196 5684
rect 42252 5740 42308 5796
rect 41916 4284 41972 4340
rect 42028 4956 42084 5012
rect 41804 4172 41860 4228
rect 41916 3052 41972 3108
rect 42140 3164 42196 3220
rect 42476 6076 42532 6132
rect 42476 4898 42532 4900
rect 42476 4846 42478 4898
rect 42478 4846 42530 4898
rect 42530 4846 42532 4898
rect 42476 4844 42532 4846
rect 42476 4620 42532 4676
rect 42812 6690 42868 6692
rect 42812 6638 42814 6690
rect 42814 6638 42866 6690
rect 42866 6638 42868 6690
rect 42812 6636 42868 6638
rect 42812 6412 42868 6468
rect 44044 13020 44100 13076
rect 43932 12684 43988 12740
rect 44268 12348 44324 12404
rect 43148 9660 43204 9716
rect 43708 11116 43764 11172
rect 43708 10498 43764 10500
rect 43708 10446 43710 10498
rect 43710 10446 43762 10498
rect 43762 10446 43764 10498
rect 43708 10444 43764 10446
rect 43708 9660 43764 9716
rect 43372 9548 43428 9604
rect 43596 9100 43652 9156
rect 43484 8764 43540 8820
rect 43148 7308 43204 7364
rect 43036 7084 43092 7140
rect 42924 5404 42980 5460
rect 42812 4620 42868 4676
rect 42700 4172 42756 4228
rect 42476 3388 42532 3444
rect 42700 2940 42756 2996
rect 42364 2828 42420 2884
rect 43148 5628 43204 5684
rect 43036 4060 43092 4116
rect 42252 1260 42308 1316
rect 42028 1148 42084 1204
rect 43148 3724 43204 3780
rect 43148 3388 43204 3444
rect 43372 6412 43428 6468
rect 43820 8540 43876 8596
rect 43596 7308 43652 7364
rect 43820 7756 43876 7812
rect 43596 5628 43652 5684
rect 43708 6524 43764 6580
rect 44380 11228 44436 11284
rect 44380 9602 44436 9604
rect 44380 9550 44382 9602
rect 44382 9550 44434 9602
rect 44434 9550 44436 9602
rect 44380 9548 44436 9550
rect 44380 8652 44436 8708
rect 44156 8092 44212 8148
rect 44044 7980 44100 8036
rect 44044 7308 44100 7364
rect 44268 7756 44324 7812
rect 44268 6972 44324 7028
rect 44380 7420 44436 7476
rect 44044 6748 44100 6804
rect 44156 6636 44212 6692
rect 44044 6412 44100 6468
rect 43820 6076 43876 6132
rect 43932 6188 43988 6244
rect 43372 3612 43428 3668
rect 43708 5180 43764 5236
rect 43596 4620 43652 4676
rect 43708 4898 43764 4900
rect 43708 4846 43710 4898
rect 43710 4846 43762 4898
rect 43762 4846 43764 4898
rect 43708 4844 43764 4846
rect 43932 4898 43988 4900
rect 43932 4846 43934 4898
rect 43934 4846 43986 4898
rect 43986 4846 43988 4898
rect 43932 4844 43988 4846
rect 43820 4620 43876 4676
rect 44380 6188 44436 6244
rect 44380 6018 44436 6020
rect 44380 5966 44382 6018
rect 44382 5966 44434 6018
rect 44434 5966 44436 6018
rect 44380 5964 44436 5966
rect 44268 4844 44324 4900
rect 44380 5628 44436 5684
rect 44156 4732 44212 4788
rect 43708 4284 43764 4340
rect 43820 4172 43876 4228
rect 43708 3948 43764 4004
rect 44044 4338 44100 4340
rect 44044 4286 44046 4338
rect 44046 4286 44098 4338
rect 44098 4286 44100 4338
rect 44044 4284 44100 4286
rect 44380 4060 44436 4116
rect 44156 3500 44212 3556
rect 44940 11170 44996 11172
rect 44940 11118 44942 11170
rect 44942 11118 44994 11170
rect 44994 11118 44996 11170
rect 44940 11116 44996 11118
rect 44828 10444 44884 10500
rect 44828 10108 44884 10164
rect 44716 8930 44772 8932
rect 44716 8878 44718 8930
rect 44718 8878 44770 8930
rect 44770 8878 44772 8930
rect 44716 8876 44772 8878
rect 45164 10444 45220 10500
rect 45612 12290 45668 12292
rect 45612 12238 45614 12290
rect 45614 12238 45666 12290
rect 45666 12238 45668 12290
rect 45612 12236 45668 12238
rect 45724 11340 45780 11396
rect 45612 11116 45668 11172
rect 45388 10220 45444 10276
rect 45388 9884 45444 9940
rect 45948 11228 46004 11284
rect 44940 8652 44996 8708
rect 45276 8540 45332 8596
rect 44604 7980 44660 8036
rect 44716 7644 44772 7700
rect 44604 6524 44660 6580
rect 44716 6972 44772 7028
rect 44604 6076 44660 6132
rect 45164 8204 45220 8260
rect 45052 8034 45108 8036
rect 45052 7982 45054 8034
rect 45054 7982 45106 8034
rect 45106 7982 45108 8034
rect 45052 7980 45108 7982
rect 45052 7644 45108 7700
rect 44828 6076 44884 6132
rect 44940 5852 44996 5908
rect 44828 5794 44884 5796
rect 44828 5742 44830 5794
rect 44830 5742 44882 5794
rect 44882 5742 44884 5794
rect 44828 5740 44884 5742
rect 44828 4956 44884 5012
rect 44828 4620 44884 4676
rect 44716 3724 44772 3780
rect 44492 3500 44548 3556
rect 44044 3276 44100 3332
rect 43372 1596 43428 1652
rect 43148 924 43204 980
rect 44940 3612 44996 3668
rect 44828 3388 44884 3444
rect 45836 9100 45892 9156
rect 45836 8930 45892 8932
rect 45836 8878 45838 8930
rect 45838 8878 45890 8930
rect 45890 8878 45892 8930
rect 45836 8876 45892 8878
rect 45836 8146 45892 8148
rect 45836 8094 45838 8146
rect 45838 8094 45890 8146
rect 45890 8094 45892 8146
rect 45836 8092 45892 8094
rect 45724 7586 45780 7588
rect 45724 7534 45726 7586
rect 45726 7534 45778 7586
rect 45778 7534 45780 7586
rect 45724 7532 45780 7534
rect 45500 6524 45556 6580
rect 45724 6300 45780 6356
rect 45836 5740 45892 5796
rect 45276 5404 45332 5460
rect 45612 5404 45668 5460
rect 45276 4620 45332 4676
rect 45388 4844 45444 4900
rect 45388 4508 45444 4564
rect 45276 3948 45332 4004
rect 45052 3276 45108 3332
rect 44940 3164 44996 3220
rect 45276 3052 45332 3108
rect 45388 3836 45444 3892
rect 44716 2940 44772 2996
rect 44268 1596 44324 1652
rect 43820 1260 43876 1316
rect 45052 2492 45108 2548
rect 46172 13074 46228 13076
rect 46172 13022 46174 13074
rect 46174 13022 46226 13074
rect 46226 13022 46228 13074
rect 46172 13020 46228 13022
rect 46172 12460 46228 12516
rect 46172 11340 46228 11396
rect 46396 12124 46452 12180
rect 46060 5516 46116 5572
rect 45612 5010 45668 5012
rect 45612 4958 45614 5010
rect 45614 4958 45666 5010
rect 45666 4958 45668 5010
rect 45612 4956 45668 4958
rect 45948 4732 46004 4788
rect 45948 4508 46004 4564
rect 45500 3276 45556 3332
rect 45500 3052 45556 3108
rect 46172 10892 46228 10948
rect 48076 12572 48132 12628
rect 47516 11564 47572 11620
rect 46956 11116 47012 11172
rect 46396 7980 46452 8036
rect 46396 7644 46452 7700
rect 46956 10332 47012 10388
rect 47068 10108 47124 10164
rect 47068 9772 47124 9828
rect 46732 8204 46788 8260
rect 46844 8316 46900 8372
rect 46620 8092 46676 8148
rect 46508 6972 46564 7028
rect 46396 6636 46452 6692
rect 46396 6300 46452 6356
rect 47180 8652 47236 8708
rect 47404 8876 47460 8932
rect 47068 7644 47124 7700
rect 47180 8092 47236 8148
rect 47292 7532 47348 7588
rect 47068 6412 47124 6468
rect 46396 6076 46452 6132
rect 46732 6076 46788 6132
rect 46508 5852 46564 5908
rect 46732 5852 46788 5908
rect 46284 5404 46340 5460
rect 46172 4396 46228 4452
rect 46172 4060 46228 4116
rect 45836 3330 45892 3332
rect 45836 3278 45838 3330
rect 45838 3278 45890 3330
rect 45890 3278 45892 3330
rect 45836 3276 45892 3278
rect 46060 3612 46116 3668
rect 46284 3442 46340 3444
rect 46284 3390 46286 3442
rect 46286 3390 46338 3442
rect 46338 3390 46340 3442
rect 46284 3388 46340 3390
rect 46172 3276 46228 3332
rect 46844 5628 46900 5684
rect 46956 6300 47012 6356
rect 46732 5404 46788 5460
rect 46620 5180 46676 5236
rect 47180 6076 47236 6132
rect 46844 5234 46900 5236
rect 46844 5182 46846 5234
rect 46846 5182 46898 5234
rect 46898 5182 46900 5234
rect 46844 5180 46900 5182
rect 46620 4620 46676 4676
rect 46844 4508 46900 4564
rect 46620 4396 46676 4452
rect 46844 4284 46900 4340
rect 47180 4284 47236 4340
rect 46732 3948 46788 4004
rect 47068 3948 47124 4004
rect 46732 3276 46788 3332
rect 46620 3052 46676 3108
rect 45612 924 45668 980
rect 45836 978 45892 980
rect 45836 926 45838 978
rect 45838 926 45890 978
rect 45890 926 45892 978
rect 45836 924 45892 926
rect 46956 3388 47012 3444
rect 46844 1372 46900 1428
rect 47628 11116 47684 11172
rect 47628 10332 47684 10388
rect 48076 10556 48132 10612
rect 47628 9324 47684 9380
rect 48076 9660 48132 9716
rect 47740 9154 47796 9156
rect 47740 9102 47742 9154
rect 47742 9102 47794 9154
rect 47794 9102 47796 9154
rect 47740 9100 47796 9102
rect 47852 8652 47908 8708
rect 47964 8540 48020 8596
rect 47852 8092 47908 8148
rect 47628 7420 47684 7476
rect 47516 6860 47572 6916
rect 47516 6188 47572 6244
rect 47628 5964 47684 6020
rect 47404 3948 47460 4004
rect 47404 3724 47460 3780
rect 48188 9100 48244 9156
rect 47852 6860 47908 6916
rect 48076 7698 48132 7700
rect 48076 7646 48078 7698
rect 48078 7646 48130 7698
rect 48130 7646 48132 7698
rect 48076 7644 48132 7646
rect 49512 16490 49568 16492
rect 49512 16438 49514 16490
rect 49514 16438 49566 16490
rect 49566 16438 49568 16490
rect 49512 16436 49568 16438
rect 49616 16490 49672 16492
rect 49616 16438 49618 16490
rect 49618 16438 49670 16490
rect 49670 16438 49672 16490
rect 49616 16436 49672 16438
rect 49720 16490 49776 16492
rect 49720 16438 49722 16490
rect 49722 16438 49774 16490
rect 49774 16438 49776 16490
rect 49720 16436 49776 16438
rect 48524 15820 48580 15876
rect 48412 10444 48468 10500
rect 48412 9548 48468 9604
rect 48412 8316 48468 8372
rect 48188 7084 48244 7140
rect 47740 4620 47796 4676
rect 47628 3612 47684 3668
rect 47964 6188 48020 6244
rect 47964 4508 48020 4564
rect 48300 5964 48356 6020
rect 48188 5068 48244 5124
rect 48188 4620 48244 4676
rect 48076 3388 48132 3444
rect 51436 15484 51492 15540
rect 54236 15260 54292 15316
rect 49512 14922 49568 14924
rect 49512 14870 49514 14922
rect 49514 14870 49566 14922
rect 49566 14870 49568 14922
rect 49512 14868 49568 14870
rect 49616 14922 49672 14924
rect 49616 14870 49618 14922
rect 49618 14870 49670 14922
rect 49670 14870 49672 14922
rect 49616 14868 49672 14870
rect 49720 14922 49776 14924
rect 49720 14870 49722 14922
rect 49722 14870 49774 14922
rect 49774 14870 49776 14922
rect 49720 14868 49776 14870
rect 49512 13354 49568 13356
rect 49512 13302 49514 13354
rect 49514 13302 49566 13354
rect 49566 13302 49568 13354
rect 49512 13300 49568 13302
rect 49616 13354 49672 13356
rect 49616 13302 49618 13354
rect 49618 13302 49670 13354
rect 49670 13302 49672 13354
rect 49616 13300 49672 13302
rect 49720 13354 49776 13356
rect 49720 13302 49722 13354
rect 49722 13302 49774 13354
rect 49774 13302 49776 13354
rect 49720 13300 49776 13302
rect 48748 11788 48804 11844
rect 48860 11900 48916 11956
rect 48636 11116 48692 11172
rect 48748 11228 48804 11284
rect 48748 10332 48804 10388
rect 48860 9548 48916 9604
rect 49512 11786 49568 11788
rect 49512 11734 49514 11786
rect 49514 11734 49566 11786
rect 49566 11734 49568 11786
rect 49512 11732 49568 11734
rect 49616 11786 49672 11788
rect 49616 11734 49618 11786
rect 49618 11734 49670 11786
rect 49670 11734 49672 11786
rect 49616 11732 49672 11734
rect 49720 11786 49776 11788
rect 49720 11734 49722 11786
rect 49722 11734 49774 11786
rect 49774 11734 49776 11786
rect 49720 11732 49776 11734
rect 50316 12066 50372 12068
rect 50316 12014 50318 12066
rect 50318 12014 50370 12066
rect 50370 12014 50372 12066
rect 50316 12012 50372 12014
rect 49756 10498 49812 10500
rect 49756 10446 49758 10498
rect 49758 10446 49810 10498
rect 49810 10446 49812 10498
rect 49756 10444 49812 10446
rect 49196 10108 49252 10164
rect 49308 10332 49364 10388
rect 49512 10218 49568 10220
rect 49512 10166 49514 10218
rect 49514 10166 49566 10218
rect 49566 10166 49568 10218
rect 49512 10164 49568 10166
rect 49616 10218 49672 10220
rect 49616 10166 49618 10218
rect 49618 10166 49670 10218
rect 49670 10166 49672 10218
rect 49616 10164 49672 10166
rect 49720 10218 49776 10220
rect 49720 10166 49722 10218
rect 49722 10166 49774 10218
rect 49774 10166 49776 10218
rect 49720 10164 49776 10166
rect 49980 9884 50036 9940
rect 50092 11506 50148 11508
rect 50092 11454 50094 11506
rect 50094 11454 50146 11506
rect 50146 11454 50148 11506
rect 50092 11452 50148 11454
rect 48972 9436 49028 9492
rect 49308 9436 49364 9492
rect 48860 9154 48916 9156
rect 48860 9102 48862 9154
rect 48862 9102 48914 9154
rect 48914 9102 48916 9154
rect 48860 9100 48916 9102
rect 48636 8540 48692 8596
rect 48972 8540 49028 8596
rect 48748 8316 48804 8372
rect 48636 7980 48692 8036
rect 48748 7586 48804 7588
rect 48748 7534 48750 7586
rect 48750 7534 48802 7586
rect 48802 7534 48804 7586
rect 48748 7532 48804 7534
rect 48636 7084 48692 7140
rect 48636 6524 48692 6580
rect 49420 8764 49476 8820
rect 49644 8988 49700 9044
rect 49644 8764 49700 8820
rect 49308 8540 49364 8596
rect 49512 8650 49568 8652
rect 49512 8598 49514 8650
rect 49514 8598 49566 8650
rect 49566 8598 49568 8650
rect 49512 8596 49568 8598
rect 49616 8650 49672 8652
rect 49616 8598 49618 8650
rect 49618 8598 49670 8650
rect 49670 8598 49672 8650
rect 49616 8596 49672 8598
rect 49720 8650 49776 8652
rect 49720 8598 49722 8650
rect 49722 8598 49774 8650
rect 49774 8598 49776 8650
rect 49720 8596 49776 8598
rect 50764 10722 50820 10724
rect 50764 10670 50766 10722
rect 50766 10670 50818 10722
rect 50818 10670 50820 10722
rect 50764 10668 50820 10670
rect 50540 10332 50596 10388
rect 50876 10444 50932 10500
rect 50428 9996 50484 10052
rect 49308 8316 49364 8372
rect 48972 7698 49028 7700
rect 48972 7646 48974 7698
rect 48974 7646 49026 7698
rect 49026 7646 49028 7698
rect 48972 7644 49028 7646
rect 49084 7474 49140 7476
rect 49084 7422 49086 7474
rect 49086 7422 49138 7474
rect 49138 7422 49140 7474
rect 49084 7420 49140 7422
rect 49980 8540 50036 8596
rect 50092 8316 50148 8372
rect 50204 8988 50260 9044
rect 49644 8146 49700 8148
rect 49644 8094 49646 8146
rect 49646 8094 49698 8146
rect 49698 8094 49700 8146
rect 49644 8092 49700 8094
rect 49532 7532 49588 7588
rect 49196 6524 49252 6580
rect 49196 6300 49252 6356
rect 48860 5906 48916 5908
rect 48860 5854 48862 5906
rect 48862 5854 48914 5906
rect 48914 5854 48916 5906
rect 48860 5852 48916 5854
rect 48972 5628 49028 5684
rect 48972 5180 49028 5236
rect 48748 3500 48804 3556
rect 49196 5852 49252 5908
rect 49196 5516 49252 5572
rect 49980 7980 50036 8036
rect 49756 7308 49812 7364
rect 49868 7532 49924 7588
rect 49512 7082 49568 7084
rect 49512 7030 49514 7082
rect 49514 7030 49566 7082
rect 49566 7030 49568 7082
rect 49512 7028 49568 7030
rect 49616 7082 49672 7084
rect 49616 7030 49618 7082
rect 49618 7030 49670 7082
rect 49670 7030 49672 7082
rect 49616 7028 49672 7030
rect 49720 7082 49776 7084
rect 49720 7030 49722 7082
rect 49722 7030 49774 7082
rect 49774 7030 49776 7082
rect 49720 7028 49776 7030
rect 49756 5628 49812 5684
rect 49512 5514 49568 5516
rect 49512 5462 49514 5514
rect 49514 5462 49566 5514
rect 49566 5462 49568 5514
rect 49512 5460 49568 5462
rect 49616 5514 49672 5516
rect 49616 5462 49618 5514
rect 49618 5462 49670 5514
rect 49670 5462 49672 5514
rect 49616 5460 49672 5462
rect 49720 5514 49776 5516
rect 49720 5462 49722 5514
rect 49722 5462 49774 5514
rect 49774 5462 49776 5514
rect 49720 5460 49776 5462
rect 49644 5292 49700 5348
rect 49756 4956 49812 5012
rect 49420 4172 49476 4228
rect 49512 3946 49568 3948
rect 49512 3894 49514 3946
rect 49514 3894 49566 3946
rect 49566 3894 49568 3946
rect 49512 3892 49568 3894
rect 49616 3946 49672 3948
rect 49616 3894 49618 3946
rect 49618 3894 49670 3946
rect 49670 3894 49672 3946
rect 49616 3892 49672 3894
rect 49720 3946 49776 3948
rect 49720 3894 49722 3946
rect 49722 3894 49774 3946
rect 49774 3894 49776 3946
rect 49720 3892 49776 3894
rect 50092 7420 50148 7476
rect 50540 9436 50596 9492
rect 50652 9100 50708 9156
rect 50764 8988 50820 9044
rect 50764 8652 50820 8708
rect 50428 8258 50484 8260
rect 50428 8206 50430 8258
rect 50430 8206 50482 8258
rect 50482 8206 50484 8258
rect 50428 8204 50484 8206
rect 50204 5516 50260 5572
rect 50316 5292 50372 5348
rect 50316 4844 50372 4900
rect 49308 1484 49364 1540
rect 50204 3330 50260 3332
rect 50204 3278 50206 3330
rect 50206 3278 50258 3330
rect 50258 3278 50260 3330
rect 50204 3276 50260 3278
rect 50652 7644 50708 7700
rect 50764 7308 50820 7364
rect 50540 3836 50596 3892
rect 50652 6636 50708 6692
rect 50428 3554 50484 3556
rect 50428 3502 50430 3554
rect 50430 3502 50482 3554
rect 50482 3502 50484 3554
rect 50428 3500 50484 3502
rect 50316 2828 50372 2884
rect 51548 11282 51604 11284
rect 51548 11230 51550 11282
rect 51550 11230 51602 11282
rect 51602 11230 51604 11282
rect 51548 11228 51604 11230
rect 51548 9996 51604 10052
rect 51324 9884 51380 9940
rect 50988 9212 51044 9268
rect 51100 8764 51156 8820
rect 51100 8428 51156 8484
rect 50988 6636 51044 6692
rect 50204 1708 50260 1764
rect 50204 1036 50260 1092
rect 50988 6466 51044 6468
rect 50988 6414 50990 6466
rect 50990 6414 51042 6466
rect 51042 6414 51044 6466
rect 50988 6412 51044 6414
rect 50988 6188 51044 6244
rect 50764 2716 50820 2772
rect 50876 5628 50932 5684
rect 51100 6076 51156 6132
rect 51100 4620 51156 4676
rect 51548 8876 51604 8932
rect 51548 8540 51604 8596
rect 51324 7980 51380 8036
rect 53228 13132 53284 13188
rect 52332 11004 52388 11060
rect 51324 7308 51380 7364
rect 51996 10108 52052 10164
rect 51996 9660 52052 9716
rect 52220 8930 52276 8932
rect 52220 8878 52222 8930
rect 52222 8878 52274 8930
rect 52274 8878 52276 8930
rect 52220 8876 52276 8878
rect 52220 8428 52276 8484
rect 51884 8258 51940 8260
rect 51884 8206 51886 8258
rect 51886 8206 51938 8258
rect 51938 8206 51940 8258
rect 51884 8204 51940 8206
rect 51548 6636 51604 6692
rect 51884 7980 51940 8036
rect 51772 7308 51828 7364
rect 51772 6412 51828 6468
rect 51660 5516 51716 5572
rect 51996 7644 52052 7700
rect 51884 6188 51940 6244
rect 51884 5794 51940 5796
rect 51884 5742 51886 5794
rect 51886 5742 51938 5794
rect 51938 5742 51940 5794
rect 51884 5740 51940 5742
rect 52108 6802 52164 6804
rect 52108 6750 52110 6802
rect 52110 6750 52162 6802
rect 52162 6750 52164 6802
rect 52108 6748 52164 6750
rect 51996 5516 52052 5572
rect 51772 5180 51828 5236
rect 51996 5292 52052 5348
rect 51548 3836 51604 3892
rect 51548 3330 51604 3332
rect 51548 3278 51550 3330
rect 51550 3278 51602 3330
rect 51602 3278 51604 3330
rect 51548 3276 51604 3278
rect 51436 1820 51492 1876
rect 52332 8316 52388 8372
rect 52556 10498 52612 10500
rect 52556 10446 52558 10498
rect 52558 10446 52610 10498
rect 52610 10446 52612 10498
rect 52556 10444 52612 10446
rect 53004 10108 53060 10164
rect 53004 9772 53060 9828
rect 52668 9602 52724 9604
rect 52668 9550 52670 9602
rect 52670 9550 52722 9602
rect 52722 9550 52724 9602
rect 52668 9548 52724 9550
rect 52556 9324 52612 9380
rect 52892 9436 52948 9492
rect 52556 7980 52612 8036
rect 52332 6860 52388 6916
rect 52220 5292 52276 5348
rect 53116 9212 53172 9268
rect 53004 8092 53060 8148
rect 53788 10892 53844 10948
rect 53564 8652 53620 8708
rect 53676 9548 53732 9604
rect 53228 7644 53284 7700
rect 53228 5906 53284 5908
rect 53228 5854 53230 5906
rect 53230 5854 53282 5906
rect 53282 5854 53284 5906
rect 53228 5852 53284 5854
rect 52780 5516 52836 5572
rect 52220 5068 52276 5124
rect 52444 4732 52500 4788
rect 52332 4620 52388 4676
rect 52220 3666 52276 3668
rect 52220 3614 52222 3666
rect 52222 3614 52274 3666
rect 52274 3614 52276 3666
rect 52220 3612 52276 3614
rect 52108 2940 52164 2996
rect 51884 2380 51940 2436
rect 52668 4620 52724 4676
rect 52780 5292 52836 5348
rect 52668 4284 52724 4340
rect 52556 4226 52612 4228
rect 52556 4174 52558 4226
rect 52558 4174 52610 4226
rect 52610 4174 52612 4226
rect 52556 4172 52612 4174
rect 52556 3666 52612 3668
rect 52556 3614 52558 3666
rect 52558 3614 52610 3666
rect 52610 3614 52612 3666
rect 52556 3612 52612 3614
rect 53452 5628 53508 5684
rect 53452 5234 53508 5236
rect 53452 5182 53454 5234
rect 53454 5182 53506 5234
rect 53506 5182 53508 5234
rect 53452 5180 53508 5182
rect 53004 4284 53060 4340
rect 53116 4956 53172 5012
rect 53004 3948 53060 4004
rect 53340 4508 53396 4564
rect 53340 4060 53396 4116
rect 53564 4114 53620 4116
rect 53564 4062 53566 4114
rect 53566 4062 53618 4114
rect 53618 4062 53620 4114
rect 53564 4060 53620 4062
rect 54012 10498 54068 10500
rect 54012 10446 54014 10498
rect 54014 10446 54066 10498
rect 54066 10446 54068 10498
rect 54012 10444 54068 10446
rect 53900 9042 53956 9044
rect 53900 8990 53902 9042
rect 53902 8990 53954 9042
rect 53954 8990 53956 9042
rect 53900 8988 53956 8990
rect 53788 8370 53844 8372
rect 53788 8318 53790 8370
rect 53790 8318 53842 8370
rect 53842 8318 53844 8370
rect 53788 8316 53844 8318
rect 53676 3948 53732 4004
rect 53788 7980 53844 8036
rect 53676 3666 53732 3668
rect 53676 3614 53678 3666
rect 53678 3614 53730 3666
rect 53730 3614 53732 3666
rect 53676 3612 53732 3614
rect 53676 3388 53732 3444
rect 53340 2604 53396 2660
rect 53900 6636 53956 6692
rect 68832 18058 68888 18060
rect 68832 18006 68834 18058
rect 68834 18006 68886 18058
rect 68886 18006 68888 18058
rect 68832 18004 68888 18006
rect 68936 18058 68992 18060
rect 68936 18006 68938 18058
rect 68938 18006 68990 18058
rect 68990 18006 68992 18058
rect 68936 18004 68992 18006
rect 69040 18058 69096 18060
rect 69040 18006 69042 18058
rect 69042 18006 69094 18058
rect 69094 18006 69096 18058
rect 69040 18004 69096 18006
rect 67116 17388 67172 17444
rect 59172 17274 59228 17276
rect 59172 17222 59174 17274
rect 59174 17222 59226 17274
rect 59226 17222 59228 17274
rect 59172 17220 59228 17222
rect 59276 17274 59332 17276
rect 59276 17222 59278 17274
rect 59278 17222 59330 17274
rect 59330 17222 59332 17274
rect 59276 17220 59332 17222
rect 59380 17274 59436 17276
rect 59380 17222 59382 17274
rect 59382 17222 59434 17274
rect 59434 17222 59436 17274
rect 59380 17220 59436 17222
rect 56028 16940 56084 16996
rect 59172 15706 59228 15708
rect 59172 15654 59174 15706
rect 59174 15654 59226 15706
rect 59226 15654 59228 15706
rect 59172 15652 59228 15654
rect 59276 15706 59332 15708
rect 59276 15654 59278 15706
rect 59278 15654 59330 15706
rect 59330 15654 59332 15706
rect 59276 15652 59332 15654
rect 59380 15706 59436 15708
rect 59380 15654 59382 15706
rect 59382 15654 59434 15706
rect 59434 15654 59436 15706
rect 59380 15652 59436 15654
rect 57372 15372 57428 15428
rect 55692 13580 55748 13636
rect 54348 8930 54404 8932
rect 54348 8878 54350 8930
rect 54350 8878 54402 8930
rect 54402 8878 54404 8930
rect 54348 8876 54404 8878
rect 54348 7698 54404 7700
rect 54348 7646 54350 7698
rect 54350 7646 54402 7698
rect 54402 7646 54404 7698
rect 54348 7644 54404 7646
rect 54684 10444 54740 10500
rect 54684 9772 54740 9828
rect 54572 8540 54628 8596
rect 54012 4732 54068 4788
rect 54460 6860 54516 6916
rect 54124 4508 54180 4564
rect 54236 5740 54292 5796
rect 53900 4338 53956 4340
rect 53900 4286 53902 4338
rect 53902 4286 53954 4338
rect 53954 4286 53956 4338
rect 53900 4284 53956 4286
rect 54236 4060 54292 4116
rect 54348 5516 54404 5572
rect 54908 10444 54964 10500
rect 54796 8204 54852 8260
rect 54796 7698 54852 7700
rect 54796 7646 54798 7698
rect 54798 7646 54850 7698
rect 54850 7646 54852 7698
rect 54796 7644 54852 7646
rect 54684 5740 54740 5796
rect 54572 3612 54628 3668
rect 54684 5180 54740 5236
rect 54796 4844 54852 4900
rect 55020 9602 55076 9604
rect 55020 9550 55022 9602
rect 55022 9550 55074 9602
rect 55074 9550 55076 9602
rect 55020 9548 55076 9550
rect 55468 9154 55524 9156
rect 55468 9102 55470 9154
rect 55470 9102 55522 9154
rect 55522 9102 55524 9154
rect 55468 9100 55524 9102
rect 55356 8988 55412 9044
rect 55244 8092 55300 8148
rect 55468 7698 55524 7700
rect 55468 7646 55470 7698
rect 55470 7646 55522 7698
rect 55522 7646 55524 7698
rect 55468 7644 55524 7646
rect 54908 4732 54964 4788
rect 54908 4284 54964 4340
rect 55244 5740 55300 5796
rect 56252 13468 56308 13524
rect 56140 8876 56196 8932
rect 55804 8204 55860 8260
rect 56028 8092 56084 8148
rect 55916 8034 55972 8036
rect 55916 7982 55918 8034
rect 55918 7982 55970 8034
rect 55970 7982 55972 8034
rect 55916 7980 55972 7982
rect 55804 7868 55860 7924
rect 55804 7420 55860 7476
rect 56028 6972 56084 7028
rect 55916 5794 55972 5796
rect 55916 5742 55918 5794
rect 55918 5742 55970 5794
rect 55970 5742 55972 5794
rect 55916 5740 55972 5742
rect 55916 5516 55972 5572
rect 55692 5292 55748 5348
rect 55468 4956 55524 5012
rect 55356 4732 55412 4788
rect 55020 4114 55076 4116
rect 55020 4062 55022 4114
rect 55022 4062 55074 4114
rect 55074 4062 55076 4114
rect 55020 4060 55076 4062
rect 55020 3836 55076 3892
rect 56028 5404 56084 5460
rect 56364 6860 56420 6916
rect 56364 5740 56420 5796
rect 56140 5068 56196 5124
rect 55468 4620 55524 4676
rect 56140 4508 56196 4564
rect 56252 4732 56308 4788
rect 55468 4060 55524 4116
rect 55356 3388 55412 3444
rect 55692 2716 55748 2772
rect 55916 3666 55972 3668
rect 55916 3614 55918 3666
rect 55918 3614 55970 3666
rect 55970 3614 55972 3666
rect 55916 3612 55972 3614
rect 56588 8876 56644 8932
rect 57148 8930 57204 8932
rect 57148 8878 57150 8930
rect 57150 8878 57202 8930
rect 57202 8878 57204 8930
rect 57148 8876 57204 8878
rect 56700 8652 56756 8708
rect 56588 7698 56644 7700
rect 56588 7646 56590 7698
rect 56590 7646 56642 7698
rect 56642 7646 56644 7698
rect 56588 7644 56644 7646
rect 56700 7532 56756 7588
rect 56588 6972 56644 7028
rect 56924 7586 56980 7588
rect 56924 7534 56926 7586
rect 56926 7534 56978 7586
rect 56978 7534 56980 7586
rect 56924 7532 56980 7534
rect 57036 7420 57092 7476
rect 56924 6860 56980 6916
rect 56924 4844 56980 4900
rect 56924 3836 56980 3892
rect 55692 924 55748 980
rect 55804 1708 55860 1764
rect 56476 3724 56532 3780
rect 56140 1596 56196 1652
rect 56028 1260 56084 1316
rect 59172 14138 59228 14140
rect 59172 14086 59174 14138
rect 59174 14086 59226 14138
rect 59226 14086 59228 14138
rect 59172 14084 59228 14086
rect 59276 14138 59332 14140
rect 59276 14086 59278 14138
rect 59278 14086 59330 14138
rect 59330 14086 59332 14138
rect 59276 14084 59332 14086
rect 59380 14138 59436 14140
rect 59380 14086 59382 14138
rect 59382 14086 59434 14138
rect 59434 14086 59436 14138
rect 59380 14084 59436 14086
rect 59172 12570 59228 12572
rect 59172 12518 59174 12570
rect 59174 12518 59226 12570
rect 59226 12518 59228 12570
rect 59172 12516 59228 12518
rect 59276 12570 59332 12572
rect 59276 12518 59278 12570
rect 59278 12518 59330 12570
rect 59330 12518 59332 12570
rect 59276 12516 59332 12518
rect 59380 12570 59436 12572
rect 59380 12518 59382 12570
rect 59382 12518 59434 12570
rect 59434 12518 59436 12570
rect 59380 12516 59436 12518
rect 58828 12124 58884 12180
rect 58044 11900 58100 11956
rect 57708 11788 57764 11844
rect 57484 10108 57540 10164
rect 57260 7084 57316 7140
rect 57484 7474 57540 7476
rect 57484 7422 57486 7474
rect 57486 7422 57538 7474
rect 57538 7422 57540 7474
rect 57484 7420 57540 7422
rect 57260 6018 57316 6020
rect 57260 5966 57262 6018
rect 57262 5966 57314 6018
rect 57314 5966 57316 6018
rect 57260 5964 57316 5966
rect 57260 3836 57316 3892
rect 57148 3724 57204 3780
rect 57820 8876 57876 8932
rect 57932 7196 57988 7252
rect 57708 5516 57764 5572
rect 57708 4844 57764 4900
rect 58268 10556 58324 10612
rect 58156 10220 58212 10276
rect 57932 4732 57988 4788
rect 57484 4396 57540 4452
rect 57932 4508 57988 4564
rect 57036 3612 57092 3668
rect 56812 3052 56868 3108
rect 56700 2716 56756 2772
rect 57820 3724 57876 3780
rect 57596 3666 57652 3668
rect 57596 3614 57598 3666
rect 57598 3614 57650 3666
rect 57650 3614 57652 3666
rect 57596 3612 57652 3614
rect 57484 3164 57540 3220
rect 57372 2268 57428 2324
rect 58716 9548 58772 9604
rect 58492 8316 58548 8372
rect 66556 11788 66612 11844
rect 59052 11564 59108 11620
rect 58940 9548 58996 9604
rect 59172 11002 59228 11004
rect 59172 10950 59174 11002
rect 59174 10950 59226 11002
rect 59226 10950 59228 11002
rect 59172 10948 59228 10950
rect 59276 11002 59332 11004
rect 59276 10950 59278 11002
rect 59278 10950 59330 11002
rect 59330 10950 59332 11002
rect 59276 10948 59332 10950
rect 59380 11002 59436 11004
rect 59380 10950 59382 11002
rect 59382 10950 59434 11002
rect 59434 10950 59436 11002
rect 59380 10948 59436 10950
rect 60844 10892 60900 10948
rect 59500 10780 59556 10836
rect 59172 9434 59228 9436
rect 59172 9382 59174 9434
rect 59174 9382 59226 9434
rect 59226 9382 59228 9434
rect 59172 9380 59228 9382
rect 59276 9434 59332 9436
rect 59276 9382 59278 9434
rect 59278 9382 59330 9434
rect 59330 9382 59332 9434
rect 59276 9380 59332 9382
rect 59380 9434 59436 9436
rect 59380 9382 59382 9434
rect 59382 9382 59434 9434
rect 59434 9382 59436 9434
rect 59380 9380 59436 9382
rect 59052 8764 59108 8820
rect 60172 9548 60228 9604
rect 62076 10780 62132 10836
rect 61180 9772 61236 9828
rect 59724 8652 59780 8708
rect 60060 8764 60116 8820
rect 58380 7586 58436 7588
rect 58380 7534 58382 7586
rect 58382 7534 58434 7586
rect 58434 7534 58436 7586
rect 58380 7532 58436 7534
rect 58492 7362 58548 7364
rect 58492 7310 58494 7362
rect 58494 7310 58546 7362
rect 58546 7310 58548 7362
rect 58492 7308 58548 7310
rect 58380 7196 58436 7252
rect 59724 8204 59780 8260
rect 59948 8428 60004 8484
rect 58940 7756 58996 7812
rect 59172 7866 59228 7868
rect 59172 7814 59174 7866
rect 59174 7814 59226 7866
rect 59226 7814 59228 7866
rect 59172 7812 59228 7814
rect 59276 7866 59332 7868
rect 59276 7814 59278 7866
rect 59278 7814 59330 7866
rect 59330 7814 59332 7866
rect 59276 7812 59332 7814
rect 59380 7866 59436 7868
rect 59380 7814 59382 7866
rect 59382 7814 59434 7866
rect 59434 7814 59436 7866
rect 59380 7812 59436 7814
rect 59276 7586 59332 7588
rect 59276 7534 59278 7586
rect 59278 7534 59330 7586
rect 59330 7534 59332 7586
rect 59276 7532 59332 7534
rect 59052 7250 59108 7252
rect 59052 7198 59054 7250
rect 59054 7198 59106 7250
rect 59106 7198 59108 7250
rect 59052 7196 59108 7198
rect 59276 7308 59332 7364
rect 59276 6748 59332 6804
rect 58940 6690 58996 6692
rect 58940 6638 58942 6690
rect 58942 6638 58994 6690
rect 58994 6638 58996 6690
rect 58940 6636 58996 6638
rect 58268 5964 58324 6020
rect 59724 7084 59780 7140
rect 59612 6972 59668 7028
rect 58380 6412 58436 6468
rect 58604 6076 58660 6132
rect 58380 5628 58436 5684
rect 58492 5852 58548 5908
rect 58044 2492 58100 2548
rect 58828 5964 58884 6020
rect 59172 6298 59228 6300
rect 59172 6246 59174 6298
rect 59174 6246 59226 6298
rect 59226 6246 59228 6298
rect 59172 6244 59228 6246
rect 59276 6298 59332 6300
rect 59276 6246 59278 6298
rect 59278 6246 59330 6298
rect 59330 6246 59332 6298
rect 59276 6244 59332 6246
rect 59380 6298 59436 6300
rect 59380 6246 59382 6298
rect 59382 6246 59434 6298
rect 59434 6246 59436 6298
rect 59380 6244 59436 6246
rect 59612 6300 59668 6356
rect 59724 6188 59780 6244
rect 58716 5180 58772 5236
rect 58940 5628 58996 5684
rect 58716 4844 58772 4900
rect 58716 3388 58772 3444
rect 59500 5906 59556 5908
rect 59500 5854 59502 5906
rect 59502 5854 59554 5906
rect 59554 5854 59556 5906
rect 59500 5852 59556 5854
rect 59500 5628 59556 5684
rect 59388 4844 59444 4900
rect 59172 4730 59228 4732
rect 59172 4678 59174 4730
rect 59174 4678 59226 4730
rect 59226 4678 59228 4730
rect 59172 4676 59228 4678
rect 59276 4730 59332 4732
rect 59276 4678 59278 4730
rect 59278 4678 59330 4730
rect 59330 4678 59332 4730
rect 59276 4676 59332 4678
rect 59380 4730 59436 4732
rect 59380 4678 59382 4730
rect 59382 4678 59434 4730
rect 59434 4678 59436 4730
rect 59380 4676 59436 4678
rect 59388 4172 59444 4228
rect 59052 3724 59108 3780
rect 59164 4060 59220 4116
rect 58940 3276 58996 3332
rect 59724 4620 59780 4676
rect 59172 3162 59228 3164
rect 59172 3110 59174 3162
rect 59174 3110 59226 3162
rect 59226 3110 59228 3162
rect 59172 3108 59228 3110
rect 59276 3162 59332 3164
rect 59276 3110 59278 3162
rect 59278 3110 59330 3162
rect 59330 3110 59332 3162
rect 59276 3108 59332 3110
rect 59380 3162 59436 3164
rect 59380 3110 59382 3162
rect 59382 3110 59434 3162
rect 59434 3110 59436 3162
rect 59380 3108 59436 3110
rect 59724 3500 59780 3556
rect 59948 7308 60004 7364
rect 59948 6972 60004 7028
rect 60060 6748 60116 6804
rect 59948 6636 60004 6692
rect 60172 5964 60228 6020
rect 60396 8652 60452 8708
rect 60396 5964 60452 6020
rect 60396 5794 60452 5796
rect 60396 5742 60398 5794
rect 60398 5742 60450 5794
rect 60450 5742 60452 5794
rect 60396 5740 60452 5742
rect 60060 5628 60116 5684
rect 59948 5404 60004 5460
rect 60284 5404 60340 5460
rect 59948 4732 60004 4788
rect 59612 2940 59668 2996
rect 59052 1148 59108 1204
rect 59836 3164 59892 3220
rect 60172 3554 60228 3556
rect 60172 3502 60174 3554
rect 60174 3502 60226 3554
rect 60226 3502 60228 3554
rect 60172 3500 60228 3502
rect 60396 2940 60452 2996
rect 60060 2828 60116 2884
rect 60732 8764 60788 8820
rect 60732 8092 60788 8148
rect 60732 7868 60788 7924
rect 61292 9660 61348 9716
rect 61292 8652 61348 8708
rect 61404 8988 61460 9044
rect 61180 8428 61236 8484
rect 60844 7756 60900 7812
rect 60732 7644 60788 7700
rect 60732 6524 60788 6580
rect 60732 5628 60788 5684
rect 60620 5404 60676 5460
rect 60620 5234 60676 5236
rect 60620 5182 60622 5234
rect 60622 5182 60674 5234
rect 60674 5182 60676 5234
rect 60620 5180 60676 5182
rect 60620 3948 60676 4004
rect 60956 7196 61012 7252
rect 60956 6188 61012 6244
rect 61068 6972 61124 7028
rect 60956 5852 61012 5908
rect 61180 7756 61236 7812
rect 61068 5122 61124 5124
rect 61068 5070 61070 5122
rect 61070 5070 61122 5122
rect 61122 5070 61124 5122
rect 61068 5068 61124 5070
rect 61068 4172 61124 4228
rect 61180 3948 61236 4004
rect 61180 3724 61236 3780
rect 61740 8428 61796 8484
rect 61516 7532 61572 7588
rect 61740 7420 61796 7476
rect 61852 8204 61908 8260
rect 61516 7362 61572 7364
rect 61516 7310 61518 7362
rect 61518 7310 61570 7362
rect 61570 7310 61572 7362
rect 61516 7308 61572 7310
rect 61740 6972 61796 7028
rect 61516 6860 61572 6916
rect 61852 6524 61908 6580
rect 61740 6412 61796 6468
rect 61964 6300 62020 6356
rect 62748 10332 62804 10388
rect 62300 8876 62356 8932
rect 62300 8428 62356 8484
rect 62188 8204 62244 8260
rect 62188 7980 62244 8036
rect 62188 7644 62244 7700
rect 62188 7308 62244 7364
rect 62076 6076 62132 6132
rect 62188 7084 62244 7140
rect 62300 6748 62356 6804
rect 62524 9042 62580 9044
rect 62524 8990 62526 9042
rect 62526 8990 62578 9042
rect 62578 8990 62580 9042
rect 62524 8988 62580 8990
rect 62636 8428 62692 8484
rect 62524 8258 62580 8260
rect 62524 8206 62526 8258
rect 62526 8206 62578 8258
rect 62578 8206 62580 8258
rect 62524 8204 62580 8206
rect 62412 6524 62468 6580
rect 62524 7532 62580 7588
rect 62524 6412 62580 6468
rect 61740 5628 61796 5684
rect 61404 5180 61460 5236
rect 61516 5516 61572 5572
rect 62076 5404 62132 5460
rect 60732 3164 60788 3220
rect 60956 3276 61012 3332
rect 62076 3948 62132 4004
rect 61740 2940 61796 2996
rect 61852 3276 61908 3332
rect 61964 1708 62020 1764
rect 62524 6076 62580 6132
rect 62300 4732 62356 4788
rect 62412 4396 62468 4452
rect 63532 10108 63588 10164
rect 63084 9826 63140 9828
rect 63084 9774 63086 9826
rect 63086 9774 63138 9826
rect 63138 9774 63140 9826
rect 63084 9772 63140 9774
rect 62860 8876 62916 8932
rect 63196 8764 63252 8820
rect 63532 8428 63588 8484
rect 62860 7586 62916 7588
rect 62860 7534 62862 7586
rect 62862 7534 62914 7586
rect 62914 7534 62916 7586
rect 62860 7532 62916 7534
rect 62748 7084 62804 7140
rect 63084 6636 63140 6692
rect 62972 6524 63028 6580
rect 62636 5292 62692 5348
rect 62748 6300 62804 6356
rect 62412 4060 62468 4116
rect 62188 3276 62244 3332
rect 62300 3612 62356 3668
rect 62524 3388 62580 3444
rect 62860 5964 62916 6020
rect 62860 4172 62916 4228
rect 62748 3724 62804 3780
rect 62860 3948 62916 4004
rect 62636 3164 62692 3220
rect 63084 5906 63140 5908
rect 63084 5854 63086 5906
rect 63086 5854 63138 5906
rect 63138 5854 63140 5906
rect 63084 5852 63140 5854
rect 63868 8428 63924 8484
rect 63644 8316 63700 8372
rect 63532 8258 63588 8260
rect 63532 8206 63534 8258
rect 63534 8206 63586 8258
rect 63586 8206 63588 8258
rect 63532 8204 63588 8206
rect 63868 8258 63924 8260
rect 63868 8206 63870 8258
rect 63870 8206 63922 8258
rect 63922 8206 63924 8258
rect 63868 8204 63924 8206
rect 64428 9436 64484 9492
rect 64092 8092 64148 8148
rect 64204 9324 64260 9380
rect 63980 7868 64036 7924
rect 63868 7756 63924 7812
rect 64204 7532 64260 7588
rect 63532 7362 63588 7364
rect 63532 7310 63534 7362
rect 63534 7310 63586 7362
rect 63586 7310 63588 7362
rect 63532 7308 63588 7310
rect 63420 7250 63476 7252
rect 63420 7198 63422 7250
rect 63422 7198 63474 7250
rect 63474 7198 63476 7250
rect 63420 7196 63476 7198
rect 63420 6802 63476 6804
rect 63420 6750 63422 6802
rect 63422 6750 63474 6802
rect 63474 6750 63476 6802
rect 63420 6748 63476 6750
rect 63308 6412 63364 6468
rect 63868 6972 63924 7028
rect 63756 6860 63812 6916
rect 63084 1484 63140 1540
rect 63644 6748 63700 6804
rect 64204 6860 64260 6916
rect 63644 6300 63700 6356
rect 63756 6466 63812 6468
rect 63756 6414 63758 6466
rect 63758 6414 63810 6466
rect 63810 6414 63812 6466
rect 63756 6412 63812 6414
rect 63868 6300 63924 6356
rect 63532 4620 63588 4676
rect 63756 5906 63812 5908
rect 63756 5854 63758 5906
rect 63758 5854 63810 5906
rect 63810 5854 63812 5906
rect 63756 5852 63812 5854
rect 64652 9266 64708 9268
rect 64652 9214 64654 9266
rect 64654 9214 64706 9266
rect 64706 9214 64708 9266
rect 64652 9212 64708 9214
rect 64540 7474 64596 7476
rect 64540 7422 64542 7474
rect 64542 7422 64594 7474
rect 64594 7422 64596 7474
rect 64540 7420 64596 7422
rect 64652 8428 64708 8484
rect 64428 7308 64484 7364
rect 64428 6748 64484 6804
rect 64540 6578 64596 6580
rect 64540 6526 64542 6578
rect 64542 6526 64594 6578
rect 64594 6526 64596 6578
rect 64540 6524 64596 6526
rect 64316 6412 64372 6468
rect 63980 5292 64036 5348
rect 64204 5404 64260 5460
rect 64092 5180 64148 5236
rect 63644 4508 63700 4564
rect 63756 4732 63812 4788
rect 63420 4396 63476 4452
rect 63980 4620 64036 4676
rect 63868 4226 63924 4228
rect 63868 4174 63870 4226
rect 63870 4174 63922 4226
rect 63922 4174 63924 4226
rect 63868 4172 63924 4174
rect 64204 2716 64260 2772
rect 64652 6188 64708 6244
rect 64540 4620 64596 4676
rect 64652 5964 64708 6020
rect 64428 4508 64484 4564
rect 64540 4450 64596 4452
rect 64540 4398 64542 4450
rect 64542 4398 64594 4450
rect 64594 4398 64596 4450
rect 64540 4396 64596 4398
rect 64876 8428 64932 8484
rect 64988 8988 65044 9044
rect 64988 8258 65044 8260
rect 64988 8206 64990 8258
rect 64990 8206 65042 8258
rect 65042 8206 65044 8258
rect 64988 8204 65044 8206
rect 64988 7420 65044 7476
rect 64876 7084 64932 7140
rect 64876 6636 64932 6692
rect 64764 5180 64820 5236
rect 64652 4060 64708 4116
rect 64540 3724 64596 3780
rect 64876 3500 64932 3556
rect 65212 9884 65268 9940
rect 65324 9436 65380 9492
rect 65212 8764 65268 8820
rect 65324 8428 65380 8484
rect 65548 10444 65604 10500
rect 78492 17274 78548 17276
rect 78492 17222 78494 17274
rect 78494 17222 78546 17274
rect 78546 17222 78548 17274
rect 78492 17220 78548 17222
rect 78596 17274 78652 17276
rect 78596 17222 78598 17274
rect 78598 17222 78650 17274
rect 78650 17222 78652 17274
rect 78596 17220 78652 17222
rect 78700 17274 78756 17276
rect 78700 17222 78702 17274
rect 78702 17222 78754 17274
rect 78754 17222 78756 17274
rect 78700 17220 78756 17222
rect 68832 16490 68888 16492
rect 68832 16438 68834 16490
rect 68834 16438 68886 16490
rect 68886 16438 68888 16490
rect 68832 16436 68888 16438
rect 68936 16490 68992 16492
rect 68936 16438 68938 16490
rect 68938 16438 68990 16490
rect 68990 16438 68992 16490
rect 68936 16436 68992 16438
rect 69040 16490 69096 16492
rect 69040 16438 69042 16490
rect 69042 16438 69094 16490
rect 69094 16438 69096 16490
rect 69040 16436 69096 16438
rect 78492 15706 78548 15708
rect 78492 15654 78494 15706
rect 78494 15654 78546 15706
rect 78546 15654 78548 15706
rect 78492 15652 78548 15654
rect 78596 15706 78652 15708
rect 78596 15654 78598 15706
rect 78598 15654 78650 15706
rect 78650 15654 78652 15706
rect 78596 15652 78652 15654
rect 78700 15706 78756 15708
rect 78700 15654 78702 15706
rect 78702 15654 78754 15706
rect 78754 15654 78756 15706
rect 78700 15652 78756 15654
rect 69804 15148 69860 15204
rect 68832 14922 68888 14924
rect 68832 14870 68834 14922
rect 68834 14870 68886 14922
rect 68886 14870 68888 14922
rect 68832 14868 68888 14870
rect 68936 14922 68992 14924
rect 68936 14870 68938 14922
rect 68938 14870 68990 14922
rect 68990 14870 68992 14922
rect 68936 14868 68992 14870
rect 69040 14922 69096 14924
rect 69040 14870 69042 14922
rect 69042 14870 69094 14922
rect 69094 14870 69096 14922
rect 69040 14868 69096 14870
rect 68832 13354 68888 13356
rect 68832 13302 68834 13354
rect 68834 13302 68886 13354
rect 68886 13302 68888 13354
rect 68832 13300 68888 13302
rect 68936 13354 68992 13356
rect 68936 13302 68938 13354
rect 68938 13302 68990 13354
rect 68990 13302 68992 13354
rect 68936 13300 68992 13302
rect 69040 13354 69096 13356
rect 69040 13302 69042 13354
rect 69042 13302 69094 13354
rect 69094 13302 69096 13354
rect 69040 13300 69096 13302
rect 67116 11452 67172 11508
rect 67452 11900 67508 11956
rect 66556 9996 66612 10052
rect 66668 10220 66724 10276
rect 65660 9212 65716 9268
rect 65548 8988 65604 9044
rect 65660 8764 65716 8820
rect 65324 8034 65380 8036
rect 65324 7982 65326 8034
rect 65326 7982 65378 8034
rect 65378 7982 65380 8034
rect 65324 7980 65380 7982
rect 65548 8258 65604 8260
rect 65548 8206 65550 8258
rect 65550 8206 65602 8258
rect 65602 8206 65604 8258
rect 65548 8204 65604 8206
rect 65100 6300 65156 6356
rect 65100 5180 65156 5236
rect 65212 3724 65268 3780
rect 65548 7756 65604 7812
rect 65436 6748 65492 6804
rect 65660 6412 65716 6468
rect 66108 9212 66164 9268
rect 66780 9714 66836 9716
rect 66780 9662 66782 9714
rect 66782 9662 66834 9714
rect 66834 9662 66836 9714
rect 66780 9660 66836 9662
rect 65996 8988 66052 9044
rect 65996 8316 66052 8372
rect 65884 8204 65940 8260
rect 65884 7756 65940 7812
rect 65884 7308 65940 7364
rect 65996 7532 66052 7588
rect 66332 8316 66388 8372
rect 66668 8540 66724 8596
rect 66556 8204 66612 8260
rect 66220 7196 66276 7252
rect 66332 7084 66388 7140
rect 65548 4508 65604 4564
rect 65548 3836 65604 3892
rect 65436 3276 65492 3332
rect 65772 4396 65828 4452
rect 65884 4956 65940 5012
rect 65772 4172 65828 4228
rect 65660 3276 65716 3332
rect 65660 2492 65716 2548
rect 66108 6188 66164 6244
rect 67228 9660 67284 9716
rect 66668 7698 66724 7700
rect 66668 7646 66670 7698
rect 66670 7646 66722 7698
rect 66722 7646 66724 7698
rect 66668 7644 66724 7646
rect 66556 7532 66612 7588
rect 66668 7308 66724 7364
rect 66556 6972 66612 7028
rect 66892 8316 66948 8372
rect 66892 7756 66948 7812
rect 66780 6412 66836 6468
rect 66892 7084 66948 7140
rect 66668 4732 66724 4788
rect 66780 5068 66836 5124
rect 66444 4396 66500 4452
rect 68832 11786 68888 11788
rect 68832 11734 68834 11786
rect 68834 11734 68886 11786
rect 68886 11734 68888 11786
rect 68832 11732 68888 11734
rect 68936 11786 68992 11788
rect 68936 11734 68938 11786
rect 68938 11734 68990 11786
rect 68990 11734 68992 11786
rect 68936 11732 68992 11734
rect 69040 11786 69096 11788
rect 69040 11734 69042 11786
rect 69042 11734 69094 11786
rect 69094 11734 69096 11786
rect 69040 11732 69096 11734
rect 68908 11452 68964 11508
rect 69356 10668 69412 10724
rect 67228 8204 67284 8260
rect 67116 7308 67172 7364
rect 67116 6524 67172 6580
rect 67340 7586 67396 7588
rect 67340 7534 67342 7586
rect 67342 7534 67394 7586
rect 67394 7534 67396 7586
rect 67340 7532 67396 7534
rect 67340 7196 67396 7252
rect 67452 6636 67508 6692
rect 67452 6300 67508 6356
rect 67228 5404 67284 5460
rect 66892 4172 66948 4228
rect 66892 3500 66948 3556
rect 67228 4508 67284 4564
rect 67340 4620 67396 4676
rect 67228 4060 67284 4116
rect 67452 4508 67508 4564
rect 67900 9154 67956 9156
rect 67900 9102 67902 9154
rect 67902 9102 67954 9154
rect 67954 9102 67956 9154
rect 67900 9100 67956 9102
rect 67788 7980 67844 8036
rect 67900 8540 67956 8596
rect 68348 10444 68404 10500
rect 69132 10498 69188 10500
rect 69132 10446 69134 10498
rect 69134 10446 69186 10498
rect 69186 10446 69188 10498
rect 69132 10444 69188 10446
rect 68348 8540 68404 8596
rect 68348 8370 68404 8372
rect 68348 8318 68350 8370
rect 68350 8318 68402 8370
rect 68402 8318 68404 8370
rect 68348 8316 68404 8318
rect 68236 8204 68292 8260
rect 68124 8092 68180 8148
rect 68348 7980 68404 8036
rect 67900 7532 67956 7588
rect 67900 6972 67956 7028
rect 67788 6636 67844 6692
rect 67788 6018 67844 6020
rect 67788 5966 67790 6018
rect 67790 5966 67842 6018
rect 67842 5966 67844 6018
rect 67788 5964 67844 5966
rect 68012 5964 68068 6020
rect 67788 4956 67844 5012
rect 67900 4844 67956 4900
rect 67788 4732 67844 4788
rect 67564 4396 67620 4452
rect 67676 4172 67732 4228
rect 67452 3388 67508 3444
rect 68236 7532 68292 7588
rect 68832 10218 68888 10220
rect 68832 10166 68834 10218
rect 68834 10166 68886 10218
rect 68886 10166 68888 10218
rect 68832 10164 68888 10166
rect 68936 10218 68992 10220
rect 68936 10166 68938 10218
rect 68938 10166 68990 10218
rect 68990 10166 68992 10218
rect 68936 10164 68992 10166
rect 69040 10218 69096 10220
rect 69040 10166 69042 10218
rect 69042 10166 69094 10218
rect 69094 10166 69096 10218
rect 69040 10164 69096 10166
rect 69244 9996 69300 10052
rect 68460 7644 68516 7700
rect 68572 6972 68628 7028
rect 68572 6578 68628 6580
rect 68572 6526 68574 6578
rect 68574 6526 68626 6578
rect 68626 6526 68628 6578
rect 68572 6524 68628 6526
rect 68124 4956 68180 5012
rect 68124 4620 68180 4676
rect 68236 6412 68292 6468
rect 68124 4284 68180 4340
rect 68572 6188 68628 6244
rect 68348 6018 68404 6020
rect 68348 5966 68350 6018
rect 68350 5966 68402 6018
rect 68402 5966 68404 6018
rect 68348 5964 68404 5966
rect 68460 5010 68516 5012
rect 68460 4958 68462 5010
rect 68462 4958 68514 5010
rect 68514 4958 68516 5010
rect 68460 4956 68516 4958
rect 68348 4732 68404 4788
rect 68796 9100 68852 9156
rect 68832 8650 68888 8652
rect 68832 8598 68834 8650
rect 68834 8598 68886 8650
rect 68886 8598 68888 8650
rect 68832 8596 68888 8598
rect 68936 8650 68992 8652
rect 68936 8598 68938 8650
rect 68938 8598 68990 8650
rect 68990 8598 68992 8650
rect 68936 8596 68992 8598
rect 69040 8650 69096 8652
rect 69040 8598 69042 8650
rect 69042 8598 69094 8650
rect 69094 8598 69096 8650
rect 69040 8596 69096 8598
rect 68908 8092 68964 8148
rect 69020 7362 69076 7364
rect 69020 7310 69022 7362
rect 69022 7310 69074 7362
rect 69074 7310 69076 7362
rect 69020 7308 69076 7310
rect 68908 7196 68964 7252
rect 69356 8146 69412 8148
rect 69356 8094 69358 8146
rect 69358 8094 69410 8146
rect 69410 8094 69412 8146
rect 69356 8092 69412 8094
rect 68832 7082 68888 7084
rect 68832 7030 68834 7082
rect 68834 7030 68886 7082
rect 68886 7030 68888 7082
rect 68832 7028 68888 7030
rect 68936 7082 68992 7084
rect 68936 7030 68938 7082
rect 68938 7030 68990 7082
rect 68990 7030 68992 7082
rect 68936 7028 68992 7030
rect 69040 7082 69096 7084
rect 69040 7030 69042 7082
rect 69042 7030 69094 7082
rect 69094 7030 69096 7082
rect 69040 7028 69096 7030
rect 68832 5514 68888 5516
rect 68832 5462 68834 5514
rect 68834 5462 68886 5514
rect 68886 5462 68888 5514
rect 68832 5460 68888 5462
rect 68936 5514 68992 5516
rect 68936 5462 68938 5514
rect 68938 5462 68990 5514
rect 68990 5462 68992 5514
rect 68936 5460 68992 5462
rect 69040 5514 69096 5516
rect 69040 5462 69042 5514
rect 69042 5462 69094 5514
rect 69094 5462 69096 5514
rect 69040 5460 69096 5462
rect 69020 4956 69076 5012
rect 69244 4844 69300 4900
rect 68460 4060 68516 4116
rect 68796 4060 68852 4116
rect 68832 3946 68888 3948
rect 68832 3894 68834 3946
rect 68834 3894 68886 3946
rect 68886 3894 68888 3946
rect 68832 3892 68888 3894
rect 68936 3946 68992 3948
rect 68936 3894 68938 3946
rect 68938 3894 68990 3946
rect 68990 3894 68992 3946
rect 68936 3892 68992 3894
rect 69040 3946 69096 3948
rect 69040 3894 69042 3946
rect 69042 3894 69094 3946
rect 69094 3894 69096 3946
rect 69040 3892 69096 3894
rect 69020 3500 69076 3556
rect 78492 14138 78548 14140
rect 78492 14086 78494 14138
rect 78494 14086 78546 14138
rect 78546 14086 78548 14138
rect 78492 14084 78548 14086
rect 78596 14138 78652 14140
rect 78596 14086 78598 14138
rect 78598 14086 78650 14138
rect 78650 14086 78652 14138
rect 78596 14084 78652 14086
rect 78700 14138 78756 14140
rect 78700 14086 78702 14138
rect 78702 14086 78754 14138
rect 78754 14086 78756 14138
rect 78700 14084 78756 14086
rect 78492 12570 78548 12572
rect 78492 12518 78494 12570
rect 78494 12518 78546 12570
rect 78546 12518 78548 12570
rect 78492 12516 78548 12518
rect 78596 12570 78652 12572
rect 78596 12518 78598 12570
rect 78598 12518 78650 12570
rect 78650 12518 78652 12570
rect 78596 12516 78652 12518
rect 78700 12570 78756 12572
rect 78700 12518 78702 12570
rect 78702 12518 78754 12570
rect 78754 12518 78756 12570
rect 78700 12516 78756 12518
rect 69804 9772 69860 9828
rect 70252 10722 70308 10724
rect 70252 10670 70254 10722
rect 70254 10670 70306 10722
rect 70306 10670 70308 10722
rect 70252 10668 70308 10670
rect 70140 10556 70196 10612
rect 69580 9042 69636 9044
rect 69580 8990 69582 9042
rect 69582 8990 69634 9042
rect 69634 8990 69636 9042
rect 69580 8988 69636 8990
rect 69580 8540 69636 8596
rect 70140 8540 70196 8596
rect 70252 8652 70308 8708
rect 70140 8204 70196 8260
rect 70028 7420 70084 7476
rect 69916 7084 69972 7140
rect 69804 6972 69860 7028
rect 70028 6860 70084 6916
rect 69580 6076 69636 6132
rect 69692 5740 69748 5796
rect 69468 4956 69524 5012
rect 69580 5180 69636 5236
rect 69468 4396 69524 4452
rect 69804 4844 69860 4900
rect 69804 4396 69860 4452
rect 69132 3052 69188 3108
rect 70140 5964 70196 6020
rect 70700 10332 70756 10388
rect 70476 9772 70532 9828
rect 70588 8988 70644 9044
rect 70476 6076 70532 6132
rect 71260 9826 71316 9828
rect 71260 9774 71262 9826
rect 71262 9774 71314 9826
rect 71314 9774 71316 9826
rect 71260 9772 71316 9774
rect 71372 9436 71428 9492
rect 71484 9212 71540 9268
rect 71260 9154 71316 9156
rect 71260 9102 71262 9154
rect 71262 9102 71314 9154
rect 71314 9102 71316 9154
rect 71260 9100 71316 9102
rect 71148 9042 71204 9044
rect 71148 8990 71150 9042
rect 71150 8990 71202 9042
rect 71202 8990 71204 9042
rect 71148 8988 71204 8990
rect 71036 8652 71092 8708
rect 71036 8428 71092 8484
rect 70700 7644 70756 7700
rect 70476 5628 70532 5684
rect 70588 5234 70644 5236
rect 70588 5182 70590 5234
rect 70590 5182 70642 5234
rect 70642 5182 70644 5234
rect 70588 5180 70644 5182
rect 70364 5068 70420 5124
rect 71148 7474 71204 7476
rect 71148 7422 71150 7474
rect 71150 7422 71202 7474
rect 71202 7422 71204 7474
rect 71148 7420 71204 7422
rect 70812 5852 70868 5908
rect 71148 7196 71204 7252
rect 71036 6076 71092 6132
rect 70476 4956 70532 5012
rect 70364 4844 70420 4900
rect 70812 5628 70868 5684
rect 70924 5516 70980 5572
rect 70924 4396 70980 4452
rect 71036 3724 71092 3780
rect 71260 7084 71316 7140
rect 71484 6748 71540 6804
rect 71484 4396 71540 4452
rect 71708 9324 71764 9380
rect 71708 8540 71764 8596
rect 71932 10556 71988 10612
rect 71932 8540 71988 8596
rect 72044 8316 72100 8372
rect 71596 4284 71652 4340
rect 71708 5404 71764 5460
rect 71932 7308 71988 7364
rect 72380 9602 72436 9604
rect 72380 9550 72382 9602
rect 72382 9550 72434 9602
rect 72434 9550 72436 9602
rect 72380 9548 72436 9550
rect 72268 9212 72324 9268
rect 72268 8930 72324 8932
rect 72268 8878 72270 8930
rect 72270 8878 72322 8930
rect 72322 8878 72324 8930
rect 72268 8876 72324 8878
rect 72380 7196 72436 7252
rect 72604 9436 72660 9492
rect 72604 7644 72660 7700
rect 72604 7420 72660 7476
rect 72044 4956 72100 5012
rect 72380 6636 72436 6692
rect 72380 6018 72436 6020
rect 72380 5966 72382 6018
rect 72382 5966 72434 6018
rect 72434 5966 72436 6018
rect 72380 5964 72436 5966
rect 72380 5180 72436 5236
rect 71820 2492 71876 2548
rect 71932 3724 71988 3780
rect 72044 3276 72100 3332
rect 72156 3388 72212 3444
rect 72492 4620 72548 4676
rect 72828 10610 72884 10612
rect 72828 10558 72830 10610
rect 72830 10558 72882 10610
rect 72882 10558 72884 10610
rect 72828 10556 72884 10558
rect 72940 8876 72996 8932
rect 72828 7084 72884 7140
rect 72828 6802 72884 6804
rect 72828 6750 72830 6802
rect 72830 6750 72882 6802
rect 72882 6750 72884 6802
rect 72828 6748 72884 6750
rect 72716 6636 72772 6692
rect 73388 8764 73444 8820
rect 73276 8540 73332 8596
rect 73164 8370 73220 8372
rect 73164 8318 73166 8370
rect 73166 8318 73218 8370
rect 73218 8318 73220 8370
rect 73164 8316 73220 8318
rect 73724 8428 73780 8484
rect 73276 7308 73332 7364
rect 73388 7980 73444 8036
rect 73164 6636 73220 6692
rect 73276 6076 73332 6132
rect 72828 5852 72884 5908
rect 72828 5628 72884 5684
rect 72828 4956 72884 5012
rect 73276 5068 73332 5124
rect 73164 4284 73220 4340
rect 73164 2828 73220 2884
rect 73724 7362 73780 7364
rect 73724 7310 73726 7362
rect 73726 7310 73778 7362
rect 73778 7310 73780 7362
rect 73724 7308 73780 7310
rect 73724 7084 73780 7140
rect 73612 6636 73668 6692
rect 73612 5852 73668 5908
rect 74172 6524 74228 6580
rect 74508 9548 74564 9604
rect 74508 8764 74564 8820
rect 74396 4956 74452 5012
rect 74956 9602 75012 9604
rect 74956 9550 74958 9602
rect 74958 9550 75010 9602
rect 75010 9550 75012 9602
rect 74956 9548 75012 9550
rect 74732 5516 74788 5572
rect 74284 4620 74340 4676
rect 73836 4508 73892 4564
rect 73612 4060 73668 4116
rect 74284 4060 74340 4116
rect 75628 9660 75684 9716
rect 75516 6860 75572 6916
rect 75628 7420 75684 7476
rect 75852 9772 75908 9828
rect 75740 6524 75796 6580
rect 75180 5628 75236 5684
rect 75628 5964 75684 6020
rect 75180 4450 75236 4452
rect 75180 4398 75182 4450
rect 75182 4398 75234 4450
rect 75234 4398 75236 4450
rect 75180 4396 75236 4398
rect 74956 3500 75012 3556
rect 76636 9212 76692 9268
rect 76188 8652 76244 8708
rect 76188 8092 76244 8148
rect 76300 6578 76356 6580
rect 76300 6526 76302 6578
rect 76302 6526 76354 6578
rect 76354 6526 76356 6578
rect 76300 6524 76356 6526
rect 76860 10780 76916 10836
rect 78492 11002 78548 11004
rect 78492 10950 78494 11002
rect 78494 10950 78546 11002
rect 78546 10950 78548 11002
rect 78492 10948 78548 10950
rect 78596 11002 78652 11004
rect 78596 10950 78598 11002
rect 78598 10950 78650 11002
rect 78650 10950 78652 11002
rect 78596 10948 78652 10950
rect 78700 11002 78756 11004
rect 78700 10950 78702 11002
rect 78702 10950 78754 11002
rect 78754 10950 78756 11002
rect 78700 10948 78756 10950
rect 77308 10892 77364 10948
rect 77532 9884 77588 9940
rect 76860 9154 76916 9156
rect 76860 9102 76862 9154
rect 76862 9102 76914 9154
rect 76914 9102 76916 9154
rect 76860 9100 76916 9102
rect 76748 5852 76804 5908
rect 76860 7532 76916 7588
rect 76300 5180 76356 5236
rect 75964 5068 76020 5124
rect 76076 4508 76132 4564
rect 77084 9212 77140 9268
rect 77420 8988 77476 9044
rect 77084 7868 77140 7924
rect 76972 6972 77028 7028
rect 77084 6748 77140 6804
rect 77196 5404 77252 5460
rect 77532 7084 77588 7140
rect 77756 7196 77812 7252
rect 78092 8316 78148 8372
rect 77980 8034 78036 8036
rect 77980 7982 77982 8034
rect 77982 7982 78034 8034
rect 78034 7982 78036 8034
rect 77980 7980 78036 7982
rect 77980 7474 78036 7476
rect 77980 7422 77982 7474
rect 77982 7422 78034 7474
rect 78034 7422 78036 7474
rect 77980 7420 78036 7422
rect 78092 7308 78148 7364
rect 77980 6466 78036 6468
rect 77980 6414 77982 6466
rect 77982 6414 78034 6466
rect 78034 6414 78036 6466
rect 77980 6412 78036 6414
rect 77868 6018 77924 6020
rect 77868 5966 77870 6018
rect 77870 5966 77922 6018
rect 77922 5966 77924 6018
rect 77868 5964 77924 5966
rect 77532 5292 77588 5348
rect 77644 5852 77700 5908
rect 75628 3164 75684 3220
rect 78092 3724 78148 3780
rect 78428 9660 78484 9716
rect 78492 9434 78548 9436
rect 78492 9382 78494 9434
rect 78494 9382 78546 9434
rect 78546 9382 78548 9434
rect 78492 9380 78548 9382
rect 78596 9434 78652 9436
rect 78596 9382 78598 9434
rect 78598 9382 78650 9434
rect 78650 9382 78652 9434
rect 78596 9380 78652 9382
rect 78700 9434 78756 9436
rect 78700 9382 78702 9434
rect 78702 9382 78754 9434
rect 78754 9382 78756 9434
rect 78700 9380 78756 9382
rect 78492 7866 78548 7868
rect 78492 7814 78494 7866
rect 78494 7814 78546 7866
rect 78546 7814 78548 7866
rect 78492 7812 78548 7814
rect 78596 7866 78652 7868
rect 78596 7814 78598 7866
rect 78598 7814 78650 7866
rect 78650 7814 78652 7866
rect 78596 7812 78652 7814
rect 78700 7866 78756 7868
rect 78700 7814 78702 7866
rect 78702 7814 78754 7866
rect 78754 7814 78756 7866
rect 78700 7812 78756 7814
rect 78492 6298 78548 6300
rect 78492 6246 78494 6298
rect 78494 6246 78546 6298
rect 78546 6246 78548 6298
rect 78492 6244 78548 6246
rect 78596 6298 78652 6300
rect 78596 6246 78598 6298
rect 78598 6246 78650 6298
rect 78650 6246 78652 6298
rect 78596 6244 78652 6246
rect 78700 6298 78756 6300
rect 78700 6246 78702 6298
rect 78702 6246 78754 6298
rect 78754 6246 78756 6298
rect 78700 6244 78756 6246
rect 78492 4730 78548 4732
rect 78492 4678 78494 4730
rect 78494 4678 78546 4730
rect 78546 4678 78548 4730
rect 78492 4676 78548 4678
rect 78596 4730 78652 4732
rect 78596 4678 78598 4730
rect 78598 4678 78650 4730
rect 78650 4678 78652 4730
rect 78596 4676 78652 4678
rect 78700 4730 78756 4732
rect 78700 4678 78702 4730
rect 78702 4678 78754 4730
rect 78754 4678 78756 4730
rect 78700 4676 78756 4678
rect 78092 3388 78148 3444
rect 78492 3162 78548 3164
rect 78492 3110 78494 3162
rect 78494 3110 78546 3162
rect 78546 3110 78548 3162
rect 78492 3108 78548 3110
rect 78596 3162 78652 3164
rect 78596 3110 78598 3162
rect 78598 3110 78650 3162
rect 78650 3110 78652 3162
rect 78596 3108 78652 3110
rect 78700 3162 78756 3164
rect 78700 3110 78702 3162
rect 78702 3110 78754 3162
rect 78754 3110 78756 3162
rect 78700 3108 78756 3110
rect 77980 2940 78036 2996
<< metal3 >>
rect 10862 36820 10872 36876
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 11136 36820 11146 36876
rect 30182 36820 30192 36876
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30456 36820 30466 36876
rect 49502 36820 49512 36876
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49776 36820 49786 36876
rect 68822 36820 68832 36876
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 69096 36820 69106 36876
rect 20522 36036 20532 36092
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20796 36036 20806 36092
rect 39842 36036 39852 36092
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 40116 36036 40126 36092
rect 59162 36036 59172 36092
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59436 36036 59446 36092
rect 78482 36036 78492 36092
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78756 36036 78766 36092
rect 10862 35252 10872 35308
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 11136 35252 11146 35308
rect 30182 35252 30192 35308
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30456 35252 30466 35308
rect 49502 35252 49512 35308
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49776 35252 49786 35308
rect 68822 35252 68832 35308
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 69096 35252 69106 35308
rect 20522 34468 20532 34524
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20796 34468 20806 34524
rect 39842 34468 39852 34524
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 40116 34468 40126 34524
rect 59162 34468 59172 34524
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59436 34468 59446 34524
rect 78482 34468 78492 34524
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78756 34468 78766 34524
rect 10862 33684 10872 33740
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 11136 33684 11146 33740
rect 30182 33684 30192 33740
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30456 33684 30466 33740
rect 49502 33684 49512 33740
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49776 33684 49786 33740
rect 68822 33684 68832 33740
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 69096 33684 69106 33740
rect 20522 32900 20532 32956
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20796 32900 20806 32956
rect 39842 32900 39852 32956
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 40116 32900 40126 32956
rect 59162 32900 59172 32956
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59436 32900 59446 32956
rect 78482 32900 78492 32956
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78756 32900 78766 32956
rect 10862 32116 10872 32172
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 11136 32116 11146 32172
rect 30182 32116 30192 32172
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30456 32116 30466 32172
rect 49502 32116 49512 32172
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49776 32116 49786 32172
rect 68822 32116 68832 32172
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 69096 32116 69106 32172
rect 20522 31332 20532 31388
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20796 31332 20806 31388
rect 39842 31332 39852 31388
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 40116 31332 40126 31388
rect 59162 31332 59172 31388
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59436 31332 59446 31388
rect 78482 31332 78492 31388
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78756 31332 78766 31388
rect 10862 30548 10872 30604
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 11136 30548 11146 30604
rect 30182 30548 30192 30604
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30456 30548 30466 30604
rect 49502 30548 49512 30604
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49776 30548 49786 30604
rect 68822 30548 68832 30604
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 69096 30548 69106 30604
rect 20522 29764 20532 29820
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20796 29764 20806 29820
rect 39842 29764 39852 29820
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 40116 29764 40126 29820
rect 59162 29764 59172 29820
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59436 29764 59446 29820
rect 78482 29764 78492 29820
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78756 29764 78766 29820
rect 10862 28980 10872 29036
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 11136 28980 11146 29036
rect 30182 28980 30192 29036
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30456 28980 30466 29036
rect 49502 28980 49512 29036
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49776 28980 49786 29036
rect 68822 28980 68832 29036
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 69096 28980 69106 29036
rect 20522 28196 20532 28252
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20796 28196 20806 28252
rect 39842 28196 39852 28252
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 40116 28196 40126 28252
rect 59162 28196 59172 28252
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59436 28196 59446 28252
rect 78482 28196 78492 28252
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78756 28196 78766 28252
rect 10862 27412 10872 27468
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 11136 27412 11146 27468
rect 30182 27412 30192 27468
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30456 27412 30466 27468
rect 49502 27412 49512 27468
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49776 27412 49786 27468
rect 68822 27412 68832 27468
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69096 27412 69106 27468
rect 20522 26628 20532 26684
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20796 26628 20806 26684
rect 39842 26628 39852 26684
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 40116 26628 40126 26684
rect 59162 26628 59172 26684
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59436 26628 59446 26684
rect 78482 26628 78492 26684
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78756 26628 78766 26684
rect 10862 25844 10872 25900
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 11136 25844 11146 25900
rect 30182 25844 30192 25900
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30456 25844 30466 25900
rect 49502 25844 49512 25900
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49776 25844 49786 25900
rect 68822 25844 68832 25900
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 69096 25844 69106 25900
rect 20522 25060 20532 25116
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20796 25060 20806 25116
rect 39842 25060 39852 25116
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 40116 25060 40126 25116
rect 59162 25060 59172 25116
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59436 25060 59446 25116
rect 78482 25060 78492 25116
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78756 25060 78766 25116
rect 10862 24276 10872 24332
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11136 24276 11146 24332
rect 30182 24276 30192 24332
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30456 24276 30466 24332
rect 49502 24276 49512 24332
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49776 24276 49786 24332
rect 68822 24276 68832 24332
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 69096 24276 69106 24332
rect 20522 23492 20532 23548
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20796 23492 20806 23548
rect 39842 23492 39852 23548
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 40116 23492 40126 23548
rect 59162 23492 59172 23548
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59436 23492 59446 23548
rect 78482 23492 78492 23548
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78756 23492 78766 23548
rect 10862 22708 10872 22764
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 11136 22708 11146 22764
rect 30182 22708 30192 22764
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30456 22708 30466 22764
rect 49502 22708 49512 22764
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49776 22708 49786 22764
rect 68822 22708 68832 22764
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 69096 22708 69106 22764
rect 20522 21924 20532 21980
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20796 21924 20806 21980
rect 39842 21924 39852 21980
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 40116 21924 40126 21980
rect 59162 21924 59172 21980
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59436 21924 59446 21980
rect 78482 21924 78492 21980
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78756 21924 78766 21980
rect 10862 21140 10872 21196
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 11136 21140 11146 21196
rect 30182 21140 30192 21196
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30456 21140 30466 21196
rect 49502 21140 49512 21196
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49776 21140 49786 21196
rect 68822 21140 68832 21196
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 69096 21140 69106 21196
rect 20522 20356 20532 20412
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20796 20356 20806 20412
rect 39842 20356 39852 20412
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 40116 20356 40126 20412
rect 59162 20356 59172 20412
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59436 20356 59446 20412
rect 78482 20356 78492 20412
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78756 20356 78766 20412
rect 10862 19572 10872 19628
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 11136 19572 11146 19628
rect 30182 19572 30192 19628
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30456 19572 30466 19628
rect 49502 19572 49512 19628
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49776 19572 49786 19628
rect 68822 19572 68832 19628
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 69096 19572 69106 19628
rect 20522 18788 20532 18844
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20796 18788 20806 18844
rect 39842 18788 39852 18844
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 40116 18788 40126 18844
rect 59162 18788 59172 18844
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59436 18788 59446 18844
rect 78482 18788 78492 18844
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78756 18788 78766 18844
rect 16706 18508 16716 18564
rect 16772 18508 54572 18564
rect 54628 18508 54638 18564
rect 10862 18004 10872 18060
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 11136 18004 11146 18060
rect 30182 18004 30192 18060
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30456 18004 30466 18060
rect 49502 18004 49512 18060
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49776 18004 49786 18060
rect 68822 18004 68832 18060
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 69096 18004 69106 18060
rect 4834 17388 4844 17444
rect 4900 17388 67116 17444
rect 67172 17388 67182 17444
rect 20522 17220 20532 17276
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20796 17220 20806 17276
rect 39842 17220 39852 17276
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40116 17220 40126 17276
rect 59162 17220 59172 17276
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59436 17220 59446 17276
rect 78482 17220 78492 17276
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78756 17220 78766 17276
rect 22540 17164 37772 17220
rect 37828 17164 37838 17220
rect 22540 17108 22596 17164
rect 20178 17052 20188 17108
rect 20244 17052 22596 17108
rect 27570 17052 27580 17108
rect 27636 17052 48300 17108
rect 48356 17052 48366 17108
rect 28802 16940 28812 16996
rect 28868 16940 56028 16996
rect 56084 16940 56094 16996
rect 23762 16828 23772 16884
rect 23828 16828 42252 16884
rect 42308 16828 42318 16884
rect 10862 16436 10872 16492
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11136 16436 11146 16492
rect 30182 16436 30192 16492
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30456 16436 30466 16492
rect 49502 16436 49512 16492
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49776 16436 49786 16492
rect 68822 16436 68832 16492
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 69096 16436 69106 16492
rect 27346 15820 27356 15876
rect 27412 15820 31836 15876
rect 31892 15820 48524 15876
rect 48580 15820 48590 15876
rect 31938 15708 31948 15764
rect 32004 15708 35028 15764
rect 20522 15652 20532 15708
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20796 15652 20806 15708
rect 28242 15596 28252 15652
rect 28308 15596 32228 15652
rect 32498 15596 32508 15652
rect 32564 15596 34748 15652
rect 34804 15596 34814 15652
rect 31266 15484 31276 15540
rect 31332 15484 31948 15540
rect 32004 15484 32014 15540
rect 32172 15428 32228 15596
rect 34972 15540 35028 15708
rect 39842 15652 39852 15708
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40116 15652 40126 15708
rect 59162 15652 59172 15708
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59436 15652 59446 15708
rect 78482 15652 78492 15708
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78756 15652 78766 15708
rect 34972 15484 51436 15540
rect 51492 15484 51502 15540
rect 32172 15372 57372 15428
rect 57428 15372 57438 15428
rect 4946 15260 4956 15316
rect 5012 15260 54236 15316
rect 54292 15260 54302 15316
rect 6402 15148 6412 15204
rect 6468 15148 69804 15204
rect 69860 15148 69870 15204
rect 10862 14868 10872 14924
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 11136 14868 11146 14924
rect 30182 14868 30192 14924
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30456 14868 30466 14924
rect 49502 14868 49512 14924
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49776 14868 49786 14924
rect 68822 14868 68832 14924
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 69096 14868 69106 14924
rect 20522 14084 20532 14140
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20796 14084 20806 14140
rect 39842 14084 39852 14140
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 40116 14084 40126 14140
rect 59162 14084 59172 14140
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59436 14084 59446 14140
rect 78482 14084 78492 14140
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78756 14084 78766 14140
rect 30930 14028 30940 14084
rect 30996 14028 35756 14084
rect 35812 14028 35822 14084
rect 19282 13916 19292 13972
rect 19348 13916 46060 13972
rect 46116 13916 46126 13972
rect 33394 13804 33404 13860
rect 33460 13804 35308 13860
rect 35364 13804 35374 13860
rect 38098 13804 38108 13860
rect 38164 13804 39900 13860
rect 39956 13804 39966 13860
rect 10434 13692 10444 13748
rect 10500 13692 28924 13748
rect 28980 13692 28990 13748
rect 33282 13692 33292 13748
rect 33348 13692 34524 13748
rect 34580 13692 37100 13748
rect 37156 13692 37166 13748
rect 40562 13580 40572 13636
rect 40628 13580 55692 13636
rect 55748 13580 55758 13636
rect 14914 13468 14924 13524
rect 14980 13468 41468 13524
rect 41524 13468 41534 13524
rect 43362 13468 43372 13524
rect 43428 13468 56252 13524
rect 56308 13468 56318 13524
rect 32162 13356 32172 13412
rect 32228 13356 37548 13412
rect 37604 13356 37614 13412
rect 10862 13300 10872 13356
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 11136 13300 11146 13356
rect 30182 13300 30192 13356
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30456 13300 30466 13356
rect 49502 13300 49512 13356
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49776 13300 49786 13356
rect 68822 13300 68832 13356
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 69096 13300 69106 13356
rect 31602 13244 31612 13300
rect 31668 13244 41076 13300
rect 41020 13188 41076 13244
rect 17938 13132 17948 13188
rect 18004 13132 40236 13188
rect 40292 13132 40302 13188
rect 41020 13132 53228 13188
rect 53284 13132 53294 13188
rect 37762 13020 37772 13076
rect 37828 13020 38892 13076
rect 38948 13020 38958 13076
rect 44034 13020 44044 13076
rect 44100 13020 46172 13076
rect 46228 13020 46238 13076
rect 9538 12908 9548 12964
rect 9604 12908 10108 12964
rect 10164 12908 13244 12964
rect 13300 12908 13310 12964
rect 36306 12908 36316 12964
rect 36372 12908 36988 12964
rect 37044 12908 37054 12964
rect 40226 12796 40236 12852
rect 40292 12796 41356 12852
rect 41412 12796 41422 12852
rect 18274 12684 18284 12740
rect 18340 12684 20860 12740
rect 20916 12684 22540 12740
rect 22596 12684 24108 12740
rect 24164 12684 24174 12740
rect 24994 12684 25004 12740
rect 25060 12684 25900 12740
rect 25956 12684 25966 12740
rect 31602 12684 31612 12740
rect 31668 12684 33292 12740
rect 33348 12684 37660 12740
rect 37716 12684 37726 12740
rect 38612 12684 40516 12740
rect 41570 12684 41580 12740
rect 41636 12684 43932 12740
rect 43988 12684 43998 12740
rect 38612 12628 38668 12684
rect 40460 12628 40516 12684
rect 35410 12572 35420 12628
rect 35476 12572 38668 12628
rect 40450 12572 40460 12628
rect 40516 12572 42364 12628
rect 42420 12572 42812 12628
rect 42868 12572 48076 12628
rect 48132 12572 48142 12628
rect 20522 12516 20532 12572
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20796 12516 20806 12572
rect 39842 12516 39852 12572
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 40116 12516 40126 12572
rect 59162 12516 59172 12572
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59436 12516 59446 12572
rect 78482 12516 78492 12572
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78756 12516 78766 12572
rect 37202 12460 37212 12516
rect 37268 12460 38556 12516
rect 38612 12460 38622 12516
rect 40572 12460 46172 12516
rect 46228 12460 46238 12516
rect 40572 12404 40628 12460
rect 9762 12348 9772 12404
rect 9828 12348 21028 12404
rect 24210 12348 24220 12404
rect 24276 12348 25452 12404
rect 25508 12348 40628 12404
rect 40786 12348 40796 12404
rect 40852 12348 42028 12404
rect 42084 12348 44268 12404
rect 44324 12348 44334 12404
rect 20972 12292 21028 12348
rect 19618 12236 19628 12292
rect 19684 12236 20300 12292
rect 20356 12236 20366 12292
rect 20972 12236 30044 12292
rect 30100 12236 30110 12292
rect 30268 12236 31836 12292
rect 31892 12236 32340 12292
rect 43250 12236 43260 12292
rect 43316 12236 45612 12292
rect 45668 12236 45678 12292
rect 13682 12124 13692 12180
rect 13748 12124 15260 12180
rect 15316 12124 17500 12180
rect 17556 12124 17566 12180
rect 30268 12068 30324 12236
rect 32284 12180 32340 12236
rect 31154 12124 31164 12180
rect 31220 12124 31724 12180
rect 31780 12124 31790 12180
rect 32274 12124 32284 12180
rect 32340 12124 35532 12180
rect 35588 12124 35598 12180
rect 40338 12124 40348 12180
rect 40404 12124 40572 12180
rect 40628 12124 41580 12180
rect 41636 12124 41646 12180
rect 46386 12124 46396 12180
rect 46452 12124 58828 12180
rect 58884 12124 58894 12180
rect 26226 12012 26236 12068
rect 26292 12012 26796 12068
rect 26852 12012 30324 12068
rect 30482 12012 30492 12068
rect 30548 12012 31388 12068
rect 31444 12012 31454 12068
rect 32386 12012 32396 12068
rect 32452 12012 33852 12068
rect 33908 12012 33918 12068
rect 37314 12012 37324 12068
rect 37380 12012 38892 12068
rect 38948 12012 38958 12068
rect 41234 12012 41244 12068
rect 41300 12012 42476 12068
rect 42532 12012 50316 12068
rect 50372 12012 50382 12068
rect 25778 11900 25788 11956
rect 25844 11900 26684 11956
rect 26740 11900 31052 11956
rect 31108 11900 31724 11956
rect 31780 11900 31790 11956
rect 33506 11900 33516 11956
rect 33572 11900 39116 11956
rect 39172 11900 39182 11956
rect 39890 11900 39900 11956
rect 39956 11900 48860 11956
rect 48916 11900 48926 11956
rect 58034 11900 58044 11956
rect 58100 11900 67452 11956
rect 67508 11900 67518 11956
rect 11666 11788 11676 11844
rect 11732 11788 12908 11844
rect 12964 11788 12974 11844
rect 22642 11788 22652 11844
rect 22708 11788 25340 11844
rect 25396 11788 25406 11844
rect 34626 11788 34636 11844
rect 34692 11788 35980 11844
rect 36036 11788 36046 11844
rect 37650 11788 37660 11844
rect 37716 11788 40908 11844
rect 40964 11788 40974 11844
rect 43138 11788 43148 11844
rect 43204 11788 48748 11844
rect 48804 11788 48814 11844
rect 57698 11788 57708 11844
rect 57764 11788 66556 11844
rect 66612 11788 66622 11844
rect 10862 11732 10872 11788
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 11136 11732 11146 11788
rect 30182 11732 30192 11788
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30456 11732 30466 11788
rect 49502 11732 49512 11788
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49776 11732 49786 11788
rect 68822 11732 68832 11788
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 69096 11732 69106 11788
rect 37090 11676 37100 11732
rect 37156 11676 37884 11732
rect 37940 11676 37950 11732
rect 16930 11564 16940 11620
rect 16996 11564 44212 11620
rect 47506 11564 47516 11620
rect 47572 11564 59052 11620
rect 59108 11564 59118 11620
rect 21746 11452 21756 11508
rect 21812 11452 23436 11508
rect 23492 11452 23502 11508
rect 26114 11452 26124 11508
rect 26180 11452 28252 11508
rect 28308 11452 28318 11508
rect 19842 11340 19852 11396
rect 19908 11340 21420 11396
rect 21476 11340 21486 11396
rect 32834 11340 32844 11396
rect 32900 11340 35308 11396
rect 35364 11340 36316 11396
rect 36372 11340 36382 11396
rect 12114 11228 12124 11284
rect 12180 11228 13132 11284
rect 13188 11228 14700 11284
rect 14756 11228 14766 11284
rect 15138 11228 15148 11284
rect 15204 11228 16492 11284
rect 16548 11228 16558 11284
rect 18162 11228 18172 11284
rect 18228 11228 20412 11284
rect 20468 11228 20478 11284
rect 22194 11228 22204 11284
rect 22260 11228 22540 11284
rect 22596 11228 22606 11284
rect 22764 11228 23324 11284
rect 23380 11228 23390 11284
rect 29922 11228 29932 11284
rect 29988 11228 31164 11284
rect 31220 11228 31230 11284
rect 38210 11228 38220 11284
rect 38276 11228 41916 11284
rect 41972 11228 41982 11284
rect 22764 11172 22820 11228
rect 44156 11172 44212 11564
rect 47012 11452 50092 11508
rect 50148 11452 50158 11508
rect 67106 11452 67116 11508
rect 67172 11452 68908 11508
rect 68964 11452 68974 11508
rect 47012 11396 47068 11452
rect 45714 11340 45724 11396
rect 45780 11340 46172 11396
rect 46228 11340 47068 11396
rect 44370 11228 44380 11284
rect 44436 11228 45948 11284
rect 46004 11228 46014 11284
rect 48738 11228 48748 11284
rect 48804 11228 51548 11284
rect 51604 11228 51614 11284
rect 12338 11116 12348 11172
rect 12404 11116 13580 11172
rect 13636 11116 13646 11172
rect 18834 11116 18844 11172
rect 18900 11116 22764 11172
rect 22820 11116 22830 11172
rect 23090 11116 23100 11172
rect 23156 11116 24444 11172
rect 24500 11116 26236 11172
rect 26292 11116 26302 11172
rect 27234 11116 27244 11172
rect 27300 11116 28588 11172
rect 28644 11116 28654 11172
rect 29250 11116 29260 11172
rect 29316 11116 39676 11172
rect 39732 11116 42140 11172
rect 42196 11116 42812 11172
rect 42868 11116 43708 11172
rect 43764 11116 43774 11172
rect 44156 11116 44940 11172
rect 44996 11116 45612 11172
rect 45668 11116 46956 11172
rect 47012 11116 47022 11172
rect 47618 11116 47628 11172
rect 47684 11116 48636 11172
rect 48692 11116 48702 11172
rect 22306 11004 22316 11060
rect 22372 11004 26908 11060
rect 32946 11004 32956 11060
rect 33012 11004 33852 11060
rect 33908 11004 35420 11060
rect 35476 11004 35486 11060
rect 40236 11004 52332 11060
rect 52388 11004 52398 11060
rect 20522 10948 20532 11004
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20796 10948 20806 11004
rect 26852 10948 26908 11004
rect 39842 10948 39852 11004
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 40116 10948 40126 11004
rect 26852 10892 35364 10948
rect 35634 10892 35644 10948
rect 35700 10892 37548 10948
rect 37604 10892 37614 10948
rect 19292 10780 29148 10836
rect 29204 10780 33628 10836
rect 33684 10780 33694 10836
rect 19292 10724 19348 10780
rect 14466 10668 14476 10724
rect 14532 10668 15820 10724
rect 15876 10668 19348 10724
rect 24546 10668 24556 10724
rect 24612 10668 25228 10724
rect 25284 10668 25294 10724
rect 27794 10668 27804 10724
rect 27860 10668 30604 10724
rect 30660 10668 30670 10724
rect 29810 10556 29820 10612
rect 29876 10556 31164 10612
rect 31220 10556 31230 10612
rect 11732 10444 12236 10500
rect 12292 10444 14028 10500
rect 14084 10444 16380 10500
rect 16436 10444 16828 10500
rect 16884 10444 17500 10500
rect 17556 10444 18284 10500
rect 18340 10444 18350 10500
rect 26226 10444 26236 10500
rect 26292 10444 27244 10500
rect 27300 10444 27310 10500
rect 29250 10444 29260 10500
rect 29316 10444 30828 10500
rect 30884 10444 32844 10500
rect 32900 10444 32910 10500
rect 10862 10164 10872 10220
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 11136 10164 11146 10220
rect 11732 10164 11788 10444
rect 35308 10388 35364 10892
rect 40236 10836 40292 11004
rect 59162 10948 59172 11004
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59436 10948 59446 11004
rect 78482 10948 78492 11004
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78756 10948 78766 11004
rect 41010 10892 41020 10948
rect 41076 10892 41356 10948
rect 41412 10892 41422 10948
rect 46162 10892 46172 10948
rect 46228 10892 53788 10948
rect 53844 10892 53854 10948
rect 60834 10892 60844 10948
rect 60900 10892 77308 10948
rect 77364 10892 77374 10948
rect 38994 10780 39004 10836
rect 39060 10780 40292 10836
rect 59490 10780 59500 10836
rect 59556 10780 62076 10836
rect 62132 10780 76860 10836
rect 76916 10780 76926 10836
rect 50372 10668 50764 10724
rect 50820 10668 50830 10724
rect 69346 10668 69356 10724
rect 69412 10668 70252 10724
rect 70308 10668 70318 10724
rect 50372 10612 50428 10668
rect 40338 10556 40348 10612
rect 40404 10556 42476 10612
rect 42532 10556 42542 10612
rect 48066 10556 48076 10612
rect 48132 10556 50428 10612
rect 58258 10556 58268 10612
rect 58324 10556 70140 10612
rect 70196 10556 70206 10612
rect 71922 10556 71932 10612
rect 71988 10556 72828 10612
rect 72884 10556 72894 10612
rect 35522 10444 35532 10500
rect 35588 10444 36652 10500
rect 36708 10444 41468 10500
rect 41524 10444 43708 10500
rect 43764 10444 44828 10500
rect 44884 10444 45164 10500
rect 45220 10444 45230 10500
rect 48402 10444 48412 10500
rect 48468 10444 49756 10500
rect 49812 10444 49822 10500
rect 50866 10444 50876 10500
rect 50932 10444 52556 10500
rect 52612 10444 52622 10500
rect 54002 10444 54012 10500
rect 54068 10444 54684 10500
rect 54740 10444 54750 10500
rect 54898 10444 54908 10500
rect 54964 10444 65548 10500
rect 65604 10444 65614 10500
rect 68338 10444 68348 10500
rect 68404 10444 69132 10500
rect 69188 10444 69198 10500
rect 32274 10332 32284 10388
rect 32340 10332 33068 10388
rect 33124 10332 33134 10388
rect 35308 10332 37996 10388
rect 38052 10332 39452 10388
rect 39508 10332 39518 10388
rect 45612 10332 46956 10388
rect 47012 10332 47628 10388
rect 47684 10332 48748 10388
rect 48804 10332 48814 10388
rect 49298 10332 49308 10388
rect 49364 10332 50540 10388
rect 50596 10332 50606 10388
rect 62738 10332 62748 10388
rect 62804 10332 70700 10388
rect 70756 10332 70766 10388
rect 13570 10220 13580 10276
rect 13636 10220 22876 10276
rect 22932 10220 22942 10276
rect 25778 10220 25788 10276
rect 25844 10220 26460 10276
rect 26516 10220 26526 10276
rect 41234 10220 41244 10276
rect 41300 10220 45388 10276
rect 45444 10220 45454 10276
rect 30182 10164 30192 10220
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30456 10164 30466 10220
rect 45612 10164 45668 10332
rect 58146 10220 58156 10276
rect 58212 10220 66668 10276
rect 66724 10220 66734 10276
rect 49502 10164 49512 10220
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49776 10164 49786 10220
rect 68822 10164 68832 10220
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 69096 10164 69106 10220
rect 11228 10108 11788 10164
rect 13234 10108 13244 10164
rect 13300 10108 13310 10164
rect 16258 10108 16268 10164
rect 16324 10108 18172 10164
rect 18228 10108 18238 10164
rect 21298 10108 21308 10164
rect 21364 10108 21980 10164
rect 22036 10108 22046 10164
rect 25218 10108 25228 10164
rect 25284 10108 25900 10164
rect 25956 10108 25966 10164
rect 28018 10108 28028 10164
rect 28084 10108 29820 10164
rect 29876 10108 29886 10164
rect 39330 10108 39340 10164
rect 39396 10108 39406 10164
rect 40226 10108 40236 10164
rect 40292 10108 42028 10164
rect 42084 10108 42094 10164
rect 44818 10108 44828 10164
rect 44884 10108 45668 10164
rect 47058 10108 47068 10164
rect 47124 10108 49196 10164
rect 49252 10108 49262 10164
rect 51986 10108 51996 10164
rect 52052 10108 53004 10164
rect 53060 10108 53070 10164
rect 57474 10108 57484 10164
rect 57540 10108 63532 10164
rect 63588 10108 63598 10164
rect 11228 10052 11284 10108
rect 9538 9996 9548 10052
rect 9604 9996 11284 10052
rect 13244 10052 13300 10108
rect 13244 9996 15260 10052
rect 15316 9996 18732 10052
rect 18788 9996 20300 10052
rect 20356 9996 20972 10052
rect 21028 9996 21420 10052
rect 21476 9996 21868 10052
rect 21924 9996 23100 10052
rect 23156 9996 23166 10052
rect 24434 9996 24444 10052
rect 24500 9996 27916 10052
rect 27972 9996 27982 10052
rect 28690 9996 28700 10052
rect 28756 9996 30492 10052
rect 30548 9996 31500 10052
rect 31556 9996 31566 10052
rect 32162 9996 32172 10052
rect 32228 9996 34972 10052
rect 35028 9996 35038 10052
rect 35746 9996 35756 10052
rect 35812 9996 36428 10052
rect 36484 9996 37100 10052
rect 37156 9996 37166 10052
rect 39340 9940 39396 10108
rect 41010 9996 41020 10052
rect 41076 9996 41086 10052
rect 50418 9996 50428 10052
rect 50484 9996 51548 10052
rect 51604 9996 51614 10052
rect 66546 9996 66556 10052
rect 66612 9996 69244 10052
rect 69300 9996 69310 10052
rect 41020 9940 41076 9996
rect 15092 9884 26908 9940
rect 26964 9884 26974 9940
rect 27570 9884 27580 9940
rect 27636 9884 29932 9940
rect 29988 9884 29998 9940
rect 34402 9884 34412 9940
rect 34468 9884 35868 9940
rect 35924 9884 35934 9940
rect 37212 9884 39396 9940
rect 39554 9884 39564 9940
rect 39620 9884 41076 9940
rect 45378 9884 45388 9940
rect 45444 9884 49980 9940
rect 50036 9884 50820 9940
rect 51314 9884 51324 9940
rect 51380 9884 65212 9940
rect 65268 9884 65278 9940
rect 65436 9884 77532 9940
rect 77588 9884 77598 9940
rect 15092 9716 15148 9884
rect 26908 9828 26964 9884
rect 19852 9772 24444 9828
rect 24500 9772 24510 9828
rect 26908 9772 28140 9828
rect 28196 9772 32396 9828
rect 32452 9772 33292 9828
rect 33348 9772 33358 9828
rect 33506 9772 33516 9828
rect 33572 9772 36988 9828
rect 37044 9772 37054 9828
rect 11442 9660 11452 9716
rect 11508 9660 13356 9716
rect 13412 9660 15148 9716
rect 16146 9660 16156 9716
rect 16212 9660 17500 9716
rect 17556 9660 17566 9716
rect 11554 9548 11564 9604
rect 11620 9548 12908 9604
rect 12964 9548 12974 9604
rect 19852 9492 19908 9772
rect 37212 9716 37268 9884
rect 50764 9828 50820 9884
rect 65436 9828 65492 9884
rect 39218 9772 39228 9828
rect 39284 9772 39676 9828
rect 39732 9772 41020 9828
rect 41076 9772 41086 9828
rect 42354 9772 42364 9828
rect 42420 9772 47068 9828
rect 47124 9772 47134 9828
rect 50764 9772 53004 9828
rect 53060 9772 53070 9828
rect 54674 9772 54684 9828
rect 54740 9772 61180 9828
rect 61236 9772 61246 9828
rect 63074 9772 63084 9828
rect 63140 9772 65492 9828
rect 69794 9772 69804 9828
rect 69860 9772 70476 9828
rect 70532 9772 70542 9828
rect 71250 9772 71260 9828
rect 71316 9772 75852 9828
rect 75908 9772 75918 9828
rect 23762 9660 23772 9716
rect 23828 9660 34188 9716
rect 34244 9660 34254 9716
rect 37202 9660 37212 9716
rect 37268 9660 37278 9716
rect 40114 9660 40124 9716
rect 40180 9660 41692 9716
rect 41748 9660 41758 9716
rect 43138 9660 43148 9716
rect 43204 9660 43708 9716
rect 43764 9660 43774 9716
rect 48066 9660 48076 9716
rect 48132 9660 51996 9716
rect 52052 9660 52062 9716
rect 55020 9660 61292 9716
rect 61348 9660 61358 9716
rect 66770 9660 66780 9716
rect 66836 9660 67228 9716
rect 67284 9660 67294 9716
rect 75618 9660 75628 9716
rect 75684 9660 78428 9716
rect 78484 9660 78494 9716
rect 55020 9604 55076 9660
rect 20850 9548 20860 9604
rect 20916 9548 22876 9604
rect 22932 9548 22942 9604
rect 25778 9548 25788 9604
rect 25844 9548 26908 9604
rect 39442 9548 39452 9604
rect 39508 9548 40012 9604
rect 40068 9548 40908 9604
rect 40964 9548 40974 9604
rect 43362 9548 43372 9604
rect 43428 9548 44380 9604
rect 44436 9548 44446 9604
rect 48402 9548 48412 9604
rect 48468 9548 48860 9604
rect 48916 9548 48926 9604
rect 50372 9548 52668 9604
rect 52724 9548 52734 9604
rect 53666 9548 53676 9604
rect 53732 9548 55020 9604
rect 55076 9548 55086 9604
rect 58706 9548 58716 9604
rect 58772 9548 58940 9604
rect 58996 9548 60172 9604
rect 60228 9548 72380 9604
rect 72436 9548 72446 9604
rect 74498 9548 74508 9604
rect 74564 9548 74956 9604
rect 75012 9548 75022 9604
rect 6738 9436 6748 9492
rect 6804 9436 19852 9492
rect 19908 9436 19918 9492
rect 20522 9380 20532 9436
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20796 9380 20806 9436
rect 26852 9268 26908 9548
rect 48962 9436 48972 9492
rect 49028 9436 49308 9492
rect 49364 9436 49374 9492
rect 39842 9380 39852 9436
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 40116 9380 40126 9436
rect 50372 9380 50428 9548
rect 50530 9436 50540 9492
rect 50596 9436 52892 9492
rect 52948 9436 52958 9492
rect 64418 9436 64428 9492
rect 64484 9436 65324 9492
rect 65380 9436 65390 9492
rect 65660 9436 70588 9492
rect 71362 9436 71372 9492
rect 71428 9436 72604 9492
rect 72660 9436 72670 9492
rect 29372 9324 33740 9380
rect 33796 9324 33806 9380
rect 47618 9324 47628 9380
rect 47684 9324 50428 9380
rect 18834 9212 18844 9268
rect 18900 9212 20188 9268
rect 20244 9212 20254 9268
rect 22764 9212 23436 9268
rect 23492 9212 24220 9268
rect 24276 9212 24286 9268
rect 25330 9212 25340 9268
rect 25396 9212 26012 9268
rect 26068 9212 26078 9268
rect 26852 9212 28700 9268
rect 28756 9212 28766 9268
rect 22764 9156 22820 9212
rect 20066 9100 20076 9156
rect 20132 9100 22820 9156
rect 23090 9100 23100 9156
rect 23156 9100 24108 9156
rect 24164 9100 24174 9156
rect 25666 9100 25676 9156
rect 25732 9100 26348 9156
rect 26404 9100 26684 9156
rect 26740 9100 26750 9156
rect 29372 9044 29428 9324
rect 50540 9268 50596 9436
rect 59162 9380 59172 9436
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59436 9380 59446 9436
rect 65660 9380 65716 9436
rect 52546 9324 52556 9380
rect 52612 9324 55524 9380
rect 64194 9324 64204 9380
rect 64260 9324 65716 9380
rect 70532 9380 70588 9436
rect 78482 9380 78492 9436
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78756 9380 78766 9436
rect 70532 9324 71708 9380
rect 71764 9324 71774 9380
rect 55468 9268 55524 9324
rect 29586 9212 29596 9268
rect 29652 9212 33516 9268
rect 33572 9212 34636 9268
rect 34692 9212 36092 9268
rect 36148 9212 36158 9268
rect 49644 9212 50596 9268
rect 50978 9212 50988 9268
rect 51044 9212 53116 9268
rect 53172 9212 53182 9268
rect 55468 9212 64652 9268
rect 64708 9212 64718 9268
rect 65650 9212 65660 9268
rect 65716 9212 66108 9268
rect 66164 9212 66174 9268
rect 68796 9212 70532 9268
rect 71474 9212 71484 9268
rect 71540 9212 72268 9268
rect 72324 9212 72334 9268
rect 76626 9212 76636 9268
rect 76692 9212 77084 9268
rect 77140 9212 77150 9268
rect 49644 9156 49700 9212
rect 68796 9156 68852 9212
rect 31378 9100 31388 9156
rect 31444 9100 35532 9156
rect 35588 9100 35598 9156
rect 38098 9100 38108 9156
rect 38164 9100 40348 9156
rect 40404 9100 40414 9156
rect 43586 9100 43596 9156
rect 43652 9100 45836 9156
rect 45892 9100 45902 9156
rect 47730 9100 47740 9156
rect 47796 9100 48188 9156
rect 48244 9100 48860 9156
rect 48916 9100 49700 9156
rect 50642 9100 50652 9156
rect 50708 9100 55468 9156
rect 55524 9100 55534 9156
rect 58772 9100 67900 9156
rect 67956 9100 67966 9156
rect 68786 9100 68796 9156
rect 68852 9100 68862 9156
rect 69580 9100 70196 9156
rect 58772 9044 58828 9100
rect 69580 9044 69636 9100
rect 12114 8988 12124 9044
rect 12180 8988 14028 9044
rect 14084 8988 14094 9044
rect 23538 8988 23548 9044
rect 23604 8988 29428 9044
rect 31490 8988 31500 9044
rect 31556 8988 36316 9044
rect 36372 8988 36382 9044
rect 36642 8988 36652 9044
rect 36708 8988 37436 9044
rect 37492 8988 37502 9044
rect 38546 8988 38556 9044
rect 38612 8988 41804 9044
rect 41860 8988 41870 9044
rect 42690 8988 42700 9044
rect 42756 8988 49644 9044
rect 49700 8988 49710 9044
rect 50194 8988 50204 9044
rect 50260 8988 50764 9044
rect 50820 8988 50830 9044
rect 53890 8988 53900 9044
rect 53956 8988 54628 9044
rect 55346 8988 55356 9044
rect 55412 8988 58828 9044
rect 61394 8988 61404 9044
rect 61460 8988 62524 9044
rect 62580 8988 64988 9044
rect 65044 8988 65054 9044
rect 65538 8988 65548 9044
rect 65604 8988 65996 9044
rect 66052 8988 66062 9044
rect 69570 8988 69580 9044
rect 69636 8988 69646 9044
rect 12898 8876 12908 8932
rect 12964 8876 21028 8932
rect 21522 8876 21532 8932
rect 21588 8876 24220 8932
rect 24276 8876 24286 8932
rect 29810 8876 29820 8932
rect 29876 8876 31164 8932
rect 31220 8876 31230 8932
rect 31378 8876 31388 8932
rect 31444 8876 32620 8932
rect 32676 8876 32686 8932
rect 33394 8876 33404 8932
rect 33460 8876 34076 8932
rect 34132 8876 34142 8932
rect 35186 8876 35196 8932
rect 35252 8876 37212 8932
rect 37268 8876 37278 8932
rect 37538 8876 37548 8932
rect 37604 8876 38892 8932
rect 38948 8876 39228 8932
rect 39284 8876 39294 8932
rect 44706 8876 44716 8932
rect 44772 8876 45836 8932
rect 45892 8876 45902 8932
rect 47394 8876 47404 8932
rect 47460 8876 51548 8932
rect 51604 8876 51614 8932
rect 52210 8876 52220 8932
rect 52276 8876 54348 8932
rect 54404 8876 54414 8932
rect 20972 8820 21028 8876
rect 54572 8820 54628 8988
rect 56130 8876 56140 8932
rect 56196 8876 56588 8932
rect 56644 8876 56654 8932
rect 57138 8876 57148 8932
rect 57204 8876 57820 8932
rect 57876 8876 62300 8932
rect 62356 8876 62366 8932
rect 62850 8876 62860 8932
rect 62916 8876 62926 8932
rect 62860 8820 62916 8876
rect 70140 8820 70196 9100
rect 70476 9044 70532 9212
rect 71250 9100 71260 9156
rect 71316 9100 76860 9156
rect 76916 9100 76926 9156
rect 70476 8988 70588 9044
rect 70644 8988 70654 9044
rect 71138 8988 71148 9044
rect 71204 8988 77420 9044
rect 77476 8988 77486 9044
rect 70364 8876 72268 8932
rect 72324 8876 72334 8932
rect 72930 8876 72940 8932
rect 72996 8876 73006 8932
rect 70364 8820 70420 8876
rect 72940 8820 72996 8876
rect 9986 8764 9996 8820
rect 10052 8764 15148 8820
rect 20972 8764 22596 8820
rect 29474 8764 29484 8820
rect 29540 8764 30940 8820
rect 30996 8764 31006 8820
rect 31266 8764 31276 8820
rect 31332 8764 34860 8820
rect 34916 8764 37100 8820
rect 37156 8764 37996 8820
rect 38052 8764 38556 8820
rect 38612 8764 38622 8820
rect 41122 8764 41132 8820
rect 41188 8764 42028 8820
rect 42084 8764 42094 8820
rect 43474 8764 43484 8820
rect 43540 8764 49420 8820
rect 49476 8764 49486 8820
rect 49634 8764 49644 8820
rect 49700 8764 51100 8820
rect 51156 8764 51166 8820
rect 54572 8764 56756 8820
rect 59042 8764 59052 8820
rect 59108 8764 60060 8820
rect 60116 8764 60126 8820
rect 60722 8764 60732 8820
rect 60788 8764 62916 8820
rect 63186 8764 63196 8820
rect 63252 8764 65212 8820
rect 65268 8764 65278 8820
rect 65650 8764 65660 8820
rect 65716 8764 69860 8820
rect 70140 8764 70420 8820
rect 70532 8764 72996 8820
rect 73378 8764 73388 8820
rect 73444 8764 74508 8820
rect 74564 8764 74574 8820
rect 10862 8596 10872 8652
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 11136 8596 11146 8652
rect 15092 8596 15148 8764
rect 20860 8652 22316 8708
rect 22372 8652 22382 8708
rect 20860 8596 20916 8652
rect 15092 8540 20916 8596
rect 22540 8596 22596 8764
rect 56700 8708 56756 8764
rect 69804 8708 69860 8764
rect 22866 8652 22876 8708
rect 22932 8652 29708 8708
rect 29764 8652 29774 8708
rect 37538 8652 37548 8708
rect 37604 8652 41580 8708
rect 41636 8652 41646 8708
rect 44370 8652 44380 8708
rect 44436 8652 44940 8708
rect 44996 8652 45006 8708
rect 47170 8652 47180 8708
rect 47236 8652 47852 8708
rect 47908 8652 47918 8708
rect 50754 8652 50764 8708
rect 50820 8652 53564 8708
rect 53620 8652 53630 8708
rect 56690 8652 56700 8708
rect 56756 8652 56766 8708
rect 59714 8652 59724 8708
rect 59780 8652 60396 8708
rect 60452 8652 60462 8708
rect 61282 8652 61292 8708
rect 61348 8652 68628 8708
rect 69804 8652 70252 8708
rect 70308 8652 70318 8708
rect 30182 8596 30192 8652
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30456 8596 30466 8652
rect 49502 8596 49512 8652
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49776 8596 49786 8652
rect 22540 8540 29036 8596
rect 29092 8540 29596 8596
rect 29652 8540 29662 8596
rect 36306 8540 36316 8596
rect 36372 8540 38108 8596
rect 38164 8540 38174 8596
rect 43810 8540 43820 8596
rect 43876 8540 45276 8596
rect 45332 8540 45342 8596
rect 47954 8540 47964 8596
rect 48020 8540 48636 8596
rect 48692 8540 48702 8596
rect 48962 8540 48972 8596
rect 49028 8540 49308 8596
rect 49364 8540 49374 8596
rect 49970 8540 49980 8596
rect 50036 8540 51548 8596
rect 51604 8540 51614 8596
rect 54562 8540 54572 8596
rect 54628 8540 66668 8596
rect 66724 8540 66734 8596
rect 67890 8540 67900 8596
rect 67956 8540 68348 8596
rect 68404 8540 68414 8596
rect 13570 8428 13580 8484
rect 13636 8428 19908 8484
rect 24994 8428 25004 8484
rect 25060 8428 31948 8484
rect 32004 8428 32014 8484
rect 34402 8428 34412 8484
rect 34468 8428 51100 8484
rect 51156 8428 51166 8484
rect 52210 8428 52220 8484
rect 52276 8428 59948 8484
rect 60004 8428 60014 8484
rect 61170 8428 61180 8484
rect 61236 8428 61740 8484
rect 61796 8428 61806 8484
rect 62290 8428 62300 8484
rect 62356 8428 62636 8484
rect 62692 8428 63532 8484
rect 63588 8428 63598 8484
rect 63858 8428 63868 8484
rect 63924 8428 64652 8484
rect 64708 8428 64718 8484
rect 64866 8428 64876 8484
rect 64932 8428 65324 8484
rect 65380 8428 65390 8484
rect 19852 8372 19908 8428
rect 68572 8372 68628 8652
rect 68822 8596 68832 8652
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 69096 8596 69106 8652
rect 69570 8540 69580 8596
rect 69636 8540 70140 8596
rect 70196 8540 70206 8596
rect 70532 8372 70588 8764
rect 71026 8652 71036 8708
rect 71092 8652 76188 8708
rect 76244 8652 76254 8708
rect 71698 8540 71708 8596
rect 71764 8540 71932 8596
rect 71988 8540 73276 8596
rect 73332 8540 73342 8596
rect 71026 8428 71036 8484
rect 71092 8428 73724 8484
rect 73780 8428 73790 8484
rect 8530 8316 8540 8372
rect 8596 8316 19684 8372
rect 19852 8316 21476 8372
rect 21634 8316 21644 8372
rect 21700 8316 23660 8372
rect 23716 8316 23884 8372
rect 23940 8316 23950 8372
rect 25106 8316 25116 8372
rect 25172 8316 27132 8372
rect 27188 8316 27198 8372
rect 27906 8316 27916 8372
rect 27972 8316 28924 8372
rect 28980 8316 28990 8372
rect 30044 8316 33628 8372
rect 33684 8316 33694 8372
rect 34178 8316 34188 8372
rect 34244 8316 35868 8372
rect 35924 8316 35934 8372
rect 37426 8316 37436 8372
rect 37492 8316 39452 8372
rect 39508 8316 39518 8372
rect 39890 8316 39900 8372
rect 39956 8316 41020 8372
rect 41076 8316 41086 8372
rect 41346 8316 41356 8372
rect 41412 8316 46844 8372
rect 46900 8316 46910 8372
rect 48402 8316 48412 8372
rect 48468 8316 48748 8372
rect 48804 8316 48814 8372
rect 49298 8316 49308 8372
rect 49364 8316 50092 8372
rect 50148 8316 50158 8372
rect 52322 8316 52332 8372
rect 52388 8316 53788 8372
rect 53844 8316 53854 8372
rect 58482 8316 58492 8372
rect 58548 8316 63644 8372
rect 63700 8316 65996 8372
rect 66052 8316 66062 8372
rect 66322 8316 66332 8372
rect 66388 8316 66398 8372
rect 66882 8316 66892 8372
rect 66948 8316 68348 8372
rect 68404 8316 68414 8372
rect 68572 8316 70588 8372
rect 72034 8316 72044 8372
rect 72100 8316 72110 8372
rect 73154 8316 73164 8372
rect 73220 8316 78092 8372
rect 78148 8316 78158 8372
rect 19628 8260 19684 8316
rect 21420 8260 21476 8316
rect 9874 8204 9884 8260
rect 9940 8204 10332 8260
rect 10388 8204 10398 8260
rect 15362 8204 15372 8260
rect 15428 8204 17500 8260
rect 17556 8204 19572 8260
rect 19628 8204 21028 8260
rect 21420 8204 21868 8260
rect 21924 8204 21934 8260
rect 22082 8204 22092 8260
rect 22148 8204 22158 8260
rect 22754 8204 22764 8260
rect 22820 8204 24332 8260
rect 24388 8204 24398 8260
rect 24658 8204 24668 8260
rect 24724 8204 27244 8260
rect 27300 8204 27310 8260
rect 27682 8204 27692 8260
rect 27748 8204 28364 8260
rect 28420 8204 28430 8260
rect 19516 8148 19572 8204
rect 13794 8092 13804 8148
rect 13860 8092 15932 8148
rect 15988 8092 15998 8148
rect 16370 8092 16380 8148
rect 16436 8092 16604 8148
rect 16660 8092 17388 8148
rect 17444 8092 17454 8148
rect 19506 8092 19516 8148
rect 19572 8092 19582 8148
rect 14578 7980 14588 8036
rect 14644 7980 15260 8036
rect 15316 7980 15326 8036
rect 20522 7812 20532 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20796 7812 20806 7868
rect 20972 7812 21028 8204
rect 22092 8036 22148 8204
rect 30044 8148 30100 8316
rect 66332 8260 66388 8316
rect 30594 8204 30604 8260
rect 30660 8204 34412 8260
rect 34468 8204 34478 8260
rect 40898 8204 40908 8260
rect 40964 8204 45164 8260
rect 45220 8204 46732 8260
rect 46788 8204 50428 8260
rect 50484 8204 50494 8260
rect 51874 8204 51884 8260
rect 51940 8204 54796 8260
rect 54852 8204 54862 8260
rect 55794 8204 55804 8260
rect 55860 8204 59724 8260
rect 59780 8204 59790 8260
rect 61842 8204 61852 8260
rect 61908 8204 62188 8260
rect 62244 8204 62254 8260
rect 62514 8204 62524 8260
rect 62580 8204 63532 8260
rect 63588 8204 63598 8260
rect 63858 8204 63868 8260
rect 63924 8204 63934 8260
rect 64978 8204 64988 8260
rect 65044 8204 65548 8260
rect 65604 8204 65614 8260
rect 65874 8204 65884 8260
rect 65940 8204 66388 8260
rect 66546 8204 66556 8260
rect 66612 8204 67228 8260
rect 67284 8204 67294 8260
rect 68226 8204 68236 8260
rect 68292 8204 70140 8260
rect 70196 8204 70206 8260
rect 63868 8148 63924 8204
rect 72044 8148 72100 8316
rect 21634 7980 21644 8036
rect 21700 7980 22148 8036
rect 22316 8092 24108 8148
rect 24164 8092 24174 8148
rect 26786 8092 26796 8148
rect 26852 8092 27020 8148
rect 27076 8092 27086 8148
rect 28130 8092 28140 8148
rect 28196 8092 30100 8148
rect 32498 8092 32508 8148
rect 32564 8092 33516 8148
rect 33572 8092 33582 8148
rect 37202 8092 37212 8148
rect 37268 8092 37884 8148
rect 37940 8092 37950 8148
rect 38668 8092 39228 8148
rect 39284 8092 41748 8148
rect 44146 8092 44156 8148
rect 44212 8092 45836 8148
rect 45892 8092 45902 8148
rect 46610 8092 46620 8148
rect 46676 8092 47180 8148
rect 47236 8092 47246 8148
rect 47842 8092 47852 8148
rect 47908 8092 49644 8148
rect 49700 8092 49710 8148
rect 52994 8092 53004 8148
rect 53060 8092 55244 8148
rect 55300 8092 55310 8148
rect 56018 8092 56028 8148
rect 56084 8092 60732 8148
rect 60788 8092 60798 8148
rect 62412 8092 64092 8148
rect 64148 8092 65604 8148
rect 68114 8092 68124 8148
rect 68180 8092 68908 8148
rect 68964 8092 69356 8148
rect 69412 8092 69422 8148
rect 72044 8092 76188 8148
rect 76244 8092 76254 8148
rect 21298 7868 21308 7924
rect 21364 7868 21756 7924
rect 21812 7868 21822 7924
rect 22316 7812 22372 8092
rect 38668 8036 38724 8092
rect 41692 8036 41748 8092
rect 20972 7756 22372 7812
rect 23492 7980 27692 8036
rect 27748 7980 30268 8036
rect 30324 7980 31612 8036
rect 31668 7980 31678 8036
rect 33058 7980 33068 8036
rect 33124 7980 34412 8036
rect 34468 7980 34478 8036
rect 38658 7980 38668 8036
rect 38724 7980 38734 8036
rect 39330 7980 39340 8036
rect 39396 7980 39676 8036
rect 39732 7980 39742 8036
rect 41692 7980 44044 8036
rect 44100 7980 44110 8036
rect 44594 7980 44604 8036
rect 44660 7980 45052 8036
rect 45108 7980 45118 8036
rect 46386 7980 46396 8036
rect 46452 7980 48636 8036
rect 48692 7980 48702 8036
rect 49970 7980 49980 8036
rect 50036 7980 51324 8036
rect 51380 7980 51390 8036
rect 51874 7980 51884 8036
rect 51940 7980 52556 8036
rect 52612 7980 52622 8036
rect 53778 7980 53788 8036
rect 53844 7980 55916 8036
rect 55972 7980 55982 8036
rect 56252 7980 62188 8036
rect 62244 7980 62254 8036
rect 23492 7700 23548 7980
rect 24322 7868 24332 7924
rect 24388 7868 26796 7924
rect 26852 7868 29484 7924
rect 29540 7868 29550 7924
rect 30034 7868 30044 7924
rect 30100 7868 34860 7924
rect 34916 7868 34926 7924
rect 41346 7868 41356 7924
rect 41412 7868 42700 7924
rect 42756 7868 42766 7924
rect 43820 7868 55804 7924
rect 55860 7868 55870 7924
rect 39842 7812 39852 7868
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 40116 7812 40126 7868
rect 43820 7812 43876 7868
rect 56252 7812 56308 7980
rect 62412 7924 62468 8092
rect 64204 7980 65324 8036
rect 65380 7980 65390 8036
rect 60722 7868 60732 7924
rect 60788 7868 62468 7924
rect 63644 7868 63980 7924
rect 64036 7868 64046 7924
rect 59162 7812 59172 7868
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59436 7812 59446 7868
rect 27234 7756 27244 7812
rect 27300 7756 28924 7812
rect 28980 7756 28990 7812
rect 33180 7756 38444 7812
rect 38500 7756 38510 7812
rect 42242 7756 42252 7812
rect 42308 7756 43820 7812
rect 43876 7756 43886 7812
rect 44258 7756 44268 7812
rect 44324 7756 56308 7812
rect 58930 7756 58940 7812
rect 58996 7756 59006 7812
rect 60834 7756 60844 7812
rect 60900 7756 61180 7812
rect 61236 7756 61246 7812
rect 10434 7644 10444 7700
rect 10500 7644 11788 7700
rect 11844 7644 13468 7700
rect 13524 7644 13534 7700
rect 17714 7644 17724 7700
rect 17780 7644 19852 7700
rect 19908 7644 21756 7700
rect 21812 7644 23548 7700
rect 25676 7644 26348 7700
rect 26404 7644 26414 7700
rect 26562 7644 26572 7700
rect 26628 7644 27020 7700
rect 27076 7644 27086 7700
rect 29810 7644 29820 7700
rect 29876 7644 30716 7700
rect 30772 7644 30782 7700
rect 6066 7532 6076 7588
rect 6132 7532 22876 7588
rect 22932 7532 22942 7588
rect 23874 7532 23884 7588
rect 23940 7532 24220 7588
rect 24276 7532 24286 7588
rect 25676 7476 25732 7644
rect 25890 7532 25900 7588
rect 25956 7532 27244 7588
rect 27300 7532 27310 7588
rect 15250 7420 15260 7476
rect 15316 7420 18172 7476
rect 18228 7420 19516 7476
rect 19572 7420 19582 7476
rect 24098 7420 24108 7476
rect 24164 7420 25732 7476
rect 26002 7420 26012 7476
rect 26068 7420 27692 7476
rect 27748 7420 27758 7476
rect 25676 7364 25732 7420
rect 33180 7364 33236 7756
rect 33618 7644 33628 7700
rect 33684 7644 35084 7700
rect 35140 7644 35150 7700
rect 35858 7644 35868 7700
rect 35924 7644 38556 7700
rect 38612 7644 38622 7700
rect 40338 7644 40348 7700
rect 40404 7644 41580 7700
rect 41636 7644 41646 7700
rect 42466 7644 42476 7700
rect 42532 7644 44716 7700
rect 44772 7644 44782 7700
rect 45042 7644 45052 7700
rect 45108 7644 46396 7700
rect 46452 7644 46462 7700
rect 47058 7644 47068 7700
rect 47124 7644 48076 7700
rect 48132 7644 48142 7700
rect 48962 7644 48972 7700
rect 49028 7644 50652 7700
rect 50708 7644 50718 7700
rect 51986 7644 51996 7700
rect 52052 7644 53228 7700
rect 53284 7644 54348 7700
rect 54404 7644 54414 7700
rect 54786 7644 54796 7700
rect 54852 7644 55468 7700
rect 55524 7644 56588 7700
rect 56644 7644 56654 7700
rect 38882 7532 38892 7588
rect 38948 7532 41132 7588
rect 41188 7532 41198 7588
rect 42802 7532 42812 7588
rect 42868 7532 45724 7588
rect 45780 7532 45790 7588
rect 47282 7532 47292 7588
rect 47348 7532 48748 7588
rect 48804 7532 48814 7588
rect 49522 7532 49532 7588
rect 49588 7532 49868 7588
rect 49924 7532 49934 7588
rect 53732 7532 56700 7588
rect 56756 7532 56766 7588
rect 56914 7532 56924 7588
rect 56980 7532 58380 7588
rect 58436 7532 58446 7588
rect 53732 7476 53788 7532
rect 34402 7420 34412 7476
rect 34468 7420 36204 7476
rect 36260 7420 36764 7476
rect 36820 7420 36830 7476
rect 37874 7420 37884 7476
rect 37940 7420 39900 7476
rect 39956 7420 40908 7476
rect 40964 7420 40974 7476
rect 41682 7420 41692 7476
rect 41748 7420 44380 7476
rect 44436 7420 44446 7476
rect 47618 7420 47628 7476
rect 47684 7420 49084 7476
rect 49140 7420 50092 7476
rect 50148 7420 53788 7476
rect 55794 7420 55804 7476
rect 55860 7420 57036 7476
rect 57092 7420 57484 7476
rect 57540 7420 57550 7476
rect 58940 7364 58996 7756
rect 63644 7700 63700 7868
rect 64204 7812 64260 7980
rect 65548 7924 65604 8092
rect 67778 7980 67788 8036
rect 67844 7980 68348 8036
rect 68404 7980 68414 8036
rect 70532 7980 73220 8036
rect 73378 7980 73388 8036
rect 73444 7980 77980 8036
rect 78036 7980 78046 8036
rect 70532 7924 70588 7980
rect 65548 7868 70588 7924
rect 73164 7924 73220 7980
rect 73164 7868 77084 7924
rect 77140 7868 77150 7924
rect 78482 7812 78492 7868
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78756 7812 78766 7868
rect 63858 7756 63868 7812
rect 63924 7756 64260 7812
rect 65538 7756 65548 7812
rect 65604 7756 65884 7812
rect 65940 7756 65950 7812
rect 66882 7756 66892 7812
rect 66948 7756 70588 7812
rect 59388 7644 60732 7700
rect 60788 7644 60798 7700
rect 62178 7644 62188 7700
rect 62244 7644 64484 7700
rect 59388 7588 59444 7644
rect 64428 7588 64484 7644
rect 65772 7644 66668 7700
rect 66724 7644 66734 7700
rect 68450 7644 68460 7700
rect 68516 7644 68526 7700
rect 65772 7588 65828 7644
rect 59266 7532 59276 7588
rect 59332 7532 59444 7588
rect 61506 7532 61516 7588
rect 61572 7532 62524 7588
rect 62580 7532 62590 7588
rect 62850 7532 62860 7588
rect 62916 7532 64204 7588
rect 64260 7532 64270 7588
rect 64428 7532 65828 7588
rect 65986 7532 65996 7588
rect 66052 7532 66556 7588
rect 66612 7532 67340 7588
rect 67396 7532 67406 7588
rect 67890 7532 67900 7588
rect 67956 7532 68236 7588
rect 68292 7532 68302 7588
rect 68460 7476 68516 7644
rect 70532 7588 70588 7756
rect 70690 7644 70700 7700
rect 70756 7644 72604 7700
rect 72660 7644 72670 7700
rect 70532 7532 76860 7588
rect 76916 7532 76926 7588
rect 61730 7420 61740 7476
rect 61796 7420 64540 7476
rect 64596 7420 64606 7476
rect 64978 7420 64988 7476
rect 65044 7420 70028 7476
rect 70084 7420 70094 7476
rect 71138 7420 71148 7476
rect 71204 7420 72604 7476
rect 72660 7420 72670 7476
rect 75618 7420 75628 7476
rect 75684 7420 77980 7476
rect 78036 7420 78046 7476
rect 5842 7308 5852 7364
rect 5908 7308 6524 7364
rect 6580 7308 6590 7364
rect 16818 7308 16828 7364
rect 16884 7308 18844 7364
rect 18900 7308 18910 7364
rect 19618 7308 19628 7364
rect 19684 7308 20076 7364
rect 20132 7308 20142 7364
rect 21522 7308 21532 7364
rect 21588 7308 22988 7364
rect 23044 7308 23054 7364
rect 25676 7308 26460 7364
rect 26516 7308 26526 7364
rect 27356 7308 32340 7364
rect 33170 7308 33180 7364
rect 33236 7308 33246 7364
rect 37762 7308 37772 7364
rect 37828 7308 38220 7364
rect 38276 7308 38286 7364
rect 40338 7308 40348 7364
rect 40404 7308 41132 7364
rect 41188 7308 41198 7364
rect 42354 7308 42364 7364
rect 42420 7308 43148 7364
rect 43204 7308 43596 7364
rect 43652 7308 43662 7364
rect 44034 7308 44044 7364
rect 44100 7308 49756 7364
rect 49812 7308 49822 7364
rect 50754 7308 50764 7364
rect 50820 7308 51324 7364
rect 51380 7308 51390 7364
rect 51762 7308 51772 7364
rect 51828 7308 58492 7364
rect 58548 7308 58558 7364
rect 58940 7308 59276 7364
rect 59332 7308 59342 7364
rect 59938 7308 59948 7364
rect 60004 7308 61516 7364
rect 61572 7308 61582 7364
rect 62178 7308 62188 7364
rect 62244 7308 63532 7364
rect 63588 7308 63598 7364
rect 64418 7308 64428 7364
rect 64484 7308 65884 7364
rect 65940 7308 66668 7364
rect 66724 7308 66734 7364
rect 67106 7308 67116 7364
rect 67172 7308 69020 7364
rect 69076 7308 69086 7364
rect 71922 7308 71932 7364
rect 71988 7308 73276 7364
rect 73332 7308 73342 7364
rect 73714 7308 73724 7364
rect 73780 7308 78092 7364
rect 78148 7308 78158 7364
rect 27356 7252 27412 7308
rect 32284 7252 32340 7308
rect 19628 7196 24556 7252
rect 24612 7196 24622 7252
rect 24892 7196 25900 7252
rect 25956 7196 25966 7252
rect 27346 7196 27356 7252
rect 27412 7196 27422 7252
rect 27570 7196 27580 7252
rect 27636 7196 27916 7252
rect 27972 7196 27982 7252
rect 29596 7196 32060 7252
rect 32116 7196 32126 7252
rect 32284 7196 57932 7252
rect 57988 7196 57998 7252
rect 58370 7196 58380 7252
rect 58436 7196 59052 7252
rect 59108 7196 59118 7252
rect 60946 7196 60956 7252
rect 61012 7196 63420 7252
rect 63476 7196 63486 7252
rect 66210 7196 66220 7252
rect 66276 7196 67340 7252
rect 67396 7196 67406 7252
rect 68684 7196 68908 7252
rect 68964 7196 68974 7252
rect 71138 7196 71148 7252
rect 71204 7196 72380 7252
rect 72436 7196 72446 7252
rect 77532 7196 77756 7252
rect 77812 7196 77822 7252
rect 19628 7140 19684 7196
rect 24892 7140 24948 7196
rect 19618 7084 19628 7140
rect 19684 7084 19694 7140
rect 22866 7084 22876 7140
rect 22932 7084 23212 7140
rect 23268 7084 23278 7140
rect 23986 7084 23996 7140
rect 24052 7084 24948 7140
rect 25554 7084 25564 7140
rect 25620 7084 28140 7140
rect 28196 7084 28206 7140
rect 28466 7084 28476 7140
rect 28532 7084 29036 7140
rect 29092 7084 29102 7140
rect 10862 7028 10872 7084
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 11136 7028 11146 7084
rect 29596 7028 29652 7196
rect 68684 7140 68740 7196
rect 77532 7140 77588 7196
rect 30594 7084 30604 7140
rect 30660 7084 38668 7140
rect 38882 7084 38892 7140
rect 38948 7084 39452 7140
rect 39508 7084 39518 7140
rect 42466 7084 42476 7140
rect 42532 7084 43036 7140
rect 43092 7084 48188 7140
rect 48244 7084 48254 7140
rect 48626 7084 48636 7140
rect 48692 7084 49252 7140
rect 57250 7084 57260 7140
rect 57316 7084 59724 7140
rect 59780 7084 59790 7140
rect 62178 7084 62188 7140
rect 62244 7084 62748 7140
rect 62804 7084 62814 7140
rect 64866 7084 64876 7140
rect 64932 7084 66332 7140
rect 66388 7084 66398 7140
rect 66882 7084 66892 7140
rect 66948 7084 68740 7140
rect 69244 7084 69916 7140
rect 69972 7084 71260 7140
rect 71316 7084 71326 7140
rect 72818 7084 72828 7140
rect 72884 7084 73724 7140
rect 73780 7084 73790 7140
rect 77522 7084 77532 7140
rect 77588 7084 77598 7140
rect 30182 7028 30192 7084
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30456 7028 30466 7084
rect 11228 6972 12740 7028
rect 14354 6972 14364 7028
rect 14420 6972 15036 7028
rect 15092 6972 29596 7028
rect 29652 6972 29662 7028
rect 11228 6916 11284 6972
rect 12684 6916 12740 6972
rect 38612 6916 38668 7084
rect 42578 6972 42588 7028
rect 42644 6972 44268 7028
rect 44324 6972 44334 7028
rect 44706 6972 44716 7028
rect 44772 6972 46508 7028
rect 46564 6972 46574 7028
rect 49196 6916 49252 7084
rect 49502 7028 49512 7084
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49776 7028 49786 7084
rect 66332 7028 66388 7084
rect 68822 7028 68832 7084
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 69096 7028 69106 7084
rect 56018 6972 56028 7028
rect 56084 6972 56588 7028
rect 56644 6972 56654 7028
rect 57092 6972 59612 7028
rect 59668 6972 59678 7028
rect 59938 6972 59948 7028
rect 60004 6972 61068 7028
rect 61124 6972 61134 7028
rect 61730 6972 61740 7028
rect 61796 6972 63868 7028
rect 63924 6972 63934 7028
rect 66332 6972 66556 7028
rect 66612 6972 66622 7028
rect 67890 6972 67900 7028
rect 67956 6972 68572 7028
rect 68628 6972 68638 7028
rect 57092 6916 57148 6972
rect 69244 6916 69300 7084
rect 69794 6972 69804 7028
rect 69860 6972 76972 7028
rect 77028 6972 77038 7028
rect 5058 6860 5068 6916
rect 5124 6860 11284 6916
rect 12450 6860 12460 6916
rect 12516 6860 12526 6916
rect 12684 6860 21980 6916
rect 22036 6860 22046 6916
rect 24210 6860 24220 6916
rect 24276 6860 24556 6916
rect 24612 6860 24622 6916
rect 28018 6860 28028 6916
rect 28084 6860 28364 6916
rect 28420 6860 28430 6916
rect 28578 6860 28588 6916
rect 28644 6860 38220 6916
rect 38276 6860 38286 6916
rect 38612 6860 47516 6916
rect 47572 6860 47582 6916
rect 47842 6860 47852 6916
rect 47908 6860 47918 6916
rect 49196 6860 52332 6916
rect 52388 6860 52398 6916
rect 54450 6860 54460 6916
rect 54516 6860 56364 6916
rect 56420 6860 56430 6916
rect 56914 6860 56924 6916
rect 56980 6860 57148 6916
rect 59052 6860 61516 6916
rect 61572 6860 61582 6916
rect 62132 6860 63756 6916
rect 63812 6860 63822 6916
rect 64194 6860 64204 6916
rect 64260 6860 69300 6916
rect 70018 6860 70028 6916
rect 70084 6860 75516 6916
rect 75572 6860 75582 6916
rect 6514 6748 6524 6804
rect 6580 6748 9436 6804
rect 9492 6748 9502 6804
rect 12460 6692 12516 6860
rect 47852 6804 47908 6860
rect 59052 6804 59108 6860
rect 62132 6804 62188 6860
rect 16594 6748 16604 6804
rect 16660 6748 17276 6804
rect 17332 6748 19292 6804
rect 19348 6748 19358 6804
rect 20514 6748 20524 6804
rect 20580 6748 22092 6804
rect 22148 6748 22158 6804
rect 24434 6748 24444 6804
rect 24500 6748 25228 6804
rect 25284 6748 25294 6804
rect 27580 6748 29372 6804
rect 29428 6748 29438 6804
rect 33842 6748 33852 6804
rect 33908 6748 40012 6804
rect 40068 6748 40078 6804
rect 41010 6748 41020 6804
rect 41076 6748 44044 6804
rect 44100 6748 44110 6804
rect 47852 6748 49028 6804
rect 52098 6748 52108 6804
rect 52164 6748 59108 6804
rect 59266 6748 59276 6804
rect 59332 6748 60060 6804
rect 60116 6748 60126 6804
rect 60284 6748 62188 6804
rect 62290 6748 62300 6804
rect 62356 6748 63420 6804
rect 63476 6748 63486 6804
rect 63634 6748 63644 6804
rect 63700 6748 64428 6804
rect 64484 6748 64494 6804
rect 65426 6748 65436 6804
rect 65492 6748 71484 6804
rect 71540 6748 71550 6804
rect 72818 6748 72828 6804
rect 72884 6748 77084 6804
rect 77140 6748 77150 6804
rect 27580 6692 27636 6748
rect 5964 6636 6300 6692
rect 6356 6636 6366 6692
rect 6626 6636 6636 6692
rect 6692 6636 7756 6692
rect 7812 6636 7822 6692
rect 12460 6636 14700 6692
rect 14756 6636 14766 6692
rect 20402 6636 20412 6692
rect 20468 6636 21756 6692
rect 21812 6636 21822 6692
rect 26562 6636 26572 6692
rect 26628 6636 26638 6692
rect 26786 6636 26796 6692
rect 26852 6636 27636 6692
rect 27794 6636 27804 6692
rect 27860 6636 28028 6692
rect 28084 6636 33292 6692
rect 33348 6636 34972 6692
rect 35028 6636 35038 6692
rect 36306 6636 36316 6692
rect 36372 6636 37996 6692
rect 38052 6636 39788 6692
rect 39844 6636 41804 6692
rect 41860 6636 41870 6692
rect 42130 6636 42140 6692
rect 42196 6636 42812 6692
rect 42868 6636 42878 6692
rect 44146 6636 44156 6692
rect 44212 6636 46396 6692
rect 46452 6636 46462 6692
rect 5964 6468 6020 6636
rect 26572 6580 26628 6636
rect 7074 6524 7084 6580
rect 7140 6524 9212 6580
rect 9268 6524 9884 6580
rect 9940 6524 9950 6580
rect 13122 6524 13132 6580
rect 13188 6524 13692 6580
rect 13748 6524 13758 6580
rect 14252 6524 22988 6580
rect 23044 6524 23436 6580
rect 23492 6524 29372 6580
rect 29428 6524 29438 6580
rect 35252 6524 35980 6580
rect 36036 6524 36428 6580
rect 36484 6524 36494 6580
rect 37762 6524 37772 6580
rect 37828 6524 41580 6580
rect 41636 6524 41646 6580
rect 43698 6524 43708 6580
rect 43764 6524 44604 6580
rect 44660 6524 44670 6580
rect 45490 6524 45500 6580
rect 45556 6524 48636 6580
rect 48692 6524 48702 6580
rect 5964 6412 9660 6468
rect 9716 6412 9726 6468
rect 14252 6356 14308 6524
rect 35252 6468 35308 6524
rect 48972 6468 49028 6748
rect 50642 6636 50652 6692
rect 50708 6636 50988 6692
rect 51044 6636 51054 6692
rect 51538 6636 51548 6692
rect 51604 6636 53900 6692
rect 53956 6636 53966 6692
rect 58930 6636 58940 6692
rect 58996 6636 59948 6692
rect 60004 6636 60014 6692
rect 60284 6580 60340 6748
rect 63074 6636 63084 6692
rect 63140 6636 64876 6692
rect 64932 6636 64942 6692
rect 67442 6636 67452 6692
rect 67508 6636 67788 6692
rect 67844 6636 67854 6692
rect 72370 6636 72380 6692
rect 72436 6636 72716 6692
rect 72772 6636 72782 6692
rect 73154 6636 73164 6692
rect 73220 6636 73612 6692
rect 73668 6636 73678 6692
rect 49186 6524 49196 6580
rect 49252 6524 60340 6580
rect 60722 6524 60732 6580
rect 60788 6524 61852 6580
rect 61908 6524 61918 6580
rect 62402 6524 62412 6580
rect 62468 6524 62972 6580
rect 63028 6524 64540 6580
rect 64596 6524 64606 6580
rect 67106 6524 67116 6580
rect 67172 6524 68572 6580
rect 68628 6524 68638 6580
rect 69916 6524 74172 6580
rect 74228 6524 74238 6580
rect 75730 6524 75740 6580
rect 75796 6524 76300 6580
rect 76356 6524 76366 6580
rect 69916 6468 69972 6524
rect 14466 6412 14476 6468
rect 14532 6412 16716 6468
rect 16772 6412 16782 6468
rect 23314 6412 23324 6468
rect 23380 6412 25900 6468
rect 25956 6412 25966 6468
rect 26898 6412 26908 6468
rect 26964 6412 29260 6468
rect 29316 6412 35308 6468
rect 39330 6412 39340 6468
rect 39396 6412 42028 6468
rect 42084 6412 42094 6468
rect 42802 6412 42812 6468
rect 42868 6412 43372 6468
rect 43428 6412 43438 6468
rect 44034 6412 44044 6468
rect 44100 6412 47068 6468
rect 47124 6412 47134 6468
rect 48972 6412 50428 6468
rect 50978 6412 50988 6468
rect 51044 6412 51772 6468
rect 51828 6412 51838 6468
rect 54460 6412 58380 6468
rect 58436 6412 58446 6468
rect 60172 6412 61740 6468
rect 61796 6412 61806 6468
rect 62514 6412 62524 6468
rect 62580 6412 63308 6468
rect 63364 6412 63374 6468
rect 63746 6412 63756 6468
rect 63812 6412 64316 6468
rect 64372 6412 64382 6468
rect 65650 6412 65660 6468
rect 65716 6412 66780 6468
rect 66836 6412 66846 6468
rect 68226 6412 68236 6468
rect 68292 6412 69972 6468
rect 73892 6412 77980 6468
rect 78036 6412 78046 6468
rect 50372 6356 50428 6412
rect 54460 6356 54516 6412
rect 60172 6356 60228 6412
rect 73892 6356 73948 6412
rect 7074 6300 7084 6356
rect 7140 6300 8652 6356
rect 8708 6300 8718 6356
rect 9538 6300 9548 6356
rect 9604 6300 11452 6356
rect 11508 6300 11518 6356
rect 11732 6300 14308 6356
rect 15092 6300 16156 6356
rect 16212 6300 16222 6356
rect 16818 6300 16828 6356
rect 16884 6300 17388 6356
rect 17444 6300 19292 6356
rect 19348 6300 19358 6356
rect 21858 6300 21868 6356
rect 21924 6300 21934 6356
rect 22306 6300 22316 6356
rect 22372 6300 22988 6356
rect 23044 6300 23054 6356
rect 24658 6300 24668 6356
rect 24724 6300 25116 6356
rect 25172 6300 25182 6356
rect 25330 6300 25340 6356
rect 25396 6300 25406 6356
rect 25666 6300 25676 6356
rect 25732 6300 26796 6356
rect 26852 6300 26862 6356
rect 27346 6300 27356 6356
rect 27412 6300 28588 6356
rect 28644 6300 28654 6356
rect 43708 6300 45724 6356
rect 45780 6300 45790 6356
rect 46386 6300 46396 6356
rect 46452 6300 46788 6356
rect 46946 6300 46956 6356
rect 47012 6300 49196 6356
rect 49252 6300 49262 6356
rect 50372 6300 54516 6356
rect 59602 6300 59612 6356
rect 59668 6300 60228 6356
rect 61954 6300 61964 6356
rect 62020 6300 62580 6356
rect 62738 6300 62748 6356
rect 62804 6300 63644 6356
rect 63700 6300 63710 6356
rect 63858 6300 63868 6356
rect 63924 6300 65100 6356
rect 65156 6300 67452 6356
rect 67508 6300 67518 6356
rect 73500 6300 73948 6356
rect 11732 6244 11788 6300
rect 6066 6188 6076 6244
rect 6132 6188 7196 6244
rect 7252 6188 7262 6244
rect 7634 6188 7644 6244
rect 7700 6188 9996 6244
rect 10052 6188 11788 6244
rect 15092 6132 15148 6300
rect 20522 6244 20532 6300
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20796 6244 20806 6300
rect 21868 6244 21924 6300
rect 25340 6244 25396 6300
rect 39842 6244 39852 6300
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 40116 6244 40126 6300
rect 43708 6244 43764 6300
rect 15810 6188 15820 6244
rect 15876 6188 17500 6244
rect 17556 6188 17566 6244
rect 21868 6188 25004 6244
rect 25060 6188 25070 6244
rect 25340 6188 28476 6244
rect 28532 6188 28542 6244
rect 29484 6188 31276 6244
rect 31332 6188 31342 6244
rect 41122 6188 41132 6244
rect 41188 6188 42196 6244
rect 5954 6076 5964 6132
rect 6020 6076 6188 6132
rect 6244 6076 15148 6132
rect 16706 6076 16716 6132
rect 16772 6076 19180 6132
rect 19236 6076 19246 6132
rect 23090 6076 23100 6132
rect 23156 6076 24332 6132
rect 24388 6076 24398 6132
rect 25218 6076 25228 6132
rect 25284 6076 28028 6132
rect 28084 6076 28094 6132
rect 29484 6020 29540 6188
rect 42140 6132 42196 6188
rect 42476 6188 43764 6244
rect 43922 6188 43932 6244
rect 43988 6188 44380 6244
rect 44436 6188 44446 6244
rect 42476 6132 42532 6188
rect 46732 6132 46788 6300
rect 59162 6244 59172 6300
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59436 6244 59446 6300
rect 47506 6188 47516 6244
rect 47572 6188 47964 6244
rect 48020 6188 48030 6244
rect 50978 6188 50988 6244
rect 51044 6188 51884 6244
rect 51940 6188 51950 6244
rect 59714 6188 59724 6244
rect 59780 6188 60956 6244
rect 61012 6188 61022 6244
rect 62524 6132 62580 6300
rect 64642 6188 64652 6244
rect 64708 6188 66108 6244
rect 66164 6188 66174 6244
rect 68562 6188 68572 6244
rect 68628 6188 72660 6244
rect 29698 6076 29708 6132
rect 29764 6076 33460 6132
rect 33404 6020 33460 6076
rect 35252 6076 40236 6132
rect 40292 6076 40302 6132
rect 42140 6076 42252 6132
rect 42308 6076 42318 6132
rect 42466 6076 42476 6132
rect 42532 6076 42542 6132
rect 43810 6076 43820 6132
rect 43876 6076 44604 6132
rect 44660 6076 44670 6132
rect 44818 6076 44828 6132
rect 44884 6076 46396 6132
rect 46452 6076 46462 6132
rect 46722 6076 46732 6132
rect 46788 6076 46798 6132
rect 47170 6076 47180 6132
rect 47236 6076 51100 6132
rect 51156 6076 51166 6132
rect 58594 6076 58604 6132
rect 58660 6076 62076 6132
rect 62132 6076 62142 6132
rect 62514 6076 62524 6132
rect 62580 6076 62590 6132
rect 63308 6076 69580 6132
rect 69636 6076 69646 6132
rect 70466 6076 70476 6132
rect 70532 6076 71036 6132
rect 71092 6076 71102 6132
rect 35252 6020 35308 6076
rect 40236 6020 40292 6076
rect 44828 6020 44884 6076
rect 8866 5964 8876 6020
rect 8932 5964 10332 6020
rect 10388 5964 13916 6020
rect 13972 5964 15708 6020
rect 15764 5964 15774 6020
rect 23874 5964 23884 6020
rect 23940 5964 27804 6020
rect 27860 5964 29540 6020
rect 31042 5964 31052 6020
rect 31108 5964 33180 6020
rect 33236 5964 33246 6020
rect 33404 5964 35308 6020
rect 39442 5964 39452 6020
rect 39508 5964 39788 6020
rect 39844 5964 39854 6020
rect 40236 5964 44380 6020
rect 44436 5964 44884 6020
rect 44940 5964 47628 6020
rect 47684 5964 47694 6020
rect 48290 5964 48300 6020
rect 48356 5964 57260 6020
rect 57316 5964 57326 6020
rect 58258 5964 58268 6020
rect 58324 5964 58828 6020
rect 58884 5964 58894 6020
rect 59052 5964 60172 6020
rect 60228 5964 60238 6020
rect 60386 5964 60396 6020
rect 60452 5964 62860 6020
rect 62916 5964 62926 6020
rect 44940 5908 44996 5964
rect 59052 5908 59108 5964
rect 8978 5852 8988 5908
rect 9044 5852 16044 5908
rect 16100 5852 16110 5908
rect 17378 5852 17388 5908
rect 17444 5852 17454 5908
rect 20738 5852 20748 5908
rect 20804 5852 22764 5908
rect 22820 5852 22830 5908
rect 24658 5852 24668 5908
rect 24724 5852 29932 5908
rect 29988 5852 29998 5908
rect 38434 5852 38444 5908
rect 38500 5852 39340 5908
rect 39396 5852 44940 5908
rect 44996 5852 45006 5908
rect 45276 5852 46508 5908
rect 46564 5852 46574 5908
rect 46722 5852 46732 5908
rect 46788 5852 48860 5908
rect 48916 5852 48926 5908
rect 49186 5852 49196 5908
rect 49252 5852 53228 5908
rect 53284 5852 53294 5908
rect 58482 5852 58492 5908
rect 58548 5852 59108 5908
rect 59490 5852 59500 5908
rect 59556 5852 60788 5908
rect 60946 5852 60956 5908
rect 61012 5852 63084 5908
rect 63140 5852 63150 5908
rect 17388 5796 17444 5852
rect 12674 5740 12684 5796
rect 12740 5740 13916 5796
rect 13972 5740 17444 5796
rect 23650 5740 23660 5796
rect 23716 5740 24108 5796
rect 24164 5740 24174 5796
rect 26786 5740 26796 5796
rect 26852 5740 30604 5796
rect 30660 5740 30670 5796
rect 42242 5740 42252 5796
rect 42308 5740 44828 5796
rect 44884 5740 44894 5796
rect 45276 5684 45332 5852
rect 60732 5796 60788 5852
rect 63308 5796 63364 6076
rect 72604 6020 72660 6188
rect 73500 6132 73556 6300
rect 78482 6244 78492 6300
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78756 6244 78766 6300
rect 73266 6076 73276 6132
rect 73332 6076 73556 6132
rect 73892 6188 75460 6244
rect 73892 6020 73948 6188
rect 64642 5964 64652 6020
rect 64708 5964 67788 6020
rect 67844 5964 67854 6020
rect 68002 5964 68012 6020
rect 68068 5964 68348 6020
rect 68404 5964 68414 6020
rect 70130 5964 70140 6020
rect 70196 5964 72380 6020
rect 72436 5964 72446 6020
rect 72604 5964 73948 6020
rect 75404 5908 75460 6188
rect 75618 5964 75628 6020
rect 75684 5964 77868 6020
rect 77924 5964 77934 6020
rect 63746 5852 63756 5908
rect 63812 5852 70812 5908
rect 70868 5852 70878 5908
rect 72818 5852 72828 5908
rect 72884 5852 73612 5908
rect 73668 5852 73678 5908
rect 75404 5852 76748 5908
rect 76804 5852 77644 5908
rect 77700 5852 77710 5908
rect 5058 5628 5068 5684
rect 5124 5628 6860 5684
rect 6916 5628 6926 5684
rect 7074 5628 7084 5684
rect 7140 5628 8764 5684
rect 8820 5628 8830 5684
rect 8978 5628 8988 5684
rect 9044 5628 9772 5684
rect 9828 5628 10556 5684
rect 10612 5628 10622 5684
rect 16146 5628 16156 5684
rect 16212 5628 17724 5684
rect 17780 5628 17790 5684
rect 24210 5628 24220 5684
rect 24276 5628 24668 5684
rect 24724 5628 24734 5684
rect 25106 5628 25116 5684
rect 25172 5628 32788 5684
rect 42130 5628 42140 5684
rect 42196 5628 43148 5684
rect 43204 5628 43596 5684
rect 43652 5628 43662 5684
rect 44370 5628 44380 5684
rect 44436 5628 45332 5684
rect 45500 5740 45836 5796
rect 45892 5740 51884 5796
rect 51940 5740 51950 5796
rect 54226 5740 54236 5796
rect 54292 5740 54684 5796
rect 54740 5740 54750 5796
rect 55234 5740 55244 5796
rect 55300 5740 55916 5796
rect 55972 5740 55982 5796
rect 56354 5740 56364 5796
rect 56420 5740 60396 5796
rect 60452 5740 60462 5796
rect 60732 5740 63364 5796
rect 69682 5740 69692 5796
rect 69748 5740 73948 5796
rect 3826 5516 3836 5572
rect 3892 5516 9324 5572
rect 9380 5516 9390 5572
rect 17602 5516 17612 5572
rect 17668 5516 23548 5572
rect 23604 5516 25060 5572
rect 26562 5516 26572 5572
rect 26628 5516 27580 5572
rect 27636 5516 27646 5572
rect 10862 5460 10872 5516
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 11136 5460 11146 5516
rect 4722 5404 4732 5460
rect 4788 5404 7756 5460
rect 7812 5404 7822 5460
rect 17154 5404 17164 5460
rect 17220 5404 21084 5460
rect 21140 5404 21150 5460
rect 5618 5292 5628 5348
rect 5684 5292 7084 5348
rect 7140 5292 7150 5348
rect 10882 5292 10892 5348
rect 10948 5292 13692 5348
rect 13748 5292 13758 5348
rect 15698 5292 15708 5348
rect 15764 5292 21308 5348
rect 21364 5292 21374 5348
rect 22754 5292 22764 5348
rect 22820 5292 24780 5348
rect 24836 5292 24846 5348
rect 25004 5236 25060 5516
rect 30182 5460 30192 5516
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30456 5460 30466 5516
rect 25330 5404 25340 5460
rect 25396 5404 28364 5460
rect 28420 5404 28430 5460
rect 27020 5292 27804 5348
rect 27860 5292 27870 5348
rect 27020 5236 27076 5292
rect 5842 5180 5852 5236
rect 5908 5180 6188 5236
rect 6244 5180 9548 5236
rect 9604 5180 9614 5236
rect 16594 5180 16604 5236
rect 16660 5180 21644 5236
rect 21700 5180 21710 5236
rect 22418 5180 22428 5236
rect 22484 5180 24612 5236
rect 25004 5180 25956 5236
rect 26674 5180 26684 5236
rect 26740 5180 27076 5236
rect 27234 5180 27244 5236
rect 27300 5180 29260 5236
rect 29316 5180 29326 5236
rect 29484 5180 30492 5236
rect 30548 5180 30558 5236
rect 24556 5124 24612 5180
rect 25900 5124 25956 5180
rect 29484 5124 29540 5180
rect 32732 5124 32788 5628
rect 45500 5572 45556 5740
rect 73892 5684 73948 5740
rect 37650 5516 37660 5572
rect 37716 5516 45556 5572
rect 45612 5628 46844 5684
rect 46900 5628 48972 5684
rect 49028 5628 49038 5684
rect 49746 5628 49756 5684
rect 49812 5628 49924 5684
rect 50866 5628 50876 5684
rect 50932 5628 53452 5684
rect 53508 5628 53518 5684
rect 58370 5628 58380 5684
rect 58436 5628 58446 5684
rect 58930 5628 58940 5684
rect 58996 5628 59500 5684
rect 59556 5628 59566 5684
rect 60050 5628 60060 5684
rect 60116 5628 60732 5684
rect 60788 5628 60798 5684
rect 61730 5628 61740 5684
rect 61796 5628 70476 5684
rect 70532 5628 70542 5684
rect 70802 5628 70812 5684
rect 70868 5628 72828 5684
rect 72884 5628 72894 5684
rect 73892 5628 75180 5684
rect 75236 5628 75246 5684
rect 45612 5460 45668 5628
rect 49868 5572 49924 5628
rect 58380 5572 58436 5628
rect 46050 5516 46060 5572
rect 46116 5516 49196 5572
rect 49252 5516 49262 5572
rect 49868 5516 50204 5572
rect 50260 5516 50270 5572
rect 51650 5516 51660 5572
rect 51716 5516 51996 5572
rect 52052 5516 52062 5572
rect 52770 5516 52780 5572
rect 52836 5516 54348 5572
rect 54404 5516 54414 5572
rect 55906 5516 55916 5572
rect 55972 5516 57708 5572
rect 57764 5516 57774 5572
rect 58380 5516 61516 5572
rect 61572 5516 61582 5572
rect 70914 5516 70924 5572
rect 70980 5516 74732 5572
rect 74788 5516 74798 5572
rect 49502 5460 49512 5516
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49776 5460 49786 5516
rect 68822 5460 68832 5516
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 69096 5460 69106 5516
rect 42914 5404 42924 5460
rect 42980 5404 45276 5460
rect 45332 5404 45342 5460
rect 45602 5404 45612 5460
rect 45668 5404 45678 5460
rect 46274 5404 46284 5460
rect 46340 5404 46732 5460
rect 46788 5404 46798 5460
rect 51996 5404 56028 5460
rect 56084 5404 59948 5460
rect 60004 5404 60284 5460
rect 60340 5404 60350 5460
rect 60610 5404 60620 5460
rect 60676 5404 62076 5460
rect 62132 5404 62142 5460
rect 64194 5404 64204 5460
rect 64260 5404 67228 5460
rect 67284 5404 67294 5460
rect 71698 5404 71708 5460
rect 71764 5404 77196 5460
rect 77252 5404 77262 5460
rect 51996 5348 52052 5404
rect 37874 5292 37884 5348
rect 37940 5292 43988 5348
rect 43932 5236 43988 5292
rect 46172 5292 49644 5348
rect 49700 5292 50316 5348
rect 50372 5292 50382 5348
rect 51986 5292 51996 5348
rect 52052 5292 52062 5348
rect 52210 5292 52220 5348
rect 52276 5292 52780 5348
rect 52836 5292 52846 5348
rect 55682 5292 55692 5348
rect 55748 5292 61684 5348
rect 62626 5292 62636 5348
rect 62692 5292 63980 5348
rect 64036 5292 77532 5348
rect 77588 5292 77598 5348
rect 35970 5180 35980 5236
rect 36036 5180 37212 5236
rect 37268 5180 37278 5236
rect 41346 5180 41356 5236
rect 41412 5180 43708 5236
rect 43764 5180 43774 5236
rect 43932 5180 44996 5236
rect 44940 5124 44996 5180
rect 2594 5068 2604 5124
rect 2660 5068 6412 5124
rect 6468 5068 6478 5124
rect 9874 5068 9884 5124
rect 9940 5068 13692 5124
rect 13748 5068 13758 5124
rect 16034 5068 16044 5124
rect 16100 5068 16940 5124
rect 16996 5068 17006 5124
rect 18050 5068 18060 5124
rect 18116 5068 19964 5124
rect 20020 5068 20860 5124
rect 20916 5068 20926 5124
rect 22306 5068 22316 5124
rect 22372 5068 23436 5124
rect 23492 5068 24332 5124
rect 24388 5068 24398 5124
rect 24556 5068 25844 5124
rect 25900 5068 29540 5124
rect 29810 5068 29820 5124
rect 29876 5068 30604 5124
rect 30660 5068 30670 5124
rect 32732 5068 44884 5124
rect 44940 5068 45668 5124
rect 5730 4956 5740 5012
rect 5796 4956 7420 5012
rect 7476 4956 7486 5012
rect 16146 4956 16156 5012
rect 16212 4956 18508 5012
rect 18564 4956 18574 5012
rect 22194 4956 22204 5012
rect 22260 4956 23324 5012
rect 23380 4956 23390 5012
rect 25788 4900 25844 5068
rect 44828 5012 44884 5068
rect 45612 5012 45668 5068
rect 26002 4956 26012 5012
rect 26068 4956 28140 5012
rect 28196 4956 28206 5012
rect 42018 4956 42028 5012
rect 42084 4956 43988 5012
rect 44818 4956 44828 5012
rect 44884 4956 44894 5012
rect 45602 4956 45612 5012
rect 45668 4956 45678 5012
rect 43932 4900 43988 4956
rect 46172 4900 46228 5292
rect 46610 5180 46620 5236
rect 46676 5180 46844 5236
rect 46900 5180 46910 5236
rect 48962 5180 48972 5236
rect 49028 5180 51772 5236
rect 51828 5180 51838 5236
rect 53442 5180 53452 5236
rect 53508 5180 53518 5236
rect 54674 5180 54684 5236
rect 54740 5180 58716 5236
rect 58772 5180 58782 5236
rect 59500 5180 60620 5236
rect 60676 5180 61404 5236
rect 61460 5180 61470 5236
rect 53452 5124 53508 5180
rect 59500 5124 59556 5180
rect 61628 5124 61684 5292
rect 64082 5180 64092 5236
rect 64148 5180 64764 5236
rect 64820 5180 65100 5236
rect 65156 5180 65166 5236
rect 69570 5180 69580 5236
rect 69636 5180 70588 5236
rect 70644 5180 70654 5236
rect 72370 5180 72380 5236
rect 72436 5180 76300 5236
rect 76356 5180 76366 5236
rect 48178 5068 48188 5124
rect 48244 5068 52220 5124
rect 52276 5068 52286 5124
rect 52556 5068 53508 5124
rect 56130 5068 56140 5124
rect 56196 5068 59556 5124
rect 61058 5068 61068 5124
rect 61124 5068 61684 5124
rect 66770 5068 66780 5124
rect 66836 5068 70364 5124
rect 70420 5068 70430 5124
rect 73266 5068 73276 5124
rect 73332 5068 75964 5124
rect 76020 5068 76030 5124
rect 49746 4956 49756 5012
rect 49812 4956 49822 5012
rect 3378 4844 3388 4900
rect 3444 4844 4620 4900
rect 4676 4844 6524 4900
rect 6580 4844 6590 4900
rect 8754 4844 8764 4900
rect 8820 4844 19852 4900
rect 19908 4844 19918 4900
rect 22866 4844 22876 4900
rect 22932 4844 23772 4900
rect 23828 4844 23838 4900
rect 25788 4844 26348 4900
rect 26404 4844 26414 4900
rect 26786 4844 26796 4900
rect 26852 4844 30716 4900
rect 30772 4844 30782 4900
rect 30930 4844 30940 4900
rect 30996 4844 31948 4900
rect 32004 4844 32014 4900
rect 42466 4844 42476 4900
rect 42532 4844 43708 4900
rect 43764 4844 43774 4900
rect 43922 4844 43932 4900
rect 43988 4844 43998 4900
rect 44258 4844 44268 4900
rect 44324 4844 45388 4900
rect 45444 4844 45454 4900
rect 45724 4844 46228 4900
rect 26348 4788 26404 4844
rect 45724 4788 45780 4844
rect 49756 4788 49812 4956
rect 52556 4900 52612 5068
rect 53106 4956 53116 5012
rect 53172 4956 55468 5012
rect 55524 4956 55534 5012
rect 65874 4956 65884 5012
rect 65940 4956 67788 5012
rect 67844 4956 67854 5012
rect 68114 4956 68124 5012
rect 68180 4956 68460 5012
rect 68516 4956 68526 5012
rect 69010 4956 69020 5012
rect 69076 4956 69468 5012
rect 69524 4956 69534 5012
rect 70466 4956 70476 5012
rect 70532 4956 72044 5012
rect 72100 4956 72110 5012
rect 72818 4956 72828 5012
rect 72884 4956 74396 5012
rect 74452 4956 74462 5012
rect 50306 4844 50316 4900
rect 50372 4844 52612 4900
rect 54786 4844 54796 4900
rect 54852 4844 56924 4900
rect 56980 4844 56990 4900
rect 57698 4844 57708 4900
rect 57764 4844 58716 4900
rect 58772 4844 59388 4900
rect 59444 4844 59454 4900
rect 67890 4844 67900 4900
rect 67956 4844 69244 4900
rect 69300 4844 69310 4900
rect 69794 4844 69804 4900
rect 69860 4844 70364 4900
rect 70420 4844 70430 4900
rect 21074 4732 21084 4788
rect 21140 4732 24108 4788
rect 24164 4732 24174 4788
rect 24882 4732 24892 4788
rect 24948 4732 25788 4788
rect 25844 4732 25854 4788
rect 26348 4732 30660 4788
rect 42476 4732 44156 4788
rect 44212 4732 44222 4788
rect 44828 4732 45780 4788
rect 45938 4732 45948 4788
rect 46004 4732 49812 4788
rect 52434 4732 52444 4788
rect 52500 4732 54012 4788
rect 54068 4732 54078 4788
rect 54898 4732 54908 4788
rect 54964 4732 55356 4788
rect 55412 4732 55422 4788
rect 56242 4732 56252 4788
rect 56308 4732 57932 4788
rect 57988 4732 57998 4788
rect 59938 4732 59948 4788
rect 60004 4732 62300 4788
rect 62356 4732 62366 4788
rect 63746 4732 63756 4788
rect 63812 4732 66668 4788
rect 66724 4732 66734 4788
rect 67778 4732 67788 4788
rect 67844 4732 68348 4788
rect 68404 4732 68414 4788
rect 20522 4676 20532 4732
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20796 4676 20806 4732
rect 30604 4676 30660 4732
rect 39842 4676 39852 4732
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 40116 4676 40126 4732
rect 42476 4676 42532 4732
rect 44828 4676 44884 4732
rect 59162 4676 59172 4732
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59436 4676 59446 4732
rect 78482 4676 78492 4732
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78756 4676 78766 4732
rect 26898 4620 26908 4676
rect 26964 4620 29148 4676
rect 29204 4620 29214 4676
rect 30604 4620 33628 4676
rect 42466 4620 42476 4676
rect 42532 4620 42542 4676
rect 42802 4620 42812 4676
rect 42868 4620 43596 4676
rect 43652 4620 43662 4676
rect 43810 4620 43820 4676
rect 43876 4620 43886 4676
rect 44156 4620 44828 4676
rect 44884 4620 44894 4676
rect 45266 4620 45276 4676
rect 45332 4620 46620 4676
rect 46676 4620 46686 4676
rect 47730 4620 47740 4676
rect 47796 4620 48188 4676
rect 48244 4620 48254 4676
rect 51090 4620 51100 4676
rect 51156 4620 52332 4676
rect 52388 4620 52398 4676
rect 52658 4620 52668 4676
rect 52724 4620 55468 4676
rect 55524 4620 55534 4676
rect 59714 4620 59724 4676
rect 59780 4620 63532 4676
rect 63588 4620 63598 4676
rect 63970 4620 63980 4676
rect 64036 4620 64540 4676
rect 64596 4620 64606 4676
rect 67330 4620 67340 4676
rect 67396 4620 68124 4676
rect 68180 4620 68190 4676
rect 72482 4620 72492 4676
rect 72548 4620 74284 4676
rect 74340 4620 74350 4676
rect 33572 4564 33628 4620
rect 43820 4564 43876 4620
rect 7298 4508 7308 4564
rect 7364 4508 10668 4564
rect 10724 4508 13412 4564
rect 18386 4508 18396 4564
rect 18452 4508 20748 4564
rect 20804 4508 20814 4564
rect 23314 4508 23324 4564
rect 23380 4508 24220 4564
rect 24276 4508 24286 4564
rect 27682 4508 27692 4564
rect 27748 4508 31164 4564
rect 31220 4508 31230 4564
rect 33572 4508 33964 4564
rect 34020 4508 36652 4564
rect 36708 4508 43876 4564
rect 4274 4396 4284 4452
rect 4340 4396 13132 4452
rect 13188 4396 13198 4452
rect 13356 4340 13412 4508
rect 44156 4452 44212 4620
rect 45378 4508 45388 4564
rect 45444 4508 45948 4564
rect 46004 4508 46014 4564
rect 46834 4508 46844 4564
rect 46900 4508 46910 4564
rect 47954 4508 47964 4564
rect 48020 4508 53172 4564
rect 53330 4508 53340 4564
rect 53396 4508 54124 4564
rect 54180 4508 56140 4564
rect 56196 4508 56206 4564
rect 57922 4508 57932 4564
rect 57988 4508 63644 4564
rect 63700 4508 63710 4564
rect 64418 4508 64428 4564
rect 64484 4508 65548 4564
rect 65604 4508 67228 4564
rect 67284 4508 67294 4564
rect 67442 4508 67452 4564
rect 67508 4508 73836 4564
rect 73892 4508 76076 4564
rect 76132 4508 76142 4564
rect 46844 4452 46900 4508
rect 14914 4396 14924 4452
rect 14980 4396 22092 4452
rect 22148 4396 22158 4452
rect 25890 4396 25900 4452
rect 25956 4396 29036 4452
rect 29092 4396 29102 4452
rect 34514 4396 34524 4452
rect 34580 4396 39564 4452
rect 39620 4396 39630 4452
rect 40898 4396 40908 4452
rect 40964 4396 44212 4452
rect 44716 4396 46172 4452
rect 46228 4396 46238 4452
rect 46610 4396 46620 4452
rect 46676 4396 46900 4452
rect 53116 4452 53172 4508
rect 53116 4396 57484 4452
rect 57540 4396 57550 4452
rect 62402 4396 62412 4452
rect 62468 4396 63420 4452
rect 63476 4396 64540 4452
rect 64596 4396 64606 4452
rect 65762 4396 65772 4452
rect 65828 4396 66444 4452
rect 66500 4396 66510 4452
rect 67554 4396 67564 4452
rect 67620 4396 69468 4452
rect 69524 4396 69534 4452
rect 69794 4396 69804 4452
rect 69860 4396 70924 4452
rect 70980 4396 70990 4452
rect 71474 4396 71484 4452
rect 71540 4396 75180 4452
rect 75236 4396 75246 4452
rect 44716 4340 44772 4396
rect 2258 4284 2268 4340
rect 2324 4284 8316 4340
rect 8372 4284 8382 4340
rect 13356 4284 23100 4340
rect 23156 4284 23166 4340
rect 23874 4284 23884 4340
rect 23940 4284 26348 4340
rect 26404 4284 26414 4340
rect 27682 4284 27692 4340
rect 27748 4284 28700 4340
rect 28756 4284 28766 4340
rect 33618 4284 33628 4340
rect 33684 4284 37548 4340
rect 37604 4284 37614 4340
rect 40338 4284 40348 4340
rect 40404 4284 41916 4340
rect 41972 4284 41982 4340
rect 42476 4284 43708 4340
rect 43764 4284 44044 4340
rect 44100 4284 44110 4340
rect 44492 4284 44772 4340
rect 45332 4284 46844 4340
rect 46900 4284 46910 4340
rect 47170 4284 47180 4340
rect 47236 4284 52668 4340
rect 52724 4284 52734 4340
rect 52994 4284 53004 4340
rect 53060 4284 53900 4340
rect 53956 4284 54908 4340
rect 54964 4284 54974 4340
rect 68114 4284 68124 4340
rect 68180 4284 71596 4340
rect 71652 4284 73164 4340
rect 73220 4284 73230 4340
rect 42476 4228 42532 4284
rect 44492 4228 44548 4284
rect 45332 4228 45388 4284
rect 7858 4172 7868 4228
rect 7924 4172 8876 4228
rect 8932 4172 8942 4228
rect 24098 4172 24108 4228
rect 24164 4172 24668 4228
rect 24724 4172 25900 4228
rect 25956 4172 26124 4228
rect 26180 4172 26190 4228
rect 26674 4172 26684 4228
rect 26740 4172 29372 4228
rect 29428 4172 29438 4228
rect 41794 4172 41804 4228
rect 41860 4172 42532 4228
rect 42690 4172 42700 4228
rect 42756 4172 43820 4228
rect 43876 4172 44548 4228
rect 45052 4172 45388 4228
rect 49410 4172 49420 4228
rect 49476 4172 49486 4228
rect 52546 4172 52556 4228
rect 52612 4172 59388 4228
rect 59444 4172 61068 4228
rect 61124 4172 61134 4228
rect 62188 4172 62860 4228
rect 62916 4172 62926 4228
rect 63858 4172 63868 4228
rect 63924 4172 65772 4228
rect 65828 4172 65838 4228
rect 66882 4172 66892 4228
rect 66948 4172 67676 4228
rect 67732 4172 67742 4228
rect 4834 4060 4844 4116
rect 4900 4060 9884 4116
rect 9940 4060 9950 4116
rect 10668 4060 15148 4116
rect 23874 4060 23884 4116
rect 23940 4060 27356 4116
rect 27412 4060 27422 4116
rect 28588 4060 33068 4116
rect 33124 4060 33134 4116
rect 39890 4060 39900 4116
rect 39956 4060 41132 4116
rect 41188 4060 41198 4116
rect 41458 4060 41468 4116
rect 41524 4060 43036 4116
rect 43092 4060 43102 4116
rect 44370 4060 44380 4116
rect 44436 4060 44884 4116
rect 10668 4004 10724 4060
rect 3332 3948 5628 4004
rect 5684 3948 5694 4004
rect 9314 3948 9324 4004
rect 9380 3948 10724 4004
rect 3266 3836 3276 3892
rect 3332 3836 3388 3948
rect 10862 3892 10872 3948
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 11136 3892 11146 3948
rect 15092 3892 15148 4060
rect 24770 3948 24780 4004
rect 24836 3948 24846 4004
rect 26562 3948 26572 4004
rect 26628 3948 27580 4004
rect 27636 3948 27646 4004
rect 24780 3892 24836 3948
rect 28588 3892 28644 4060
rect 44828 4004 44884 4060
rect 45052 4004 45108 4172
rect 49420 4116 49476 4172
rect 62188 4116 62244 4172
rect 46162 4060 46172 4116
rect 46228 4060 49476 4116
rect 53330 4060 53340 4116
rect 53396 4060 53564 4116
rect 53620 4060 54236 4116
rect 54292 4060 54302 4116
rect 55010 4060 55020 4116
rect 55076 4060 55468 4116
rect 55524 4060 55534 4116
rect 59154 4060 59164 4116
rect 59220 4060 62244 4116
rect 62402 4060 62412 4116
rect 62468 4060 64652 4116
rect 64708 4060 64718 4116
rect 67218 4060 67228 4116
rect 67284 4060 68460 4116
rect 68516 4060 68526 4116
rect 68786 4060 68796 4116
rect 68852 4060 73612 4116
rect 73668 4060 74284 4116
rect 74340 4060 74350 4116
rect 33730 3948 33740 4004
rect 33796 3948 43708 4004
rect 43764 3948 43774 4004
rect 44828 3948 45108 4004
rect 45266 3948 45276 4004
rect 45332 3948 46732 4004
rect 46788 3948 46798 4004
rect 47058 3948 47068 4004
rect 47124 3948 47404 4004
rect 47460 3948 47470 4004
rect 52994 3948 53004 4004
rect 53060 3948 53676 4004
rect 53732 3948 60620 4004
rect 60676 3948 60686 4004
rect 61170 3948 61180 4004
rect 61236 3948 62076 4004
rect 62132 3948 62860 4004
rect 62916 3948 62926 4004
rect 30182 3892 30192 3948
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30456 3892 30466 3948
rect 49502 3892 49512 3948
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49776 3892 49786 3948
rect 68822 3892 68832 3948
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 69096 3892 69106 3948
rect 3490 3836 3500 3892
rect 3556 3836 9212 3892
rect 9268 3836 9278 3892
rect 15092 3836 17836 3892
rect 17892 3836 17902 3892
rect 24780 3836 28588 3892
rect 28644 3836 28654 3892
rect 38994 3836 39004 3892
rect 39060 3836 45388 3892
rect 45444 3836 45454 3892
rect 50530 3836 50540 3892
rect 50596 3836 51548 3892
rect 51604 3836 51614 3892
rect 55010 3836 55020 3892
rect 55076 3836 56924 3892
rect 56980 3836 56990 3892
rect 57250 3836 57260 3892
rect 57316 3836 65548 3892
rect 65604 3836 65614 3892
rect 2482 3724 2492 3780
rect 2548 3724 9772 3780
rect 9828 3724 9838 3780
rect 9996 3724 15484 3780
rect 15540 3724 15550 3780
rect 18162 3724 18172 3780
rect 18228 3724 23828 3780
rect 23986 3724 23996 3780
rect 24052 3724 26124 3780
rect 26180 3724 26190 3780
rect 32386 3724 32396 3780
rect 32452 3724 36988 3780
rect 37044 3724 37054 3780
rect 43138 3724 43148 3780
rect 43204 3724 44716 3780
rect 44772 3724 44782 3780
rect 44940 3724 47404 3780
rect 47460 3724 47470 3780
rect 56466 3724 56476 3780
rect 56532 3724 57148 3780
rect 57204 3724 57214 3780
rect 57810 3724 57820 3780
rect 57876 3724 59052 3780
rect 59108 3724 59118 3780
rect 61170 3724 61180 3780
rect 61236 3724 62748 3780
rect 62804 3724 62814 3780
rect 64530 3724 64540 3780
rect 64596 3724 65212 3780
rect 65268 3724 65278 3780
rect 65884 3724 71036 3780
rect 71092 3724 71102 3780
rect 71922 3724 71932 3780
rect 71988 3724 78092 3780
rect 78148 3724 78158 3780
rect 9996 3668 10052 3724
rect 23772 3668 23828 3724
rect 44940 3668 44996 3724
rect 65884 3668 65940 3724
rect 2930 3612 2940 3668
rect 2996 3612 3668 3668
rect 5618 3612 5628 3668
rect 5684 3612 10052 3668
rect 11554 3612 11564 3668
rect 11620 3612 16380 3668
rect 16436 3612 16446 3668
rect 17938 3612 17948 3668
rect 18004 3612 21868 3668
rect 21924 3612 21934 3668
rect 23772 3612 25116 3668
rect 25172 3612 25182 3668
rect 26450 3612 26460 3668
rect 26516 3612 27412 3668
rect 27570 3612 27580 3668
rect 27636 3612 28812 3668
rect 28868 3612 28878 3668
rect 34402 3612 34412 3668
rect 34468 3612 35644 3668
rect 35700 3612 35710 3668
rect 43362 3612 43372 3668
rect 43428 3612 44940 3668
rect 44996 3612 45006 3668
rect 45164 3612 46060 3668
rect 46116 3612 46126 3668
rect 46508 3612 47628 3668
rect 47684 3612 47694 3668
rect 52210 3612 52220 3668
rect 52276 3612 52556 3668
rect 52612 3612 53676 3668
rect 53732 3612 54572 3668
rect 54628 3612 55916 3668
rect 55972 3612 55982 3668
rect 57026 3612 57036 3668
rect 57092 3612 57596 3668
rect 57652 3612 57662 3668
rect 62290 3612 62300 3668
rect 62356 3612 65940 3668
rect 3612 3556 3668 3612
rect 27356 3556 27412 3612
rect 45164 3556 45220 3612
rect 2258 3500 2268 3556
rect 2324 3500 3388 3556
rect 3444 3500 3454 3556
rect 3602 3500 3612 3556
rect 3668 3500 6972 3556
rect 7028 3500 7038 3556
rect 13122 3500 13132 3556
rect 13188 3500 18172 3556
rect 18228 3500 18238 3556
rect 22530 3500 22540 3556
rect 22596 3500 24892 3556
rect 24948 3500 24958 3556
rect 25890 3500 25900 3556
rect 25956 3500 27132 3556
rect 27188 3500 27198 3556
rect 27356 3500 32284 3556
rect 32340 3500 33628 3556
rect 33684 3500 33694 3556
rect 44146 3500 44156 3556
rect 44212 3500 44492 3556
rect 44548 3500 45220 3556
rect 1922 3388 1932 3444
rect 1988 3388 4508 3444
rect 4564 3388 7196 3444
rect 7252 3388 7262 3444
rect 7746 3388 7756 3444
rect 7812 3388 14364 3444
rect 14420 3388 14430 3444
rect 14802 3388 14812 3444
rect 14868 3388 18396 3444
rect 18452 3388 18462 3444
rect 24658 3388 24668 3444
rect 24724 3388 29820 3444
rect 29876 3388 29886 3444
rect 33170 3388 33180 3444
rect 33236 3388 41020 3444
rect 41076 3388 41086 3444
rect 42466 3388 42476 3444
rect 42532 3388 43148 3444
rect 43204 3388 43214 3444
rect 44818 3388 44828 3444
rect 44884 3388 46284 3444
rect 46340 3388 46350 3444
rect 46508 3332 46564 3612
rect 48738 3500 48748 3556
rect 48804 3500 50428 3556
rect 50484 3500 50494 3556
rect 59714 3500 59724 3556
rect 59780 3500 60172 3556
rect 60228 3500 60238 3556
rect 64866 3500 64876 3556
rect 64932 3500 66892 3556
rect 66948 3500 66958 3556
rect 69010 3500 69020 3556
rect 69076 3500 74956 3556
rect 75012 3500 75022 3556
rect 46946 3388 46956 3444
rect 47012 3388 48076 3444
rect 48132 3388 48142 3444
rect 53666 3388 53676 3444
rect 53732 3388 55356 3444
rect 55412 3388 55422 3444
rect 58706 3388 58716 3444
rect 58772 3388 59668 3444
rect 13458 3276 13468 3332
rect 13524 3276 13804 3332
rect 13860 3276 13870 3332
rect 26674 3276 26684 3332
rect 26740 3276 28252 3332
rect 28308 3276 28318 3332
rect 35298 3276 35308 3332
rect 35364 3276 36316 3332
rect 36372 3276 36382 3332
rect 39218 3276 39228 3332
rect 39284 3276 44044 3332
rect 44100 3276 45052 3332
rect 45108 3276 45118 3332
rect 45490 3276 45500 3332
rect 45556 3276 45836 3332
rect 45892 3276 45902 3332
rect 46162 3276 46172 3332
rect 46228 3276 46564 3332
rect 46722 3276 46732 3332
rect 46788 3276 50204 3332
rect 50260 3276 50270 3332
rect 51538 3276 51548 3332
rect 51604 3276 58940 3332
rect 58996 3276 59006 3332
rect 27906 3164 27916 3220
rect 27972 3164 29148 3220
rect 29204 3164 29214 3220
rect 42130 3164 42140 3220
rect 42196 3164 44940 3220
rect 44996 3164 45006 3220
rect 45500 3164 57484 3220
rect 57540 3164 57550 3220
rect 20522 3108 20532 3164
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20796 3108 20806 3164
rect 39842 3108 39852 3164
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 40116 3108 40126 3164
rect 45500 3108 45556 3164
rect 59162 3108 59172 3164
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59436 3108 59446 3164
rect 59612 3108 59668 3388
rect 60956 3388 62524 3444
rect 62580 3388 62590 3444
rect 65436 3388 67452 3444
rect 67508 3388 67518 3444
rect 69020 3388 69524 3444
rect 72146 3388 72156 3444
rect 72212 3388 78092 3444
rect 78148 3388 78158 3444
rect 60956 3332 61012 3388
rect 65436 3332 65492 3388
rect 69020 3332 69076 3388
rect 60946 3276 60956 3332
rect 61012 3276 61022 3332
rect 61842 3276 61852 3332
rect 61908 3276 62188 3332
rect 62244 3276 62254 3332
rect 65426 3276 65436 3332
rect 65492 3276 65502 3332
rect 65650 3276 65660 3332
rect 65716 3276 69076 3332
rect 69468 3332 69524 3388
rect 69468 3276 72044 3332
rect 72100 3276 72110 3332
rect 59826 3164 59836 3220
rect 59892 3164 60732 3220
rect 60788 3164 60798 3220
rect 62626 3164 62636 3220
rect 62692 3164 75628 3220
rect 75684 3164 75694 3220
rect 78482 3108 78492 3164
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78756 3108 78766 3164
rect 41906 3052 41916 3108
rect 41972 3052 45276 3108
rect 45332 3052 45342 3108
rect 45490 3052 45500 3108
rect 45556 3052 45566 3108
rect 46610 3052 46620 3108
rect 46676 3052 56812 3108
rect 56868 3052 56878 3108
rect 59612 3052 69132 3108
rect 69188 3052 69198 3108
rect 9650 2940 9660 2996
rect 9716 2940 42700 2996
rect 42756 2940 42766 2996
rect 44706 2940 44716 2996
rect 44772 2940 52108 2996
rect 52164 2940 52174 2996
rect 59602 2940 59612 2996
rect 59668 2940 60396 2996
rect 60452 2940 60462 2996
rect 61730 2940 61740 2996
rect 61796 2940 77980 2996
rect 78036 2940 78046 2996
rect 16034 2828 16044 2884
rect 16100 2828 38556 2884
rect 38612 2828 38622 2884
rect 42354 2828 42364 2884
rect 42420 2828 50316 2884
rect 50372 2828 50382 2884
rect 60050 2828 60060 2884
rect 60116 2828 73164 2884
rect 73220 2828 73230 2884
rect 18610 2716 18620 2772
rect 18676 2716 50764 2772
rect 50820 2716 50830 2772
rect 55682 2716 55692 2772
rect 55748 2716 56700 2772
rect 56756 2716 64204 2772
rect 64260 2716 64270 2772
rect 4050 2604 4060 2660
rect 4116 2604 53340 2660
rect 53396 2604 53406 2660
rect 2930 2492 2940 2548
rect 2996 2492 12796 2548
rect 12852 2492 12862 2548
rect 25666 2492 25676 2548
rect 25732 2492 35308 2548
rect 35364 2492 35374 2548
rect 45042 2492 45052 2548
rect 45108 2492 58044 2548
rect 58100 2492 58110 2548
rect 65650 2492 65660 2548
rect 65716 2492 71820 2548
rect 71876 2492 71886 2548
rect 3154 2380 3164 2436
rect 3220 2380 31052 2436
rect 31108 2380 31118 2436
rect 39554 2380 39564 2436
rect 39620 2380 51884 2436
rect 51940 2380 51950 2436
rect 26338 2268 26348 2324
rect 26404 2268 57372 2324
rect 57428 2268 57438 2324
rect 50372 1820 51436 1876
rect 51492 1820 51502 1876
rect 50372 1764 50428 1820
rect 50194 1708 50204 1764
rect 50260 1708 50428 1764
rect 50764 1708 51716 1764
rect 55794 1708 55804 1764
rect 55860 1708 61964 1764
rect 62020 1708 62030 1764
rect 50764 1652 50820 1708
rect 20636 1596 33124 1652
rect 13794 1372 13804 1428
rect 13860 1372 20300 1428
rect 20356 1372 20366 1428
rect 20636 1316 20692 1596
rect 33068 1540 33124 1596
rect 38612 1596 43372 1652
rect 43428 1596 43438 1652
rect 44258 1596 44268 1652
rect 44324 1596 50820 1652
rect 51660 1652 51716 1708
rect 51660 1596 56140 1652
rect 56196 1596 56206 1652
rect 8372 1260 20692 1316
rect 20860 1484 32732 1540
rect 32788 1484 32798 1540
rect 33058 1484 33068 1540
rect 33124 1484 33134 1540
rect 8372 1092 8428 1260
rect 20860 1204 20916 1484
rect 38612 1428 38668 1596
rect 38770 1484 38780 1540
rect 38836 1484 49308 1540
rect 49364 1484 49374 1540
rect 50652 1484 63084 1540
rect 63140 1484 63150 1540
rect 50652 1428 50708 1484
rect 10098 1148 10108 1204
rect 10164 1148 20916 1204
rect 21196 1372 38668 1428
rect 46834 1372 46844 1428
rect 46900 1372 50708 1428
rect 21196 1092 21252 1372
rect 24882 1260 24892 1316
rect 24948 1260 42252 1316
rect 42308 1260 42318 1316
rect 43810 1260 43820 1316
rect 43876 1260 56028 1316
rect 56084 1260 56094 1316
rect 42018 1148 42028 1204
rect 42084 1148 59052 1204
rect 59108 1148 59118 1204
rect 5842 1036 5852 1092
rect 5908 1036 8428 1092
rect 16930 1036 16940 1092
rect 16996 1036 17006 1092
rect 20290 1036 20300 1092
rect 20356 1036 21252 1092
rect 23492 1036 32564 1092
rect 33058 1036 33068 1092
rect 33124 1036 50204 1092
rect 50260 1036 50270 1092
rect 16940 84 16996 1036
rect 18946 924 18956 980
rect 19012 924 19022 980
rect 18956 644 19012 924
rect 23492 644 23548 1036
rect 18956 588 23548 644
rect 24556 924 27132 980
rect 27188 924 27198 980
rect 28018 924 28028 980
rect 28084 924 28094 980
rect 24556 84 24612 924
rect 28028 420 28084 924
rect 32508 868 32564 1036
rect 32722 924 32732 980
rect 32788 924 40908 980
rect 40964 924 40974 980
rect 43138 924 43148 980
rect 43204 924 43214 980
rect 45332 924 45612 980
rect 45668 924 45678 980
rect 45826 924 45836 980
rect 45892 924 55692 980
rect 55748 924 55758 980
rect 43148 868 43204 924
rect 32508 812 43204 868
rect 45332 420 45388 924
rect 28028 364 45388 420
rect 16940 28 24612 84
<< via3 >>
rect 10872 36820 10928 36876
rect 10976 36820 11032 36876
rect 11080 36820 11136 36876
rect 30192 36820 30248 36876
rect 30296 36820 30352 36876
rect 30400 36820 30456 36876
rect 49512 36820 49568 36876
rect 49616 36820 49672 36876
rect 49720 36820 49776 36876
rect 68832 36820 68888 36876
rect 68936 36820 68992 36876
rect 69040 36820 69096 36876
rect 20532 36036 20588 36092
rect 20636 36036 20692 36092
rect 20740 36036 20796 36092
rect 39852 36036 39908 36092
rect 39956 36036 40012 36092
rect 40060 36036 40116 36092
rect 59172 36036 59228 36092
rect 59276 36036 59332 36092
rect 59380 36036 59436 36092
rect 78492 36036 78548 36092
rect 78596 36036 78652 36092
rect 78700 36036 78756 36092
rect 10872 35252 10928 35308
rect 10976 35252 11032 35308
rect 11080 35252 11136 35308
rect 30192 35252 30248 35308
rect 30296 35252 30352 35308
rect 30400 35252 30456 35308
rect 49512 35252 49568 35308
rect 49616 35252 49672 35308
rect 49720 35252 49776 35308
rect 68832 35252 68888 35308
rect 68936 35252 68992 35308
rect 69040 35252 69096 35308
rect 20532 34468 20588 34524
rect 20636 34468 20692 34524
rect 20740 34468 20796 34524
rect 39852 34468 39908 34524
rect 39956 34468 40012 34524
rect 40060 34468 40116 34524
rect 59172 34468 59228 34524
rect 59276 34468 59332 34524
rect 59380 34468 59436 34524
rect 78492 34468 78548 34524
rect 78596 34468 78652 34524
rect 78700 34468 78756 34524
rect 10872 33684 10928 33740
rect 10976 33684 11032 33740
rect 11080 33684 11136 33740
rect 30192 33684 30248 33740
rect 30296 33684 30352 33740
rect 30400 33684 30456 33740
rect 49512 33684 49568 33740
rect 49616 33684 49672 33740
rect 49720 33684 49776 33740
rect 68832 33684 68888 33740
rect 68936 33684 68992 33740
rect 69040 33684 69096 33740
rect 20532 32900 20588 32956
rect 20636 32900 20692 32956
rect 20740 32900 20796 32956
rect 39852 32900 39908 32956
rect 39956 32900 40012 32956
rect 40060 32900 40116 32956
rect 59172 32900 59228 32956
rect 59276 32900 59332 32956
rect 59380 32900 59436 32956
rect 78492 32900 78548 32956
rect 78596 32900 78652 32956
rect 78700 32900 78756 32956
rect 10872 32116 10928 32172
rect 10976 32116 11032 32172
rect 11080 32116 11136 32172
rect 30192 32116 30248 32172
rect 30296 32116 30352 32172
rect 30400 32116 30456 32172
rect 49512 32116 49568 32172
rect 49616 32116 49672 32172
rect 49720 32116 49776 32172
rect 68832 32116 68888 32172
rect 68936 32116 68992 32172
rect 69040 32116 69096 32172
rect 20532 31332 20588 31388
rect 20636 31332 20692 31388
rect 20740 31332 20796 31388
rect 39852 31332 39908 31388
rect 39956 31332 40012 31388
rect 40060 31332 40116 31388
rect 59172 31332 59228 31388
rect 59276 31332 59332 31388
rect 59380 31332 59436 31388
rect 78492 31332 78548 31388
rect 78596 31332 78652 31388
rect 78700 31332 78756 31388
rect 10872 30548 10928 30604
rect 10976 30548 11032 30604
rect 11080 30548 11136 30604
rect 30192 30548 30248 30604
rect 30296 30548 30352 30604
rect 30400 30548 30456 30604
rect 49512 30548 49568 30604
rect 49616 30548 49672 30604
rect 49720 30548 49776 30604
rect 68832 30548 68888 30604
rect 68936 30548 68992 30604
rect 69040 30548 69096 30604
rect 20532 29764 20588 29820
rect 20636 29764 20692 29820
rect 20740 29764 20796 29820
rect 39852 29764 39908 29820
rect 39956 29764 40012 29820
rect 40060 29764 40116 29820
rect 59172 29764 59228 29820
rect 59276 29764 59332 29820
rect 59380 29764 59436 29820
rect 78492 29764 78548 29820
rect 78596 29764 78652 29820
rect 78700 29764 78756 29820
rect 10872 28980 10928 29036
rect 10976 28980 11032 29036
rect 11080 28980 11136 29036
rect 30192 28980 30248 29036
rect 30296 28980 30352 29036
rect 30400 28980 30456 29036
rect 49512 28980 49568 29036
rect 49616 28980 49672 29036
rect 49720 28980 49776 29036
rect 68832 28980 68888 29036
rect 68936 28980 68992 29036
rect 69040 28980 69096 29036
rect 20532 28196 20588 28252
rect 20636 28196 20692 28252
rect 20740 28196 20796 28252
rect 39852 28196 39908 28252
rect 39956 28196 40012 28252
rect 40060 28196 40116 28252
rect 59172 28196 59228 28252
rect 59276 28196 59332 28252
rect 59380 28196 59436 28252
rect 78492 28196 78548 28252
rect 78596 28196 78652 28252
rect 78700 28196 78756 28252
rect 10872 27412 10928 27468
rect 10976 27412 11032 27468
rect 11080 27412 11136 27468
rect 30192 27412 30248 27468
rect 30296 27412 30352 27468
rect 30400 27412 30456 27468
rect 49512 27412 49568 27468
rect 49616 27412 49672 27468
rect 49720 27412 49776 27468
rect 68832 27412 68888 27468
rect 68936 27412 68992 27468
rect 69040 27412 69096 27468
rect 20532 26628 20588 26684
rect 20636 26628 20692 26684
rect 20740 26628 20796 26684
rect 39852 26628 39908 26684
rect 39956 26628 40012 26684
rect 40060 26628 40116 26684
rect 59172 26628 59228 26684
rect 59276 26628 59332 26684
rect 59380 26628 59436 26684
rect 78492 26628 78548 26684
rect 78596 26628 78652 26684
rect 78700 26628 78756 26684
rect 10872 25844 10928 25900
rect 10976 25844 11032 25900
rect 11080 25844 11136 25900
rect 30192 25844 30248 25900
rect 30296 25844 30352 25900
rect 30400 25844 30456 25900
rect 49512 25844 49568 25900
rect 49616 25844 49672 25900
rect 49720 25844 49776 25900
rect 68832 25844 68888 25900
rect 68936 25844 68992 25900
rect 69040 25844 69096 25900
rect 20532 25060 20588 25116
rect 20636 25060 20692 25116
rect 20740 25060 20796 25116
rect 39852 25060 39908 25116
rect 39956 25060 40012 25116
rect 40060 25060 40116 25116
rect 59172 25060 59228 25116
rect 59276 25060 59332 25116
rect 59380 25060 59436 25116
rect 78492 25060 78548 25116
rect 78596 25060 78652 25116
rect 78700 25060 78756 25116
rect 10872 24276 10928 24332
rect 10976 24276 11032 24332
rect 11080 24276 11136 24332
rect 30192 24276 30248 24332
rect 30296 24276 30352 24332
rect 30400 24276 30456 24332
rect 49512 24276 49568 24332
rect 49616 24276 49672 24332
rect 49720 24276 49776 24332
rect 68832 24276 68888 24332
rect 68936 24276 68992 24332
rect 69040 24276 69096 24332
rect 20532 23492 20588 23548
rect 20636 23492 20692 23548
rect 20740 23492 20796 23548
rect 39852 23492 39908 23548
rect 39956 23492 40012 23548
rect 40060 23492 40116 23548
rect 59172 23492 59228 23548
rect 59276 23492 59332 23548
rect 59380 23492 59436 23548
rect 78492 23492 78548 23548
rect 78596 23492 78652 23548
rect 78700 23492 78756 23548
rect 10872 22708 10928 22764
rect 10976 22708 11032 22764
rect 11080 22708 11136 22764
rect 30192 22708 30248 22764
rect 30296 22708 30352 22764
rect 30400 22708 30456 22764
rect 49512 22708 49568 22764
rect 49616 22708 49672 22764
rect 49720 22708 49776 22764
rect 68832 22708 68888 22764
rect 68936 22708 68992 22764
rect 69040 22708 69096 22764
rect 20532 21924 20588 21980
rect 20636 21924 20692 21980
rect 20740 21924 20796 21980
rect 39852 21924 39908 21980
rect 39956 21924 40012 21980
rect 40060 21924 40116 21980
rect 59172 21924 59228 21980
rect 59276 21924 59332 21980
rect 59380 21924 59436 21980
rect 78492 21924 78548 21980
rect 78596 21924 78652 21980
rect 78700 21924 78756 21980
rect 10872 21140 10928 21196
rect 10976 21140 11032 21196
rect 11080 21140 11136 21196
rect 30192 21140 30248 21196
rect 30296 21140 30352 21196
rect 30400 21140 30456 21196
rect 49512 21140 49568 21196
rect 49616 21140 49672 21196
rect 49720 21140 49776 21196
rect 68832 21140 68888 21196
rect 68936 21140 68992 21196
rect 69040 21140 69096 21196
rect 20532 20356 20588 20412
rect 20636 20356 20692 20412
rect 20740 20356 20796 20412
rect 39852 20356 39908 20412
rect 39956 20356 40012 20412
rect 40060 20356 40116 20412
rect 59172 20356 59228 20412
rect 59276 20356 59332 20412
rect 59380 20356 59436 20412
rect 78492 20356 78548 20412
rect 78596 20356 78652 20412
rect 78700 20356 78756 20412
rect 10872 19572 10928 19628
rect 10976 19572 11032 19628
rect 11080 19572 11136 19628
rect 30192 19572 30248 19628
rect 30296 19572 30352 19628
rect 30400 19572 30456 19628
rect 49512 19572 49568 19628
rect 49616 19572 49672 19628
rect 49720 19572 49776 19628
rect 68832 19572 68888 19628
rect 68936 19572 68992 19628
rect 69040 19572 69096 19628
rect 20532 18788 20588 18844
rect 20636 18788 20692 18844
rect 20740 18788 20796 18844
rect 39852 18788 39908 18844
rect 39956 18788 40012 18844
rect 40060 18788 40116 18844
rect 59172 18788 59228 18844
rect 59276 18788 59332 18844
rect 59380 18788 59436 18844
rect 78492 18788 78548 18844
rect 78596 18788 78652 18844
rect 78700 18788 78756 18844
rect 10872 18004 10928 18060
rect 10976 18004 11032 18060
rect 11080 18004 11136 18060
rect 30192 18004 30248 18060
rect 30296 18004 30352 18060
rect 30400 18004 30456 18060
rect 49512 18004 49568 18060
rect 49616 18004 49672 18060
rect 49720 18004 49776 18060
rect 68832 18004 68888 18060
rect 68936 18004 68992 18060
rect 69040 18004 69096 18060
rect 20532 17220 20588 17276
rect 20636 17220 20692 17276
rect 20740 17220 20796 17276
rect 39852 17220 39908 17276
rect 39956 17220 40012 17276
rect 40060 17220 40116 17276
rect 59172 17220 59228 17276
rect 59276 17220 59332 17276
rect 59380 17220 59436 17276
rect 78492 17220 78548 17276
rect 78596 17220 78652 17276
rect 78700 17220 78756 17276
rect 10872 16436 10928 16492
rect 10976 16436 11032 16492
rect 11080 16436 11136 16492
rect 30192 16436 30248 16492
rect 30296 16436 30352 16492
rect 30400 16436 30456 16492
rect 49512 16436 49568 16492
rect 49616 16436 49672 16492
rect 49720 16436 49776 16492
rect 68832 16436 68888 16492
rect 68936 16436 68992 16492
rect 69040 16436 69096 16492
rect 20532 15652 20588 15708
rect 20636 15652 20692 15708
rect 20740 15652 20796 15708
rect 39852 15652 39908 15708
rect 39956 15652 40012 15708
rect 40060 15652 40116 15708
rect 59172 15652 59228 15708
rect 59276 15652 59332 15708
rect 59380 15652 59436 15708
rect 78492 15652 78548 15708
rect 78596 15652 78652 15708
rect 78700 15652 78756 15708
rect 10872 14868 10928 14924
rect 10976 14868 11032 14924
rect 11080 14868 11136 14924
rect 30192 14868 30248 14924
rect 30296 14868 30352 14924
rect 30400 14868 30456 14924
rect 49512 14868 49568 14924
rect 49616 14868 49672 14924
rect 49720 14868 49776 14924
rect 68832 14868 68888 14924
rect 68936 14868 68992 14924
rect 69040 14868 69096 14924
rect 20532 14084 20588 14140
rect 20636 14084 20692 14140
rect 20740 14084 20796 14140
rect 39852 14084 39908 14140
rect 39956 14084 40012 14140
rect 40060 14084 40116 14140
rect 59172 14084 59228 14140
rect 59276 14084 59332 14140
rect 59380 14084 59436 14140
rect 78492 14084 78548 14140
rect 78596 14084 78652 14140
rect 78700 14084 78756 14140
rect 10872 13300 10928 13356
rect 10976 13300 11032 13356
rect 11080 13300 11136 13356
rect 30192 13300 30248 13356
rect 30296 13300 30352 13356
rect 30400 13300 30456 13356
rect 49512 13300 49568 13356
rect 49616 13300 49672 13356
rect 49720 13300 49776 13356
rect 68832 13300 68888 13356
rect 68936 13300 68992 13356
rect 69040 13300 69096 13356
rect 20532 12516 20588 12572
rect 20636 12516 20692 12572
rect 20740 12516 20796 12572
rect 39852 12516 39908 12572
rect 39956 12516 40012 12572
rect 40060 12516 40116 12572
rect 59172 12516 59228 12572
rect 59276 12516 59332 12572
rect 59380 12516 59436 12572
rect 78492 12516 78548 12572
rect 78596 12516 78652 12572
rect 78700 12516 78756 12572
rect 10872 11732 10928 11788
rect 10976 11732 11032 11788
rect 11080 11732 11136 11788
rect 30192 11732 30248 11788
rect 30296 11732 30352 11788
rect 30400 11732 30456 11788
rect 49512 11732 49568 11788
rect 49616 11732 49672 11788
rect 49720 11732 49776 11788
rect 68832 11732 68888 11788
rect 68936 11732 68992 11788
rect 69040 11732 69096 11788
rect 20532 10948 20588 11004
rect 20636 10948 20692 11004
rect 20740 10948 20796 11004
rect 39852 10948 39908 11004
rect 39956 10948 40012 11004
rect 40060 10948 40116 11004
rect 10872 10164 10928 10220
rect 10976 10164 11032 10220
rect 11080 10164 11136 10220
rect 59172 10948 59228 11004
rect 59276 10948 59332 11004
rect 59380 10948 59436 11004
rect 78492 10948 78548 11004
rect 78596 10948 78652 11004
rect 78700 10948 78756 11004
rect 30192 10164 30248 10220
rect 30296 10164 30352 10220
rect 30400 10164 30456 10220
rect 49512 10164 49568 10220
rect 49616 10164 49672 10220
rect 49720 10164 49776 10220
rect 68832 10164 68888 10220
rect 68936 10164 68992 10220
rect 69040 10164 69096 10220
rect 20532 9380 20588 9436
rect 20636 9380 20692 9436
rect 20740 9380 20796 9436
rect 39852 9380 39908 9436
rect 39956 9380 40012 9436
rect 40060 9380 40116 9436
rect 59172 9380 59228 9436
rect 59276 9380 59332 9436
rect 59380 9380 59436 9436
rect 78492 9380 78548 9436
rect 78596 9380 78652 9436
rect 78700 9380 78756 9436
rect 10872 8596 10928 8652
rect 10976 8596 11032 8652
rect 11080 8596 11136 8652
rect 30192 8596 30248 8652
rect 30296 8596 30352 8652
rect 30400 8596 30456 8652
rect 49512 8596 49568 8652
rect 49616 8596 49672 8652
rect 49720 8596 49776 8652
rect 68832 8596 68888 8652
rect 68936 8596 68992 8652
rect 69040 8596 69096 8652
rect 20532 7812 20588 7868
rect 20636 7812 20692 7868
rect 20740 7812 20796 7868
rect 39852 7812 39908 7868
rect 39956 7812 40012 7868
rect 40060 7812 40116 7868
rect 59172 7812 59228 7868
rect 59276 7812 59332 7868
rect 59380 7812 59436 7868
rect 78492 7812 78548 7868
rect 78596 7812 78652 7868
rect 78700 7812 78756 7868
rect 10872 7028 10928 7084
rect 10976 7028 11032 7084
rect 11080 7028 11136 7084
rect 30192 7028 30248 7084
rect 30296 7028 30352 7084
rect 30400 7028 30456 7084
rect 49512 7028 49568 7084
rect 49616 7028 49672 7084
rect 49720 7028 49776 7084
rect 68832 7028 68888 7084
rect 68936 7028 68992 7084
rect 69040 7028 69096 7084
rect 20532 6244 20588 6300
rect 20636 6244 20692 6300
rect 20740 6244 20796 6300
rect 39852 6244 39908 6300
rect 39956 6244 40012 6300
rect 40060 6244 40116 6300
rect 59172 6244 59228 6300
rect 59276 6244 59332 6300
rect 59380 6244 59436 6300
rect 78492 6244 78548 6300
rect 78596 6244 78652 6300
rect 78700 6244 78756 6300
rect 10872 5460 10928 5516
rect 10976 5460 11032 5516
rect 11080 5460 11136 5516
rect 30192 5460 30248 5516
rect 30296 5460 30352 5516
rect 30400 5460 30456 5516
rect 49512 5460 49568 5516
rect 49616 5460 49672 5516
rect 49720 5460 49776 5516
rect 68832 5460 68888 5516
rect 68936 5460 68992 5516
rect 69040 5460 69096 5516
rect 20532 4676 20588 4732
rect 20636 4676 20692 4732
rect 20740 4676 20796 4732
rect 39852 4676 39908 4732
rect 39956 4676 40012 4732
rect 40060 4676 40116 4732
rect 59172 4676 59228 4732
rect 59276 4676 59332 4732
rect 59380 4676 59436 4732
rect 78492 4676 78548 4732
rect 78596 4676 78652 4732
rect 78700 4676 78756 4732
rect 10872 3892 10928 3948
rect 10976 3892 11032 3948
rect 11080 3892 11136 3948
rect 30192 3892 30248 3948
rect 30296 3892 30352 3948
rect 30400 3892 30456 3948
rect 49512 3892 49568 3948
rect 49616 3892 49672 3948
rect 49720 3892 49776 3948
rect 68832 3892 68888 3948
rect 68936 3892 68992 3948
rect 69040 3892 69096 3948
rect 20532 3108 20588 3164
rect 20636 3108 20692 3164
rect 20740 3108 20796 3164
rect 39852 3108 39908 3164
rect 39956 3108 40012 3164
rect 40060 3108 40116 3164
rect 59172 3108 59228 3164
rect 59276 3108 59332 3164
rect 59380 3108 59436 3164
rect 78492 3108 78548 3164
rect 78596 3108 78652 3164
rect 78700 3108 78756 3164
<< metal4 >>
rect 10844 36876 11164 36908
rect 10844 36820 10872 36876
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 11136 36820 11164 36876
rect 10844 35308 11164 36820
rect 10844 35252 10872 35308
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 11136 35252 11164 35308
rect 10844 33740 11164 35252
rect 10844 33684 10872 33740
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 11136 33684 11164 33740
rect 10844 32172 11164 33684
rect 10844 32116 10872 32172
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 11136 32116 11164 32172
rect 10844 30604 11164 32116
rect 10844 30548 10872 30604
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 11136 30548 11164 30604
rect 10844 29036 11164 30548
rect 10844 28980 10872 29036
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 11136 28980 11164 29036
rect 10844 27468 11164 28980
rect 10844 27412 10872 27468
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 11136 27412 11164 27468
rect 10844 25900 11164 27412
rect 10844 25844 10872 25900
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 11136 25844 11164 25900
rect 10844 24332 11164 25844
rect 10844 24276 10872 24332
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11136 24276 11164 24332
rect 10844 22764 11164 24276
rect 10844 22708 10872 22764
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 11136 22708 11164 22764
rect 10844 21196 11164 22708
rect 10844 21140 10872 21196
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 11136 21140 11164 21196
rect 10844 19628 11164 21140
rect 10844 19572 10872 19628
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 11136 19572 11164 19628
rect 10844 18060 11164 19572
rect 10844 18004 10872 18060
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 11136 18004 11164 18060
rect 10844 16492 11164 18004
rect 10844 16436 10872 16492
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11136 16436 11164 16492
rect 10844 14924 11164 16436
rect 10844 14868 10872 14924
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 11136 14868 11164 14924
rect 10844 13356 11164 14868
rect 10844 13300 10872 13356
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 11136 13300 11164 13356
rect 10844 11788 11164 13300
rect 10844 11732 10872 11788
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 11136 11732 11164 11788
rect 10844 10220 11164 11732
rect 10844 10164 10872 10220
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 11136 10164 11164 10220
rect 10844 8652 11164 10164
rect 10844 8596 10872 8652
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 11136 8596 11164 8652
rect 10844 7084 11164 8596
rect 10844 7028 10872 7084
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 11136 7028 11164 7084
rect 10844 5516 11164 7028
rect 10844 5460 10872 5516
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 11136 5460 11164 5516
rect 10844 3948 11164 5460
rect 10844 3892 10872 3948
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 11136 3892 11164 3948
rect 10844 3076 11164 3892
rect 20504 36092 20824 36908
rect 20504 36036 20532 36092
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20796 36036 20824 36092
rect 20504 34524 20824 36036
rect 20504 34468 20532 34524
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20796 34468 20824 34524
rect 20504 32956 20824 34468
rect 20504 32900 20532 32956
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20796 32900 20824 32956
rect 20504 31388 20824 32900
rect 20504 31332 20532 31388
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20796 31332 20824 31388
rect 20504 29820 20824 31332
rect 20504 29764 20532 29820
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20796 29764 20824 29820
rect 20504 28252 20824 29764
rect 20504 28196 20532 28252
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20796 28196 20824 28252
rect 20504 26684 20824 28196
rect 20504 26628 20532 26684
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20796 26628 20824 26684
rect 20504 25116 20824 26628
rect 20504 25060 20532 25116
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20796 25060 20824 25116
rect 20504 23548 20824 25060
rect 20504 23492 20532 23548
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20796 23492 20824 23548
rect 20504 21980 20824 23492
rect 20504 21924 20532 21980
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20796 21924 20824 21980
rect 20504 20412 20824 21924
rect 20504 20356 20532 20412
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20796 20356 20824 20412
rect 20504 18844 20824 20356
rect 20504 18788 20532 18844
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20796 18788 20824 18844
rect 20504 17276 20824 18788
rect 20504 17220 20532 17276
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20796 17220 20824 17276
rect 20504 15708 20824 17220
rect 20504 15652 20532 15708
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20796 15652 20824 15708
rect 20504 14140 20824 15652
rect 20504 14084 20532 14140
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20796 14084 20824 14140
rect 20504 12572 20824 14084
rect 20504 12516 20532 12572
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20796 12516 20824 12572
rect 20504 11004 20824 12516
rect 20504 10948 20532 11004
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20796 10948 20824 11004
rect 20504 9436 20824 10948
rect 20504 9380 20532 9436
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20796 9380 20824 9436
rect 20504 7868 20824 9380
rect 20504 7812 20532 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20796 7812 20824 7868
rect 20504 6300 20824 7812
rect 20504 6244 20532 6300
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20796 6244 20824 6300
rect 20504 4732 20824 6244
rect 20504 4676 20532 4732
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20796 4676 20824 4732
rect 20504 3164 20824 4676
rect 20504 3108 20532 3164
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20796 3108 20824 3164
rect 20504 3076 20824 3108
rect 30164 36876 30484 36908
rect 30164 36820 30192 36876
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30456 36820 30484 36876
rect 30164 35308 30484 36820
rect 30164 35252 30192 35308
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30456 35252 30484 35308
rect 30164 33740 30484 35252
rect 30164 33684 30192 33740
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30456 33684 30484 33740
rect 30164 32172 30484 33684
rect 30164 32116 30192 32172
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30456 32116 30484 32172
rect 30164 30604 30484 32116
rect 30164 30548 30192 30604
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30456 30548 30484 30604
rect 30164 29036 30484 30548
rect 30164 28980 30192 29036
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30456 28980 30484 29036
rect 30164 27468 30484 28980
rect 30164 27412 30192 27468
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30456 27412 30484 27468
rect 30164 25900 30484 27412
rect 30164 25844 30192 25900
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30456 25844 30484 25900
rect 30164 24332 30484 25844
rect 30164 24276 30192 24332
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30456 24276 30484 24332
rect 30164 22764 30484 24276
rect 30164 22708 30192 22764
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30456 22708 30484 22764
rect 30164 21196 30484 22708
rect 30164 21140 30192 21196
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30456 21140 30484 21196
rect 30164 19628 30484 21140
rect 30164 19572 30192 19628
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30456 19572 30484 19628
rect 30164 18060 30484 19572
rect 30164 18004 30192 18060
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30456 18004 30484 18060
rect 30164 16492 30484 18004
rect 30164 16436 30192 16492
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30456 16436 30484 16492
rect 30164 14924 30484 16436
rect 30164 14868 30192 14924
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30456 14868 30484 14924
rect 30164 13356 30484 14868
rect 30164 13300 30192 13356
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30456 13300 30484 13356
rect 30164 11788 30484 13300
rect 30164 11732 30192 11788
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30456 11732 30484 11788
rect 30164 10220 30484 11732
rect 30164 10164 30192 10220
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30456 10164 30484 10220
rect 30164 8652 30484 10164
rect 30164 8596 30192 8652
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30456 8596 30484 8652
rect 30164 7084 30484 8596
rect 30164 7028 30192 7084
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30456 7028 30484 7084
rect 30164 5516 30484 7028
rect 30164 5460 30192 5516
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30456 5460 30484 5516
rect 30164 3948 30484 5460
rect 30164 3892 30192 3948
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30456 3892 30484 3948
rect 30164 3076 30484 3892
rect 39824 36092 40144 36908
rect 39824 36036 39852 36092
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 40116 36036 40144 36092
rect 39824 34524 40144 36036
rect 39824 34468 39852 34524
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 40116 34468 40144 34524
rect 39824 32956 40144 34468
rect 39824 32900 39852 32956
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 40116 32900 40144 32956
rect 39824 31388 40144 32900
rect 39824 31332 39852 31388
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 40116 31332 40144 31388
rect 39824 29820 40144 31332
rect 39824 29764 39852 29820
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 40116 29764 40144 29820
rect 39824 28252 40144 29764
rect 39824 28196 39852 28252
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 40116 28196 40144 28252
rect 39824 26684 40144 28196
rect 39824 26628 39852 26684
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 40116 26628 40144 26684
rect 39824 25116 40144 26628
rect 39824 25060 39852 25116
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 40116 25060 40144 25116
rect 39824 23548 40144 25060
rect 39824 23492 39852 23548
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 40116 23492 40144 23548
rect 39824 21980 40144 23492
rect 39824 21924 39852 21980
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 40116 21924 40144 21980
rect 39824 20412 40144 21924
rect 39824 20356 39852 20412
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 40116 20356 40144 20412
rect 39824 18844 40144 20356
rect 39824 18788 39852 18844
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 40116 18788 40144 18844
rect 39824 17276 40144 18788
rect 39824 17220 39852 17276
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40116 17220 40144 17276
rect 39824 15708 40144 17220
rect 39824 15652 39852 15708
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40116 15652 40144 15708
rect 39824 14140 40144 15652
rect 39824 14084 39852 14140
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 40116 14084 40144 14140
rect 39824 12572 40144 14084
rect 39824 12516 39852 12572
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 40116 12516 40144 12572
rect 39824 11004 40144 12516
rect 39824 10948 39852 11004
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 40116 10948 40144 11004
rect 39824 9436 40144 10948
rect 39824 9380 39852 9436
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 40116 9380 40144 9436
rect 39824 7868 40144 9380
rect 39824 7812 39852 7868
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 40116 7812 40144 7868
rect 39824 6300 40144 7812
rect 39824 6244 39852 6300
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 40116 6244 40144 6300
rect 39824 4732 40144 6244
rect 39824 4676 39852 4732
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 40116 4676 40144 4732
rect 39824 3164 40144 4676
rect 39824 3108 39852 3164
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 40116 3108 40144 3164
rect 39824 3076 40144 3108
rect 49484 36876 49804 36908
rect 49484 36820 49512 36876
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49776 36820 49804 36876
rect 49484 35308 49804 36820
rect 49484 35252 49512 35308
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49776 35252 49804 35308
rect 49484 33740 49804 35252
rect 49484 33684 49512 33740
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49776 33684 49804 33740
rect 49484 32172 49804 33684
rect 49484 32116 49512 32172
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49776 32116 49804 32172
rect 49484 30604 49804 32116
rect 49484 30548 49512 30604
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49776 30548 49804 30604
rect 49484 29036 49804 30548
rect 49484 28980 49512 29036
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49776 28980 49804 29036
rect 49484 27468 49804 28980
rect 49484 27412 49512 27468
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49776 27412 49804 27468
rect 49484 25900 49804 27412
rect 49484 25844 49512 25900
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49776 25844 49804 25900
rect 49484 24332 49804 25844
rect 49484 24276 49512 24332
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49776 24276 49804 24332
rect 49484 22764 49804 24276
rect 49484 22708 49512 22764
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49776 22708 49804 22764
rect 49484 21196 49804 22708
rect 49484 21140 49512 21196
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49776 21140 49804 21196
rect 49484 19628 49804 21140
rect 49484 19572 49512 19628
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49776 19572 49804 19628
rect 49484 18060 49804 19572
rect 49484 18004 49512 18060
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49776 18004 49804 18060
rect 49484 16492 49804 18004
rect 49484 16436 49512 16492
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49776 16436 49804 16492
rect 49484 14924 49804 16436
rect 49484 14868 49512 14924
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49776 14868 49804 14924
rect 49484 13356 49804 14868
rect 49484 13300 49512 13356
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49776 13300 49804 13356
rect 49484 11788 49804 13300
rect 49484 11732 49512 11788
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49776 11732 49804 11788
rect 49484 10220 49804 11732
rect 49484 10164 49512 10220
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49776 10164 49804 10220
rect 49484 8652 49804 10164
rect 49484 8596 49512 8652
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49776 8596 49804 8652
rect 49484 7084 49804 8596
rect 49484 7028 49512 7084
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49776 7028 49804 7084
rect 49484 5516 49804 7028
rect 49484 5460 49512 5516
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49776 5460 49804 5516
rect 49484 3948 49804 5460
rect 49484 3892 49512 3948
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49776 3892 49804 3948
rect 49484 3076 49804 3892
rect 59144 36092 59464 36908
rect 59144 36036 59172 36092
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59436 36036 59464 36092
rect 59144 34524 59464 36036
rect 59144 34468 59172 34524
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59436 34468 59464 34524
rect 59144 32956 59464 34468
rect 59144 32900 59172 32956
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59436 32900 59464 32956
rect 59144 31388 59464 32900
rect 59144 31332 59172 31388
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59436 31332 59464 31388
rect 59144 29820 59464 31332
rect 59144 29764 59172 29820
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59436 29764 59464 29820
rect 59144 28252 59464 29764
rect 59144 28196 59172 28252
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59436 28196 59464 28252
rect 59144 26684 59464 28196
rect 59144 26628 59172 26684
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59436 26628 59464 26684
rect 59144 25116 59464 26628
rect 59144 25060 59172 25116
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59436 25060 59464 25116
rect 59144 23548 59464 25060
rect 59144 23492 59172 23548
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59436 23492 59464 23548
rect 59144 21980 59464 23492
rect 59144 21924 59172 21980
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59436 21924 59464 21980
rect 59144 20412 59464 21924
rect 59144 20356 59172 20412
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59436 20356 59464 20412
rect 59144 18844 59464 20356
rect 59144 18788 59172 18844
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59436 18788 59464 18844
rect 59144 17276 59464 18788
rect 59144 17220 59172 17276
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59436 17220 59464 17276
rect 59144 15708 59464 17220
rect 59144 15652 59172 15708
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59436 15652 59464 15708
rect 59144 14140 59464 15652
rect 59144 14084 59172 14140
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59436 14084 59464 14140
rect 59144 12572 59464 14084
rect 59144 12516 59172 12572
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59436 12516 59464 12572
rect 59144 11004 59464 12516
rect 59144 10948 59172 11004
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59436 10948 59464 11004
rect 59144 9436 59464 10948
rect 59144 9380 59172 9436
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59436 9380 59464 9436
rect 59144 7868 59464 9380
rect 59144 7812 59172 7868
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59436 7812 59464 7868
rect 59144 6300 59464 7812
rect 59144 6244 59172 6300
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59436 6244 59464 6300
rect 59144 4732 59464 6244
rect 59144 4676 59172 4732
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59436 4676 59464 4732
rect 59144 3164 59464 4676
rect 59144 3108 59172 3164
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59436 3108 59464 3164
rect 59144 3076 59464 3108
rect 68804 36876 69124 36908
rect 68804 36820 68832 36876
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 69096 36820 69124 36876
rect 68804 35308 69124 36820
rect 68804 35252 68832 35308
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 69096 35252 69124 35308
rect 68804 33740 69124 35252
rect 68804 33684 68832 33740
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 69096 33684 69124 33740
rect 68804 32172 69124 33684
rect 68804 32116 68832 32172
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 69096 32116 69124 32172
rect 68804 30604 69124 32116
rect 68804 30548 68832 30604
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 69096 30548 69124 30604
rect 68804 29036 69124 30548
rect 68804 28980 68832 29036
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 69096 28980 69124 29036
rect 68804 27468 69124 28980
rect 68804 27412 68832 27468
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69096 27412 69124 27468
rect 68804 25900 69124 27412
rect 68804 25844 68832 25900
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 69096 25844 69124 25900
rect 68804 24332 69124 25844
rect 68804 24276 68832 24332
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 69096 24276 69124 24332
rect 68804 22764 69124 24276
rect 68804 22708 68832 22764
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 69096 22708 69124 22764
rect 68804 21196 69124 22708
rect 68804 21140 68832 21196
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 69096 21140 69124 21196
rect 68804 19628 69124 21140
rect 68804 19572 68832 19628
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 69096 19572 69124 19628
rect 68804 18060 69124 19572
rect 68804 18004 68832 18060
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 69096 18004 69124 18060
rect 68804 16492 69124 18004
rect 68804 16436 68832 16492
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 69096 16436 69124 16492
rect 68804 14924 69124 16436
rect 68804 14868 68832 14924
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 69096 14868 69124 14924
rect 68804 13356 69124 14868
rect 68804 13300 68832 13356
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 69096 13300 69124 13356
rect 68804 11788 69124 13300
rect 68804 11732 68832 11788
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 69096 11732 69124 11788
rect 68804 10220 69124 11732
rect 68804 10164 68832 10220
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 69096 10164 69124 10220
rect 68804 8652 69124 10164
rect 68804 8596 68832 8652
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 69096 8596 69124 8652
rect 68804 7084 69124 8596
rect 68804 7028 68832 7084
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 69096 7028 69124 7084
rect 68804 5516 69124 7028
rect 68804 5460 68832 5516
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 69096 5460 69124 5516
rect 68804 3948 69124 5460
rect 68804 3892 68832 3948
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 69096 3892 69124 3948
rect 68804 3076 69124 3892
rect 78464 36092 78784 36908
rect 78464 36036 78492 36092
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78756 36036 78784 36092
rect 78464 34524 78784 36036
rect 78464 34468 78492 34524
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78756 34468 78784 34524
rect 78464 32956 78784 34468
rect 78464 32900 78492 32956
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78756 32900 78784 32956
rect 78464 31388 78784 32900
rect 78464 31332 78492 31388
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78756 31332 78784 31388
rect 78464 29820 78784 31332
rect 78464 29764 78492 29820
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78756 29764 78784 29820
rect 78464 28252 78784 29764
rect 78464 28196 78492 28252
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78756 28196 78784 28252
rect 78464 26684 78784 28196
rect 78464 26628 78492 26684
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78756 26628 78784 26684
rect 78464 25116 78784 26628
rect 78464 25060 78492 25116
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78756 25060 78784 25116
rect 78464 23548 78784 25060
rect 78464 23492 78492 23548
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78756 23492 78784 23548
rect 78464 21980 78784 23492
rect 78464 21924 78492 21980
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78756 21924 78784 21980
rect 78464 20412 78784 21924
rect 78464 20356 78492 20412
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78756 20356 78784 20412
rect 78464 18844 78784 20356
rect 78464 18788 78492 18844
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78756 18788 78784 18844
rect 78464 17276 78784 18788
rect 78464 17220 78492 17276
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78756 17220 78784 17276
rect 78464 15708 78784 17220
rect 78464 15652 78492 15708
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78756 15652 78784 15708
rect 78464 14140 78784 15652
rect 78464 14084 78492 14140
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78756 14084 78784 14140
rect 78464 12572 78784 14084
rect 78464 12516 78492 12572
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78756 12516 78784 12572
rect 78464 11004 78784 12516
rect 78464 10948 78492 11004
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78756 10948 78784 11004
rect 78464 9436 78784 10948
rect 78464 9380 78492 9436
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78756 9380 78784 9436
rect 78464 7868 78784 9380
rect 78464 7812 78492 7868
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78756 7812 78784 7868
rect 78464 6300 78784 7812
rect 78464 6244 78492 6300
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78756 6244 78784 6300
rect 78464 4732 78784 6244
rect 78464 4676 78492 4732
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78756 4676 78784 4732
rect 78464 3164 78784 4676
rect 78464 3108 78492 3164
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78756 3108 78784 3164
rect 78464 3076 78784 3108
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 69888 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _189_
timestamp 1698431365
transform -1 0 55328 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 52192 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _191_
timestamp 1698431365
transform 1 0 69888 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44576 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _193_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _194_
timestamp 1698431365
transform -1 0 21840 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1698431365
transform -1 0 40992 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _196_
timestamp 1698431365
transform -1 0 42672 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _197_
timestamp 1698431365
transform 1 0 55328 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _198_
timestamp 1698431365
transform -1 0 58240 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _199_
timestamp 1698431365
transform 1 0 6048 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _200_
timestamp 1698431365
transform -1 0 53424 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _201_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 56224 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _202_
timestamp 1698431365
transform -1 0 55776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _203_
timestamp 1698431365
transform -1 0 65856 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _204_
timestamp 1698431365
transform -1 0 62048 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 64176 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _206_
timestamp 1698431365
transform -1 0 64064 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 62720 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _208_
timestamp 1698431365
transform -1 0 65184 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _209_
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 67872 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _211_
timestamp 1698431365
transform -1 0 67088 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _212_
timestamp 1698431365
transform 1 0 59136 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _213_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 63168 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _214_
timestamp 1698431365
transform -1 0 64064 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _215_
timestamp 1698431365
transform 1 0 60816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _216_
timestamp 1698431365
transform -1 0 60816 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _217_
timestamp 1698431365
transform -1 0 59808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _218_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 59360 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _219_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 55664 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _220_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _222_
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _223_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30800 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _224_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24752 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _225_
timestamp 1698431365
transform -1 0 24864 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _226_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _227_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _228_
timestamp 1698431365
transform -1 0 29680 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _229_
timestamp 1698431365
transform -1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _230_
timestamp 1698431365
transform -1 0 57232 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _231_
timestamp 1698431365
transform -1 0 27888 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _232_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30352 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _233_
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _234_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 3136
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _235_
timestamp 1698431365
transform -1 0 26208 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _236_
timestamp 1698431365
transform -1 0 58352 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _237_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _238_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _239_
timestamp 1698431365
transform 1 0 22960 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _240_
timestamp 1698431365
transform 1 0 25536 0 1 3136
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _241_
timestamp 1698431365
transform -1 0 26096 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _242_
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _243_
timestamp 1698431365
transform -1 0 58912 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _244_
timestamp 1698431365
transform 1 0 26208 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _245_
timestamp 1698431365
transform -1 0 30464 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _246_
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _247_
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _248_
timestamp 1698431365
transform -1 0 26768 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _249_
timestamp 1698431365
transform -1 0 55104 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _250_
timestamp 1698431365
transform -1 0 54208 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _251_
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _252_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _253_
timestamp 1698431365
transform -1 0 34720 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _254_
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _255_
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _256_
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _257_
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _258_
timestamp 1698431365
transform -1 0 32704 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _259_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _260_
timestamp 1698431365
transform -1 0 57120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _261_
timestamp 1698431365
transform 1 0 35728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _262_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _263_
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _264_
timestamp 1698431365
transform -1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _265_
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _266_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _267_
timestamp 1698431365
transform -1 0 34944 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _268_
timestamp 1698431365
transform -1 0 52416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _269_
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _270_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _271_
timestamp 1698431365
transform 1 0 39424 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _272_
timestamp 1698431365
transform -1 0 33712 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _273_
timestamp 1698431365
transform -1 0 46144 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _274_
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _275_
timestamp 1698431365
transform 1 0 24864 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _276_
timestamp 1698431365
transform 1 0 41440 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _277_
timestamp 1698431365
transform -1 0 37520 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _278_
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _279_
timestamp 1698431365
transform 1 0 44688 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _280_
timestamp 1698431365
transform -1 0 43680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _281_
timestamp 1698431365
transform 1 0 39200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _282_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34720 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _283_
timestamp 1698431365
transform 1 0 38304 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _284_
timestamp 1698431365
transform 1 0 39200 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _285_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _286_
timestamp 1698431365
transform -1 0 50736 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _287_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41440 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _288_
timestamp 1698431365
transform -1 0 38416 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _289_
timestamp 1698431365
transform -1 0 37632 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _290_
timestamp 1698431365
transform 1 0 36736 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _291_
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _292_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _293_
timestamp 1698431365
transform 1 0 42112 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _294_
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _295_
timestamp 1698431365
transform 1 0 47712 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _296_
timestamp 1698431365
transform 1 0 39424 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _297_
timestamp 1698431365
transform 1 0 47040 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _298_
timestamp 1698431365
transform 1 0 48496 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _299_
timestamp 1698431365
transform 1 0 51408 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _300_
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _301_
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _302_
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _303_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38304 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _304_
timestamp 1698431365
transform -1 0 41440 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _305_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37632 0 1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _306_
timestamp 1698431365
transform -1 0 41440 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _307_
timestamp 1698431365
transform 1 0 50288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _308_
timestamp 1698431365
transform 1 0 50624 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _309_
timestamp 1698431365
transform -1 0 50960 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _310_
timestamp 1698431365
transform 1 0 58464 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _311_
timestamp 1698431365
transform -1 0 49504 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _312_
timestamp 1698431365
transform -1 0 47712 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _313_
timestamp 1698431365
transform 1 0 45472 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _314_
timestamp 1698431365
transform -1 0 49280 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _315_
timestamp 1698431365
transform -1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _316_
timestamp 1698431365
transform -1 0 40544 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _317_
timestamp 1698431365
transform 1 0 41104 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _318_
timestamp 1698431365
transform -1 0 45472 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _319_
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _320_
timestamp 1698431365
transform 1 0 52416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _321_
timestamp 1698431365
transform 1 0 43680 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _322_
timestamp 1698431365
transform -1 0 43568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _323_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42672 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _324_
timestamp 1698431365
transform -1 0 48384 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _325_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _326_
timestamp 1698431365
transform -1 0 45360 0 1 3136
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _327_
timestamp 1698431365
transform 1 0 55776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _328_
timestamp 1698431365
transform 1 0 43344 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _329_
timestamp 1698431365
transform -1 0 44464 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _330_
timestamp 1698431365
transform 1 0 58912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _331_
timestamp 1698431365
transform 1 0 45360 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _332_
timestamp 1698431365
transform 1 0 46368 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _333_
timestamp 1698431365
transform -1 0 48160 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _334_
timestamp 1698431365
transform -1 0 18704 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _335_
timestamp 1698431365
transform -1 0 19824 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _336_
timestamp 1698431365
transform -1 0 17472 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _337_
timestamp 1698431365
transform -1 0 18144 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _338_
timestamp 1698431365
transform 1 0 15008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _339_
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _340_
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _341_
timestamp 1698431365
transform 1 0 7504 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _342_
timestamp 1698431365
transform 1 0 7952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _343_
timestamp 1698431365
transform -1 0 15008 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _344_
timestamp 1698431365
transform 1 0 12208 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _345_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _346_
timestamp 1698431365
transform 1 0 10864 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _347_
timestamp 1698431365
transform -1 0 10864 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _348_
timestamp 1698431365
transform 1 0 10976 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _349_
timestamp 1698431365
transform -1 0 10752 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _350_
timestamp 1698431365
transform 1 0 11760 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _351_
timestamp 1698431365
transform -1 0 11760 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _352_
timestamp 1698431365
transform 1 0 13888 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _353_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _354_
timestamp 1698431365
transform 1 0 14896 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _355_
timestamp 1698431365
transform 1 0 19936 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _356_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _357_
timestamp 1698431365
transform 1 0 19264 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _358_
timestamp 1698431365
transform 1 0 19152 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _359_
timestamp 1698431365
transform -1 0 19712 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _360_
timestamp 1698431365
transform -1 0 20608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _361_
timestamp 1698431365
transform -1 0 17920 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _362_
timestamp 1698431365
transform -1 0 16464 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _363_
timestamp 1698431365
transform 1 0 22288 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _364_
timestamp 1698431365
transform -1 0 22400 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _365_
timestamp 1698431365
transform 1 0 17360 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _366_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _367_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _368_
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _369_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _370_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _371_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _372_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _373_
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _374_
timestamp 1698431365
transform 1 0 24192 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _375_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _376_
timestamp 1698431365
transform -1 0 35728 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _377_
timestamp 1698431365
transform -1 0 33152 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _378_
timestamp 1698431365
transform -1 0 36624 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _379_
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _380_
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _381_
timestamp 1698431365
transform -1 0 42000 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _382_
timestamp 1698431365
transform -1 0 53312 0 -1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _383_
timestamp 1698431365
transform -1 0 53200 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _384_
timestamp 1698431365
transform -1 0 50288 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _385_
timestamp 1698431365
transform -1 0 45024 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _386_
timestamp 1698431365
transform -1 0 45696 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _387_
timestamp 1698431365
transform -1 0 49392 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _388_
timestamp 1698431365
transform -1 0 19152 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _389_
timestamp 1698431365
transform 1 0 6832 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _390_
timestamp 1698431365
transform -1 0 10192 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _391_
timestamp 1698431365
transform -1 0 14000 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _392_
timestamp 1698431365
transform 1 0 8960 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _393_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _394_
timestamp 1698431365
transform 1 0 9856 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _395_
timestamp 1698431365
transform 1 0 13440 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _396_
timestamp 1698431365
transform -1 0 22960 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _397_
timestamp 1698431365
transform -1 0 21280 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _398_
timestamp 1698431365
transform -1 0 22176 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _399_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _400_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _401_
timestamp 1698431365
transform 1 0 15232 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _402_
timestamp 1698431365
transform 1 0 13552 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _403_
timestamp 1698431365
transform -1 0 26544 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 69888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1698431365
transform 1 0 59472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I
timestamp 1698431365
transform 1 0 54544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A1
timestamp 1698431365
transform 1 0 60592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A2
timestamp 1698431365
transform -1 0 54096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I1
timestamp 1698431365
transform -1 0 69104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__A2
timestamp 1698431365
transform -1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I
timestamp 1698431365
transform -1 0 22848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1698431365
transform -1 0 42112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1698431365
transform 1 0 42784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__A2
timestamp 1698431365
transform -1 0 56896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1698431365
transform 1 0 65408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I
timestamp 1698431365
transform 1 0 61152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__B2
timestamp 1698431365
transform -1 0 63616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__B2
timestamp 1698431365
transform -1 0 64288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I
timestamp 1698431365
transform 1 0 62496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1698431365
transform 1 0 64512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__B2
timestamp 1698431365
transform 1 0 60144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__A1
timestamp 1698431365
transform -1 0 65184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__A2
timestamp 1698431365
transform -1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__B1
timestamp 1698431365
transform 1 0 60816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__B2
timestamp 1698431365
transform 1 0 61264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__A1
timestamp 1698431365
transform -1 0 60032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__A1
timestamp 1698431365
transform 1 0 61040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__A2
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__B
timestamp 1698431365
transform -1 0 38752 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__I
timestamp 1698431365
transform -1 0 23744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I
timestamp 1698431365
transform -1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__I
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__A1
timestamp 1698431365
transform -1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A1
timestamp 1698431365
transform -1 0 27888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A2
timestamp 1698431365
transform -1 0 28336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__I
timestamp 1698431365
transform -1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A2
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A1
timestamp 1698431365
transform -1 0 10752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__A1
timestamp 1698431365
transform -1 0 28448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__A2
timestamp 1698431365
transform -1 0 28896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A1
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__A2
timestamp 1698431365
transform -1 0 23184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A1
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A1
timestamp 1698431365
transform -1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__A1
timestamp 1698431365
transform -1 0 27664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__A2
timestamp 1698431365
transform -1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__A1
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__A2
timestamp 1698431365
transform 1 0 27216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__A3
timestamp 1698431365
transform 1 0 26656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__A1
timestamp 1698431365
transform 1 0 30464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A1
timestamp 1698431365
transform -1 0 27440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A2
timestamp 1698431365
transform -1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__A1
timestamp 1698431365
transform 1 0 26768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I
timestamp 1698431365
transform 1 0 34160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__A3
timestamp 1698431365
transform -1 0 31136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__A4
timestamp 1698431365
transform 1 0 31360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__A1
timestamp 1698431365
transform -1 0 26992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I
timestamp 1698431365
transform -1 0 25984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I
timestamp 1698431365
transform -1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__A1
timestamp 1698431365
transform 1 0 30128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__A1
timestamp 1698431365
transform -1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__A2
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A1
timestamp 1698431365
transform 1 0 31808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A1
timestamp 1698431365
transform 1 0 34384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A2
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__A1
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__B
timestamp 1698431365
transform -1 0 31808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A1
timestamp 1698431365
transform -1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__A2
timestamp 1698431365
transform -1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A1
timestamp 1698431365
transform 1 0 59920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A1
timestamp 1698431365
transform 1 0 26320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A2
timestamp 1698431365
transform -1 0 26544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__A1
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__A1
timestamp 1698431365
transform 1 0 49840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__A2
timestamp 1698431365
transform 1 0 51856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__A1
timestamp 1698431365
transform -1 0 26992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__A2
timestamp 1698431365
transform 1 0 43792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__A2
timestamp 1698431365
transform 1 0 50288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__B
timestamp 1698431365
transform 1 0 52752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A1
timestamp 1698431365
transform 1 0 37184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A2
timestamp 1698431365
transform 1 0 29232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1698431365
transform 1 0 40880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A1
timestamp 1698431365
transform 1 0 52304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A2
timestamp 1698431365
transform 1 0 49840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A2
timestamp 1698431365
transform 1 0 44240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__C2
timestamp 1698431365
transform 1 0 43904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A1
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A2
timestamp 1698431365
transform 1 0 37968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A1
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A2
timestamp 1698431365
transform 1 0 46816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__B2
timestamp 1698431365
transform 1 0 44800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1698431365
transform 1 0 48048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A1
timestamp 1698431365
transform 1 0 56672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__C2
timestamp 1698431365
transform 1 0 52976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A1
timestamp 1698431365
transform 1 0 58912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A1
timestamp 1698431365
transform 1 0 53872 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__B
timestamp 1698431365
transform 1 0 50288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__I
timestamp 1698431365
transform 1 0 38528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__I
timestamp 1698431365
transform -1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A1
timestamp 1698431365
transform 1 0 41552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A2
timestamp 1698431365
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__C2
timestamp 1698431365
transform 1 0 52528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__A1
timestamp 1698431365
transform 1 0 61040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A1
timestamp 1698431365
transform -1 0 48720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__C2
timestamp 1698431365
transform 1 0 53200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A1
timestamp 1698431365
transform 1 0 44352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__A1
timestamp 1698431365
transform -1 0 41216 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__A1
timestamp 1698431365
transform -1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A1
timestamp 1698431365
transform 1 0 54992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__B2
timestamp 1698431365
transform 1 0 49392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__A1
timestamp 1698431365
transform -1 0 45696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A1
timestamp 1698431365
transform 1 0 57120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__B2
timestamp 1698431365
transform 1 0 47264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__A1
timestamp 1698431365
transform -1 0 60816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__A1
timestamp 1698431365
transform 1 0 50064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__C2
timestamp 1698431365
transform 1 0 48832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__I
timestamp 1698431365
transform -1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__I1
timestamp 1698431365
transform -1 0 7952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__I1
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__I1
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I1
timestamp 1698431365
transform 1 0 13328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I1
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I1
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__I1
timestamp 1698431365
transform 1 0 15792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__A1
timestamp 1698431365
transform -1 0 22288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I1
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__A1
timestamp 1698431365
transform -1 0 18928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A1
timestamp 1698431365
transform -1 0 13888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__I1
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A1
timestamp 1698431365
transform 1 0 17920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A1
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__I1
timestamp 1698431365
transform -1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__CLK
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__CLK
timestamp 1698431365
transform 1 0 27216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__CLK
timestamp 1698431365
transform -1 0 24192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__CLK
timestamp 1698431365
transform 1 0 41440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__CLK
timestamp 1698431365
transform 1 0 49840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__CLK
timestamp 1698431365
transform 1 0 53424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__CLK
timestamp 1698431365
transform 1 0 49616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__CLK
timestamp 1698431365
transform -1 0 45248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__CLK
timestamp 1698431365
transform -1 0 45696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__CLK
timestamp 1698431365
transform 1 0 45136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__CLK
timestamp 1698431365
transform 1 0 18256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__CLK
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__CLK
timestamp 1698431365
transform -1 0 6048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__CLK
timestamp 1698431365
transform 1 0 14000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__CLK
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__CLK
timestamp 1698431365
transform -1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__CLK
timestamp 1698431365
transform 1 0 22512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__CLK
timestamp 1698431365
transform 1 0 21504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__CLK
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__CLK
timestamp 1698431365
transform 1 0 24416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__CLK
timestamp 1698431365
transform 1 0 18704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__CLK
timestamp 1698431365
transform 1 0 23072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_counter.clk_I
timestamp 1698431365
transform 1 0 30576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_counter.clk_I
timestamp 1698431365
transform -1 0 17808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_counter.clk_I
timestamp 1698431365
transform 1 0 27664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_counter.clk_I
timestamp 1698431365
transform 1 0 40768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_counter.clk_I
timestamp 1698431365
transform -1 0 33376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold1_I
timestamp 1698431365
transform -1 0 71792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold5_I
timestamp 1698431365
transform 1 0 74144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold9_I
timestamp 1698431365
transform 1 0 69104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold10_I
timestamp 1698431365
transform 1 0 59360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold13_I
timestamp 1698431365
transform 1 0 76944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold17_I
timestamp 1698431365
transform -1 0 73920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold18_I
timestamp 1698431365
transform 1 0 63056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold21_I
timestamp 1698431365
transform -1 0 72240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold25_I
timestamp 1698431365
transform 1 0 74592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold29_I
timestamp 1698431365
transform -1 0 66864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold33_I
timestamp 1698431365
transform -1 0 66304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold34_I
timestamp 1698431365
transform 1 0 57568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold37_I
timestamp 1698431365
transform 1 0 70672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold38_I
timestamp 1698431365
transform -1 0 50960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold41_I
timestamp 1698431365
transform 1 0 72800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold45_I
timestamp 1698431365
transform -1 0 68880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold49_I
timestamp 1698431365
transform -1 0 61824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold50_I
timestamp 1698431365
transform -1 0 57344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold53_I
timestamp 1698431365
transform -1 0 62608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold54_I
timestamp 1698431365
transform -1 0 53648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold57_I
timestamp 1698431365
transform -1 0 68208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold61_I
timestamp 1698431365
transform -1 0 70000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold65_I
timestamp 1698431365
transform -1 0 76048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold68_I
timestamp 1698431365
transform 1 0 74928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold69_I
timestamp 1698431365
transform -1 0 67760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold71_I
timestamp 1698431365
transform 1 0 72912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold72_I
timestamp 1698431365
transform 1 0 72464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold74_I
timestamp 1698431365
transform -1 0 71344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold75_I
timestamp 1698431365
transform -1 0 75264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold76_I
timestamp 1698431365
transform -1 0 70448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold77_I
timestamp 1698431365
transform 1 0 73248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold79_I
timestamp 1698431365
transform -1 0 62496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold80_I
timestamp 1698431365
transform -1 0 69552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold81_I
timestamp 1698431365
transform -1 0 60928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold82_I
timestamp 1698431365
transform 1 0 75376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold83_I
timestamp 1698431365
transform -1 0 64848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold84_I
timestamp 1698431365
transform -1 0 66304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold85_I
timestamp 1698431365
transform -1 0 68656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold86_I
timestamp 1698431365
transform -1 0 67088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold87_I
timestamp 1698431365
transform -1 0 73920 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 76720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 77728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 3472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 3024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 4592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 18592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 17808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 3920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 4368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform 1 0 19152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 7504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 10080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform -1 0 2576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform -1 0 13104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform -1 0 14224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 2128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 2016 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 2016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 5600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output60_I
timestamp 1698431365
transform 1 0 44912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1698431365
transform 1 0 49280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1698431365
transform 1 0 50288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output68_I
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output70_I
timestamp 1698431365
transform -1 0 27552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output72_I
timestamp 1698431365
transform -1 0 33824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output74_I
timestamp 1698431365
transform 1 0 27776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output75_I
timestamp 1698431365
transform 1 0 6272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_counter.clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34608 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_counter.clk
timestamp 1698431365
transform -1 0 23408 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_counter.clk
timestamp 1698431365
transform 1 0 18928 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_counter.clk
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_counter.clk
timestamp 1698431365
transform -1 0 39312 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout92
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout93
timestamp 1698431365
transform -1 0 32704 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout94
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_168
timestamp 1698431365
transform 1 0 20160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_393 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45360 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_416
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698431365
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_472
timestamp 1698431365
transform 1 0 54208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_498
timestamp 1698431365
transform 1 0 57120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_509
timestamp 1698431365
transform 1 0 58352 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_512
timestamp 1698431365
transform 1 0 58688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_539
timestamp 1698431365
transform 1 0 61712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_546
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_611
timestamp 1698431365
transform 1 0 69776 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_639
timestamp 1698431365
transform 1 0 72912 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_679
timestamp 1698431365
transform 1 0 77392 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_80
timestamp 1698431365
transform 1 0 10304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_113
timestamp 1698431365
transform 1 0 14000 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_152
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_191
timestamp 1698431365
transform 1 0 22736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_237
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_461
timestamp 1698431365
transform 1 0 52976 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_471
timestamp 1698431365
transform 1 0 54096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_499
timestamp 1698431365
transform 1 0 57232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_542
timestamp 1698431365
transform 1 0 62048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_628
timestamp 1698431365
transform 1 0 71680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_4
timestamp 1698431365
transform 1 0 1792 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_7
timestamp 1698431365
transform 1 0 2128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_11
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_15
timestamp 1698431365
transform 1 0 3024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_19
timestamp 1698431365
transform 1 0 3472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_23
timestamp 1698431365
transform 1 0 3920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_39
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_203
timestamp 1698431365
transform 1 0 24080 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_220
timestamp 1698431365
transform 1 0 25984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_225
timestamp 1698431365
transform 1 0 26544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_336
timestamp 1698431365
transform 1 0 38976 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_363
timestamp 1698431365
transform 1 0 42000 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_373
timestamp 1698431365
transform 1 0 43120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_400
timestamp 1698431365
transform 1 0 46144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_404
timestamp 1698431365
transform 1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_408
timestamp 1698431365
transform 1 0 47040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_412
timestamp 1698431365
transform 1 0 47488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_414
timestamp 1698431365
transform 1 0 47712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_427
timestamp 1698431365
transform 1 0 49168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_431
timestamp 1698431365
transform 1 0 49616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_435
timestamp 1698431365
transform 1 0 50064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_515
timestamp 1698431365
transform 1 0 59024 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_527
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_531
timestamp 1698431365
transform 1 0 60816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_535
timestamp 1698431365
transform 1 0 61264 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_593
timestamp 1698431365
transform 1 0 67760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_663
timestamp 1698431365
transform 1 0 75600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_687
timestamp 1698431365
transform 1 0 78288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_87
timestamp 1698431365
transform 1 0 11088 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_229
timestamp 1698431365
transform 1 0 26992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_231
timestamp 1698431365
transform 1 0 27216 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_234
timestamp 1698431365
transform 1 0 27552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_292
timestamp 1698431365
transform 1 0 34048 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_378
timestamp 1698431365
transform 1 0 43680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_382
timestamp 1698431365
transform 1 0 44128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_386
timestamp 1698431365
transform 1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_390
timestamp 1698431365
transform 1 0 45024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_426
timestamp 1698431365
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_430
timestamp 1698431365
transform 1 0 49504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_432
timestamp 1698431365
transform 1 0 49728 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_449
timestamp 1698431365
transform 1 0 51632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_453
timestamp 1698431365
transform 1 0 52080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_457
timestamp 1698431365
transform 1 0 52528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_461
timestamp 1698431365
transform 1 0 52976 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_465
timestamp 1698431365
transform 1 0 53424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_467
timestamp 1698431365
transform 1 0 53648 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_480
timestamp 1698431365
transform 1 0 55104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_496
timestamp 1698431365
transform 1 0 56896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_500
timestamp 1698431365
transform 1 0 57344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_504
timestamp 1698431365
transform 1 0 57792 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_509
timestamp 1698431365
transform 1 0 58352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_517
timestamp 1698431365
transform 1 0 59248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_521
timestamp 1698431365
transform 1 0 59696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_525
timestamp 1698431365
transform 1 0 60144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_542
timestamp 1698431365
transform 1 0 62048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_546
timestamp 1698431365
transform 1 0 62496 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_562
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_627
timestamp 1698431365
transform 1 0 71568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_629
timestamp 1698431365
transform 1 0 71792 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_26
timestamp 1698431365
transform 1 0 4256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_78
timestamp 1698431365
transform 1 0 10080 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_165
timestamp 1698431365
transform 1 0 19824 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_187
timestamp 1698431365
transform 1 0 22288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_220
timestamp 1698431365
transform 1 0 25984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_222
timestamp 1698431365
transform 1 0 26208 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_225
timestamp 1698431365
transform 1 0 26544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_260
timestamp 1698431365
transform 1 0 30464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_262
timestamp 1698431365
transform 1 0 30688 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_351
timestamp 1698431365
transform 1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_355
timestamp 1698431365
transform 1 0 41104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_357
timestamp 1698431365
transform 1 0 41328 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_391
timestamp 1698431365
transform 1 0 45136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_393
timestamp 1698431365
transform 1 0 45360 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_412
timestamp 1698431365
transform 1 0 47488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_414
timestamp 1698431365
transform 1 0 47712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_431
timestamp 1698431365
transform 1 0 49616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_435
timestamp 1698431365
transform 1 0 50064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_439
timestamp 1698431365
transform 1 0 50512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_454
timestamp 1698431365
transform 1 0 52192 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_459
timestamp 1698431365
transform 1 0 52752 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_516
timestamp 1698431365
transform 1 0 59136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_531
timestamp 1698431365
transform 1 0 60816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_535
timestamp 1698431365
transform 1 0 61264 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_561
timestamp 1698431365
transform 1 0 64176 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_578
timestamp 1698431365
transform 1 0 66080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_580
timestamp 1698431365
transform 1 0 66304 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_594
timestamp 1698431365
transform 1 0 67872 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_597
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_664
timestamp 1698431365
transform 1 0 75712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_687
timestamp 1698431365
transform 1 0 78288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_48
timestamp 1698431365
transform 1 0 6720 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_137
timestamp 1698431365
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_144
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_197
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_245
timestamp 1698431365
transform 1 0 28784 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_251
timestamp 1698431365
transform 1 0 29456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_255
timestamp 1698431365
transform 1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_259
timestamp 1698431365
transform 1 0 30352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_354
timestamp 1698431365
transform 1 0 40992 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_357
timestamp 1698431365
transform 1 0 41328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_377
timestamp 1698431365
transform 1 0 43568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_381
timestamp 1698431365
transform 1 0 44016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_385
timestamp 1698431365
transform 1 0 44464 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_430
timestamp 1698431365
transform 1 0 49504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_432
timestamp 1698431365
transform 1 0 49728 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_488
timestamp 1698431365
transform 1 0 56000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_528
timestamp 1698431365
transform 1 0 60480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_530
timestamp 1698431365
transform 1 0 60704 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_535
timestamp 1698431365
transform 1 0 61264 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_629
timestamp 1698431365
transform 1 0 71792 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_648
timestamp 1698431365
transform 1 0 73920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_687
timestamp 1698431365
transform 1 0 78288 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_43
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_46
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_50
timestamp 1698431365
transform 1 0 6944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_52
timestamp 1698431365
transform 1 0 7168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_55
timestamp 1698431365
transform 1 0 7504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_65
timestamp 1698431365
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_67
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_109
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_157
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_233
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_361
timestamp 1698431365
transform 1 0 41776 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_394
timestamp 1698431365
transform 1 0 45472 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_420
timestamp 1698431365
transform 1 0 48384 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_443
timestamp 1698431365
transform 1 0 50960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_463
timestamp 1698431365
transform 1 0 53200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_465
timestamp 1698431365
transform 1 0 53424 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_502
timestamp 1698431365
transform 1 0 57568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_522
timestamp 1698431365
transform 1 0 59808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_524
timestamp 1698431365
transform 1 0 60032 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_535
timestamp 1698431365
transform 1 0 61264 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_548
timestamp 1698431365
transform 1 0 62720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_550
timestamp 1698431365
transform 1 0 62944 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_560
timestamp 1698431365
transform 1 0 64064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_594
timestamp 1698431365
transform 1 0 67872 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_687
timestamp 1698431365
transform 1 0 78288 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_50
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_58
timestamp 1698431365
transform 1 0 7840 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_62
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_100
timestamp 1698431365
transform 1 0 12544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_102
timestamp 1698431365
transform 1 0 12768 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_154
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_186
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_214
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_256
timestamp 1698431365
transform 1 0 30016 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_292
timestamp 1698431365
transform 1 0 34048 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_295
timestamp 1698431365
transform 1 0 34384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_315
timestamp 1698431365
transform 1 0 36624 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_325
timestamp 1698431365
transform 1 0 37744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_329
timestamp 1698431365
transform 1 0 38192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_331
timestamp 1698431365
transform 1 0 38416 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_364
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_418
timestamp 1698431365
transform 1 0 48160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_463
timestamp 1698431365
transform 1 0 53200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_467
timestamp 1698431365
transform 1 0 53648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_471
timestamp 1698431365
transform 1 0 54096 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_488
timestamp 1698431365
transform 1 0 56000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_496
timestamp 1698431365
transform 1 0 56896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_500
timestamp 1698431365
transform 1 0 57344 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_512
timestamp 1698431365
transform 1 0 58688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_516
timestamp 1698431365
transform 1 0 59136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_520
timestamp 1698431365
transform 1 0 59584 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_524
timestamp 1698431365
transform 1 0 60032 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_527
timestamp 1698431365
transform 1 0 60368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_529
timestamp 1698431365
transform 1 0 60592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_532
timestamp 1698431365
transform 1 0 60928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_536
timestamp 1698431365
transform 1 0 61376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_544
timestamp 1698431365
transform 1 0 62272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_582
timestamp 1698431365
transform 1 0 66528 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_611
timestamp 1698431365
transform 1 0 69776 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_627
timestamp 1698431365
transform 1 0 71568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_629
timestamp 1698431365
transform 1 0 71792 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_670
timestamp 1698431365
transform 1 0 76384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_672
timestamp 1698431365
transform 1 0 76608 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_685
timestamp 1698431365
transform 1 0 78064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_687
timestamp 1698431365
transform 1 0 78288 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_71
timestamp 1698431365
transform 1 0 9296 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_74
timestamp 1698431365
transform 1 0 9632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_84
timestamp 1698431365
transform 1 0 10752 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_121
timestamp 1698431365
transform 1 0 14896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_153
timestamp 1698431365
transform 1 0 18480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_157
timestamp 1698431365
transform 1 0 18928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_161
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_167
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_206
timestamp 1698431365
transform 1 0 24416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_236
timestamp 1698431365
transform 1 0 27776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_238
timestamp 1698431365
transform 1 0 28000 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_331
timestamp 1698431365
transform 1 0 38416 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_350
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_354
timestamp 1698431365
transform 1 0 40992 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_473
timestamp 1698431365
transform 1 0 54320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_477
timestamp 1698431365
transform 1 0 54768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_481
timestamp 1698431365
transform 1 0 55216 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_513
timestamp 1698431365
transform 1 0 58800 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_524
timestamp 1698431365
transform 1 0 60032 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_533
timestamp 1698431365
transform 1 0 61040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_537
timestamp 1698431365
transform 1 0 61488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_547
timestamp 1698431365
transform 1 0 62608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_557
timestamp 1698431365
transform 1 0 63728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_559
timestamp 1698431365
transform 1 0 63952 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_562
timestamp 1698431365
transform 1 0 64288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_564
timestamp 1698431365
transform 1 0 64512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_567
timestamp 1698431365
transform 1 0 64848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_569
timestamp 1698431365
transform 1 0 65072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_576
timestamp 1698431365
transform 1 0 65856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_580
timestamp 1698431365
transform 1 0 66304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_582
timestamp 1698431365
transform 1 0 66528 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_611
timestamp 1698431365
transform 1 0 69776 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_655
timestamp 1698431365
transform 1 0 74704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_659
timestamp 1698431365
transform 1 0 75152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_663
timestamp 1698431365
transform 1 0 75600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_671
timestamp 1698431365
transform 1 0 76496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_679
timestamp 1698431365
transform 1 0 77392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_681
timestamp 1698431365
transform 1 0 77616 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_101
timestamp 1698431365
transform 1 0 12656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_105
timestamp 1698431365
transform 1 0 13104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_109
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_115
timestamp 1698431365
transform 1 0 14224 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_121
timestamp 1698431365
transform 1 0 14896 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_124
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_132
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_150
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_154
timestamp 1698431365
transform 1 0 18592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_156
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_222
timestamp 1698431365
transform 1 0 26208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_226
timestamp 1698431365
transform 1 0 26656 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_229
timestamp 1698431365
transform 1 0 26992 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_233
timestamp 1698431365
transform 1 0 27440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_288
timestamp 1698431365
transform 1 0 33600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_313
timestamp 1698431365
transform 1 0 36400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_317
timestamp 1698431365
transform 1 0 36848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_319
timestamp 1698431365
transform 1 0 37072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_430
timestamp 1698431365
transform 1 0 49504 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_455
timestamp 1698431365
transform 1 0 52304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_459
timestamp 1698431365
transform 1 0 52752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_463
timestamp 1698431365
transform 1 0 53200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_467
timestamp 1698431365
transform 1 0 53648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_471
timestamp 1698431365
transform 1 0 54096 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_487
timestamp 1698431365
transform 1 0 55888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_489
timestamp 1698431365
transform 1 0 56112 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_524
timestamp 1698431365
transform 1 0 60032 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_540
timestamp 1698431365
transform 1 0 61824 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_548
timestamp 1698431365
transform 1 0 62720 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_552
timestamp 1698431365
transform 1 0 63168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_566
timestamp 1698431365
transform 1 0 64736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_570
timestamp 1698431365
transform 1 0 65184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_574
timestamp 1698431365
transform 1 0 65632 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_580
timestamp 1698431365
transform 1 0 66304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_584
timestamp 1698431365
transform 1 0 66752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_587
timestamp 1698431365
transform 1 0 67088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_593
timestamp 1698431365
transform 1 0 67760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_597
timestamp 1698431365
transform 1 0 68208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_603
timestamp 1698431365
transform 1 0 68880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_607
timestamp 1698431365
transform 1 0 69328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_609
timestamp 1698431365
transform 1 0 69552 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_612
timestamp 1698431365
transform 1 0 69888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_628
timestamp 1698431365
transform 1 0 71680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_636
timestamp 1698431365
transform 1 0 72576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_640
timestamp 1698431365
transform 1 0 73024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_644
timestamp 1698431365
transform 1 0 73472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_648
timestamp 1698431365
transform 1 0 73920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_652
timestamp 1698431365
transform 1 0 74368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_656
timestamp 1698431365
transform 1 0 74816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_660
timestamp 1698431365
transform 1 0 75264 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_664
timestamp 1698431365
transform 1 0 75712 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_667
timestamp 1698431365
transform 1 0 76048 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_673
timestamp 1698431365
transform 1 0 76720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_677
timestamp 1698431365
transform 1 0 77168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_679
timestamp 1698431365
transform 1 0 77392 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_85
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_99
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_127
timestamp 1698431365
transform 1 0 15568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_131
timestamp 1698431365
transform 1 0 16016 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_139
timestamp 1698431365
transform 1 0 16912 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_143
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_147
timestamp 1698431365
transform 1 0 17808 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_153
timestamp 1698431365
transform 1 0 18480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_159
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_188
timestamp 1698431365
transform 1 0 22400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_192
timestamp 1698431365
transform 1 0 22848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_225
timestamp 1698431365
transform 1 0 26544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_229
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_233
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_237
timestamp 1698431365
transform 1 0 27888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_331
timestamp 1698431365
transform 1 0 38416 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_396
timestamp 1698431365
transform 1 0 45696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_429
timestamp 1698431365
transform 1 0 49392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_433
timestamp 1698431365
transform 1 0 49840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_437
timestamp 1698431365
transform 1 0 50288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_454
timestamp 1698431365
transform 1 0 52192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698431365
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_601
timestamp 1698431365
transform 1 0 68656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_605
timestamp 1698431365
transform 1 0 69104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_609
timestamp 1698431365
transform 1 0 69552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_613
timestamp 1698431365
transform 1 0 70000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_617
timestamp 1698431365
transform 1 0 70448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_621
timestamp 1698431365
transform 1 0 70896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_625
timestamp 1698431365
transform 1 0 71344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_629
timestamp 1698431365
transform 1 0 71792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_633
timestamp 1698431365
transform 1 0 72240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_637
timestamp 1698431365
transform 1 0 72688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_641
timestamp 1698431365
transform 1 0 73136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_645
timestamp 1698431365
transform 1 0 73584 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_648
timestamp 1698431365
transform 1 0 73920 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_664
timestamp 1698431365
transform 1 0 75712 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_667
timestamp 1698431365
transform 1 0 76048 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_683
timestamp 1698431365
transform 1 0 77840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_687
timestamp 1698431365
transform 1 0 78288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_86
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_137
timestamp 1698431365
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_148
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_182
timestamp 1698431365
transform 1 0 21728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_184
timestamp 1698431365
transform 1 0 21952 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_187
timestamp 1698431365
transform 1 0 22288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_191
timestamp 1698431365
transform 1 0 22736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_228
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_233
timestamp 1698431365
transform 1 0 27440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_235
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_242
timestamp 1698431365
transform 1 0 28448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_246
timestamp 1698431365
transform 1 0 28896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_264
timestamp 1698431365
transform 1 0 30912 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_270
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_339
timestamp 1698431365
transform 1 0 39312 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_358
timestamp 1698431365
transform 1 0 41440 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_390
timestamp 1698431365
transform 1 0 45024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_392
timestamp 1698431365
transform 1 0 45248 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_426
timestamp 1698431365
transform 1 0 49056 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_431
timestamp 1698431365
transform 1 0 49616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_435
timestamp 1698431365
transform 1 0 50064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_439
timestamp 1698431365
transform 1 0 50512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_443
timestamp 1698431365
transform 1 0 50960 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_475
timestamp 1698431365
transform 1 0 54544 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_483
timestamp 1698431365
transform 1 0 55440 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_487
timestamp 1698431365
transform 1 0 55888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_489
timestamp 1698431365
transform 1 0 56112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_664
timestamp 1698431365
transform 1 0 75712 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_680
timestamp 1698431365
transform 1 0 77504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_73
timestamp 1698431365
transform 1 0 9520 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_75
timestamp 1698431365
transform 1 0 9744 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_145
timestamp 1698431365
transform 1 0 17584 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_153
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_165
timestamp 1698431365
transform 1 0 19824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_183
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_197
timestamp 1698431365
transform 1 0 23408 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_200
timestamp 1698431365
transform 1 0 23744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_204
timestamp 1698431365
transform 1 0 24192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_208
timestamp 1698431365
transform 1 0 24640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_212
timestamp 1698431365
transform 1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_216
timestamp 1698431365
transform 1 0 25536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_220
timestamp 1698431365
transform 1 0 25984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_224
timestamp 1698431365
transform 1 0 26432 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_235
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_259
timestamp 1698431365
transform 1 0 30352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_262
timestamp 1698431365
transform 1 0 30688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_266
timestamp 1698431365
transform 1 0 31136 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_280
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_354
timestamp 1698431365
transform 1 0 40992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_360
timestamp 1698431365
transform 1 0 41664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_364
timestamp 1698431365
transform 1 0 42112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_368
timestamp 1698431365
transform 1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_372
timestamp 1698431365
transform 1 0 43008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_380
timestamp 1698431365
transform 1 0 43904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_389
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_392
timestamp 1698431365
transform 1 0 45248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_396
timestamp 1698431365
transform 1 0 45696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_398
timestamp 1698431365
transform 1 0 45920 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_415
timestamp 1698431365
transform 1 0 47824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_419
timestamp 1698431365
transform 1 0 48272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_423
timestamp 1698431365
transform 1 0 48720 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698431365
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698431365
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_667
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_683
timestamp 1698431365
transform 1 0 77840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_687
timestamp 1698431365
transform 1 0 78288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_107
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_260
timestamp 1698431365
transform 1 0 30464 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_268
timestamp 1698431365
transform 1 0 31360 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_272
timestamp 1698431365
transform 1 0 31808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_316
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_332
timestamp 1698431365
transform 1 0 38528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698431365
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_632
timestamp 1698431365
transform 1 0 72128 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_664
timestamp 1698431365
transform 1 0 75712 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_680
timestamp 1698431365
transform 1 0 77504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_279
timestamp 1698431365
transform 1 0 32592 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_303
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_323
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_330
timestamp 1698431365
transform 1 0 38304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_334
timestamp 1698431365
transform 1 0 38752 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_366
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_382
timestamp 1698431365
transform 1 0 44128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698431365
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698431365
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698431365
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_683
timestamp 1698431365
transform 1 0 77840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_687
timestamp 1698431365
transform 1 0 78288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_294
timestamp 1698431365
transform 1 0 34272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_296
timestamp 1698431365
transform 1 0 34496 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_313
timestamp 1698431365
transform 1 0 36400 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_664
timestamp 1698431365
transform 1 0 75712 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_680
timestamp 1698431365
transform 1 0 77504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698431365
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698431365
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698431365
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_683
timestamp 1698431365
transform 1 0 77840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_687
timestamp 1698431365
transform 1 0 78288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698431365
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_664
timestamp 1698431365
transform 1 0 75712 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_680
timestamp 1698431365
transform 1 0 77504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698431365
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698431365
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_683
timestamp 1698431365
transform 1 0 77840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_687
timestamp 1698431365
transform 1 0 78288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_632
timestamp 1698431365
transform 1 0 72128 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_664
timestamp 1698431365
transform 1 0 75712 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_680
timestamp 1698431365
transform 1 0 77504 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698431365
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_661
timestamp 1698431365
transform 1 0 75376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_667
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_683
timestamp 1698431365
transform 1 0 77840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_687
timestamp 1698431365
transform 1 0 78288 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698431365
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_664
timestamp 1698431365
transform 1 0 75712 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_680
timestamp 1698431365
transform 1 0 77504 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_521
timestamp 1698431365
transform 1 0 59696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698431365
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_661
timestamp 1698431365
transform 1 0 75376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_683
timestamp 1698431365
transform 1 0 77840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_687
timestamp 1698431365
transform 1 0 78288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698431365
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_626
timestamp 1698431365
transform 1 0 71456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_632
timestamp 1698431365
transform 1 0 72128 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_664
timestamp 1698431365
transform 1 0 75712 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_680
timestamp 1698431365
transform 1 0 77504 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_521
timestamp 1698431365
transform 1 0 59696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698431365
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_597
timestamp 1698431365
transform 1 0 68208 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_661
timestamp 1698431365
transform 1 0 75376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_667
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_683
timestamp 1698431365
transform 1 0 77840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_687
timestamp 1698431365
transform 1 0 78288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698431365
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_626
timestamp 1698431365
transform 1 0 71456 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_632
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_664
timestamp 1698431365
transform 1 0 75712 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_680
timestamp 1698431365
transform 1 0 77504 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698431365
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_661
timestamp 1698431365
transform 1 0 75376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_667
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_683
timestamp 1698431365
transform 1 0 77840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_687
timestamp 1698431365
transform 1 0 78288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_556
timestamp 1698431365
transform 1 0 63616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_632
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_664
timestamp 1698431365
transform 1 0 75712 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_680
timestamp 1698431365
transform 1 0 77504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698431365
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698431365
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_661
timestamp 1698431365
transform 1 0 75376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_667
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_683
timestamp 1698431365
transform 1 0 77840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_687
timestamp 1698431365
transform 1 0 78288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698431365
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_626
timestamp 1698431365
transform 1 0 71456 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_632
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_664
timestamp 1698431365
transform 1 0 75712 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_680
timestamp 1698431365
transform 1 0 77504 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698431365
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698431365
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_661
timestamp 1698431365
transform 1 0 75376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_667
timestamp 1698431365
transform 1 0 76048 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_683
timestamp 1698431365
transform 1 0 77840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_687
timestamp 1698431365
transform 1 0 78288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698431365
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_626
timestamp 1698431365
transform 1 0 71456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_632
timestamp 1698431365
transform 1 0 72128 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_664
timestamp 1698431365
transform 1 0 75712 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_680
timestamp 1698431365
transform 1 0 77504 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698431365
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_661
timestamp 1698431365
transform 1 0 75376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_667
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_683
timestamp 1698431365
transform 1 0 77840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_687
timestamp 1698431365
transform 1 0 78288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698431365
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_626
timestamp 1698431365
transform 1 0 71456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_632
timestamp 1698431365
transform 1 0 72128 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_664
timestamp 1698431365
transform 1 0 75712 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_680
timestamp 1698431365
transform 1 0 77504 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_521
timestamp 1698431365
transform 1 0 59696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_661
timestamp 1698431365
transform 1 0 75376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_667
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_683
timestamp 1698431365
transform 1 0 77840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_687
timestamp 1698431365
transform 1 0 78288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698431365
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_632
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_664
timestamp 1698431365
transform 1 0 75712 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_680
timestamp 1698431365
transform 1 0 77504 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_521
timestamp 1698431365
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_661
timestamp 1698431365
transform 1 0 75376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_667
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_683
timestamp 1698431365
transform 1 0 77840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_687
timestamp 1698431365
transform 1 0 78288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_626
timestamp 1698431365
transform 1 0 71456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_632
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_664
timestamp 1698431365
transform 1 0 75712 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_680
timestamp 1698431365
transform 1 0 77504 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698431365
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698431365
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698431365
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_683
timestamp 1698431365
transform 1 0 77840 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_687
timestamp 1698431365
transform 1 0 78288 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_626
timestamp 1698431365
transform 1 0 71456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_632
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_664
timestamp 1698431365
transform 1 0 75712 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_680
timestamp 1698431365
transform 1 0 77504 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_521
timestamp 1698431365
transform 1 0 59696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_661
timestamp 1698431365
transform 1 0 75376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_667
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_683
timestamp 1698431365
transform 1 0 77840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_687
timestamp 1698431365
transform 1 0 78288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698431365
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_632
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_664
timestamp 1698431365
transform 1 0 75712 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_680
timestamp 1698431365
transform 1 0 77504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_36
timestamp 1698431365
transform 1 0 5376 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_138
timestamp 1698431365
transform 1 0 16800 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_206
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_274
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_342
timestamp 1698431365
transform 1 0 39648 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_376
timestamp 1698431365
transform 1 0 43456 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_410
timestamp 1698431365
transform 1 0 47264 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_444
timestamp 1698431365
transform 1 0 51072 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_478
timestamp 1698431365
transform 1 0 54880 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_512
timestamp 1698431365
transform 1 0 58688 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_546
timestamp 1698431365
transform 1 0 62496 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_580
timestamp 1698431365
transform 1 0 66304 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_614
timestamp 1698431365
transform 1 0 70112 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_648
timestamp 1698431365
transform 1 0 73920 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_682
timestamp 1698431365
transform 1 0 77728 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_686
timestamp 1698431365
transform 1 0 78176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 71792 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 62048 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 47488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 47488 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform -1 0 75376 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform -1 0 62048 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold7
timestamp 1698431365
transform -1 0 47040 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold8
timestamp 1698431365
transform -1 0 47824 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold9
timestamp 1698431365
transform 1 0 68320 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold10
timestamp 1698431365
transform -1 0 59248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold11
timestamp 1698431365
transform -1 0 46368 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold12
timestamp 1698431365
transform -1 0 43680 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold13
timestamp 1698431365
transform -1 0 77840 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold14
timestamp 1698431365
transform -1 0 63168 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold15
timestamp 1698431365
transform 1 0 50512 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold16
timestamp 1698431365
transform -1 0 55328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold17
timestamp 1698431365
transform 1 0 73920 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold18
timestamp 1698431365
transform -1 0 63168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold19
timestamp 1698431365
transform -1 0 51632 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold20
timestamp 1698431365
transform -1 0 56000 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold21
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold22
timestamp 1698431365
transform -1 0 63168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold23
timestamp 1698431365
transform -1 0 50288 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold24
timestamp 1698431365
transform -1 0 51408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold25
timestamp 1698431365
transform -1 0 75600 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold26
timestamp 1698431365
transform -1 0 65968 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold27
timestamp 1698431365
transform 1 0 47824 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold28
timestamp 1698431365
transform -1 0 52192 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold29
timestamp 1698431365
transform 1 0 67088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold30
timestamp 1698431365
transform -1 0 59024 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold31
timestamp 1698431365
transform -1 0 43568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold32
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold33
timestamp 1698431365
transform -1 0 67760 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold34
timestamp 1698431365
transform -1 0 48384 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold35
timestamp 1698431365
transform -1 0 29792 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold36
timestamp 1698431365
transform 1 0 26992 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold37
timestamp 1698431365
transform -1 0 71680 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold38
timestamp 1698431365
transform -1 0 50064 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold39
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold40
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold41
timestamp 1698431365
transform -1 0 73920 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold42
timestamp 1698431365
transform -1 0 56224 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold43
timestamp 1698431365
transform -1 0 40544 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold44
timestamp 1698431365
transform -1 0 39200 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold45
timestamp 1698431365
transform -1 0 70672 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold46
timestamp 1698431365
transform -1 0 58464 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold47
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold48
timestamp 1698431365
transform 1 0 34944 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold49
timestamp 1698431365
transform 1 0 62272 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  hold50
timestamp 1698431365
transform -1 0 48496 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold51
timestamp 1698431365
transform -1 0 32592 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold52
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold53
timestamp 1698431365
transform 1 0 64288 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold54
timestamp 1698431365
transform -1 0 51408 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold55
timestamp 1698431365
transform -1 0 29792 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold56
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold57
timestamp 1698431365
transform -1 0 70000 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold58
timestamp 1698431365
transform -1 0 54432 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold59
timestamp 1698431365
transform -1 0 36400 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold60
timestamp 1698431365
transform 1 0 33488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold61
timestamp 1698431365
transform -1 0 71792 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold62
timestamp 1698431365
transform -1 0 55664 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold63
timestamp 1698431365
transform -1 0 36400 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold64
timestamp 1698431365
transform -1 0 36624 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold65
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold66
timestamp 1698431365
transform -1 0 77840 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  hold67
timestamp 1698431365
transform -1 0 59248 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold68
timestamp 1698431365
transform 1 0 74144 0 -1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold69
timestamp 1698431365
transform 1 0 68096 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold70
timestamp 1698431365
transform 1 0 41664 0 1 9408
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold71
timestamp 1698431365
transform -1 0 74928 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold72
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold73
timestamp 1698431365
transform 1 0 45360 0 -1 12544
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold74
timestamp 1698431365
transform -1 0 73808 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold75
timestamp 1698431365
transform 1 0 74928 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold76
timestamp 1698431365
transform 1 0 70112 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold77
timestamp 1698431365
transform 1 0 72912 0 1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold78
timestamp 1698431365
transform 1 0 45584 0 1 7840
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold79
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold80
timestamp 1698431365
transform 1 0 70112 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold81
timestamp 1698431365
transform 1 0 62608 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold82
timestamp 1698431365
transform 1 0 74928 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold83
timestamp 1698431365
transform 1 0 64848 0 -1 6272
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold84
timestamp 1698431365
transform -1 0 69104 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold85
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold86
timestamp 1698431365
transform 1 0 67088 0 -1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold87
timestamp 1698431365
transform -1 0 76720 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 66080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 64064 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 65856 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 65184 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 67200 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 68432 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 67312 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 69776 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 67984 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 77392 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 72240 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 78400 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 74256 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 71232 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 78400 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 78400 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 77392 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 78064 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 69776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 63392 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 65856 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 66528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698431365
transform -1 0 66528 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 67872 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform -1 0 73696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 71344 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 77392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 69104 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 71568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 72912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 78400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input32
timestamp 1698431365
transform -1 0 73584 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 78288 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 77616 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 78400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 76384 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input37
timestamp 1698431365
transform 1 0 4368 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input38
timestamp 1698431365
transform 1 0 3360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 4592 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input40
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input41
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 19040 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input43
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input45
timestamp 1698431365
transform 1 0 18480 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 6832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 9520 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 9520 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform 1 0 10192 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 2688 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform 1 0 13104 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 22064 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 2016 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform 1 0 2016 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input57
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29792 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform -1 0 39984 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform -1 0 40544 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698431365
transform -1 0 42000 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698431365
transform -1 0 43680 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698431365
transform 1 0 30800 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698431365
transform 1 0 28896 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698431365
transform 1 0 29792 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698431365
transform 1 0 30800 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output70
timestamp 1698431365
transform -1 0 36624 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output71
timestamp 1698431365
transform -1 0 37072 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output72
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output73
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output74
timestamp 1698431365
transform 1 0 34720 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output75
timestamp 1698431365
transform -1 0 6272 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output76
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output77
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output78
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output79
timestamp 1698431365
transform -1 0 20160 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output80
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output81
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output82
timestamp 1698431365
transform -1 0 22064 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform -1 0 6272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform -1 0 13776 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform -1 0 16688 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_106
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_107
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_108
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_109
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_110
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_115
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_121
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_122
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_123
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_124
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_126
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_127
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_128
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_129
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_130
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_131
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_134
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_135
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_136
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_137
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_149
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_150
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_151
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_152
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_155
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_156
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_157
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_158
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_160
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_161
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_162
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_163
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_164
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_165
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_170
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_171
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_174
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_175
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_176
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_177
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_178
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_179
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_180
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_181
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_182
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_183
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_184
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_185
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_186
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_187
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_188
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_189
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_190
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_191
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_192
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_193
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_194
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_195
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_196
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_197
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_198
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_199
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_200
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_201
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_202
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_203
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_204
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_205
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_206
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_207
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_208
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_209
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_210
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_211
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_212
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_213
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_214
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_215
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_216
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_217
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_218
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_219
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_220
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_221
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_222
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_223
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_224
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_225
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_226
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_227
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_228
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_229
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_230
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_231
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_232
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_233
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_234
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_235
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_236
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_237
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_238
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_239
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_240
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_241
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_242
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_243
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_244
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_245
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_246
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_247
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_248
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_249
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_250
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_251
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_252
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_253
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_254
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_258
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_259
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_260
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_261
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_267
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_268
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_276
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_283
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_284
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_285
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_290
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_291
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_292
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_293
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_294
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_295
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_297
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_298
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_299
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_300
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_301
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_302
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_303
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_304
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_305
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_306
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_307
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_308
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_309
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_310
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_311
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_312
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_313
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_314
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_315
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_316
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_317
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_318
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_319
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_320
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_321
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_322
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_323
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_324
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_325
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_326
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_327
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_328
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_329
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_330
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_331
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_332
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_333
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_334
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_335
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_336
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_337
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_338
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_339
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_340
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_341
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_342
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_343
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_344
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_345
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_346
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_347
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_348
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_349
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_350
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_351
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_352
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_353
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_354
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_355
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_356
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_357
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_358
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_359
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_360
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_361
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_362
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_363
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_364
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_365
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_366
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_367
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_371
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_372
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_377
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_378
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_379
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_380
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_382
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_383
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_384
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_385
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_386
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_387
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_388
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_389
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_390
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_391
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_392
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_393
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_394
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_395
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_396
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_397
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_398
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_399
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_400
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_401
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_402
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_403
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_404
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_405
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_406
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_407
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_408
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_409
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_410
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_411
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_412
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_413
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_414
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_415
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_416
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_417
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_418
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_419
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_420
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_421
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_422
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_423
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_424
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_425
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_426
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_427
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_428
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_429
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_430
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_431
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_432
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_433
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_434
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_435
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_436
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_437
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_438
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_439
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_440
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_441
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_442
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_443
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_444
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_445
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_446
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_447
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_448
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_449
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_450
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_451
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_452
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_453
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_454
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_455
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_456
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_457
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_458
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_459
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_460
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_461
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_462
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_463
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_464
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_465
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_466
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_467
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_468
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_469
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_470
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_471
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_472
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_473
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_474
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_475
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_476
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_477
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_478
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_479
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_480
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_481
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_482
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_483
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_484
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_485
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_486
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_487
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_488
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_489
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_490
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_491
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_492
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_493
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_494
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_495
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_496
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_497
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_498
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_499
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_500
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_501
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_502
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_503
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_504
timestamp 1698431365
transform 1 0 39424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_505
timestamp 1698431365
transform 1 0 43232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_506
timestamp 1698431365
transform 1 0 47040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_507
timestamp 1698431365
transform 1 0 50848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_508
timestamp 1698431365
transform 1 0 54656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_509
timestamp 1698431365
transform 1 0 58464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_510
timestamp 1698431365
transform 1 0 62272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_511
timestamp 1698431365
transform 1 0 66080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_512
timestamp 1698431365
transform 1 0 69888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_513
timestamp 1698431365
transform 1 0 73696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_514
timestamp 1698431365
transform 1 0 77504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_95 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_96
timestamp 1698431365
transform -1 0 52304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_97
timestamp 1698431365
transform -1 0 52976 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_98
timestamp 1698431365
transform -1 0 49616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_99
timestamp 1698431365
transform -1 0 51856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_100
timestamp 1698431365
transform -1 0 53424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_101
timestamp 1698431365
transform -1 0 52304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_102
timestamp 1698431365
transform -1 0 53872 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_103
timestamp 1698431365
transform -1 0 54320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_104
timestamp 1698431365
transform -1 0 55776 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_105
timestamp 1698431365
transform -1 0 56224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_106
timestamp 1698431365
transform -1 0 56672 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_107
timestamp 1698431365
transform -1 0 57120 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_108
timestamp 1698431365
transform -1 0 62272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_109
timestamp 1698431365
transform -1 0 57568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_110
timestamp 1698431365
transform -1 0 60032 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_111
timestamp 1698431365
transform -1 0 59360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_112
timestamp 1698431365
transform -1 0 60480 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_113
timestamp 1698431365
transform -1 0 59808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_114
timestamp 1698431365
transform -1 0 61264 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_115
timestamp 1698431365
transform -1 0 62272 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_116
timestamp 1698431365
transform 1 0 60816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_117
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_118
timestamp 1698431365
transform -1 0 68096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_119
timestamp 1698431365
transform -1 0 63728 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_120
timestamp 1698431365
transform -1 0 64848 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_121
timestamp 1698431365
transform -1 0 65632 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_122
timestamp 1698431365
transform -1 0 71792 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_123
timestamp 1698431365
transform -1 0 67760 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_124
timestamp 1698431365
transform -1 0 67312 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_125
timestamp 1698431365
transform -1 0 68880 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_126
timestamp 1698431365
transform -1 0 69328 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_127
timestamp 1698431365
transform -1 0 69776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_128
timestamp 1698431365
transform -1 0 70560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_129
timestamp 1698431365
transform -1 0 75824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_130
timestamp 1698431365
transform -1 0 71680 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_131
timestamp 1698431365
transform -1 0 72576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_132
timestamp 1698431365
transform -1 0 78288 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_133
timestamp 1698431365
transform -1 0 74704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_134
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_135
timestamp 1698431365
transform -1 0 22400 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_136
timestamp 1698431365
transform -1 0 23968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_137
timestamp 1698431365
transform -1 0 23296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_138
timestamp 1698431365
transform -1 0 22848 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_139
timestamp 1698431365
transform -1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_140
timestamp 1698431365
transform 1 0 22400 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_141
timestamp 1698431365
transform -1 0 26208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_142
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_143
timestamp 1698431365
transform 1 0 24640 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_144
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_145
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_146
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_147
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_148
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_149
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_150
timestamp 1698431365
transform -1 0 78288 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_151
timestamp 1698431365
transform -1 0 76496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_152
timestamp 1698431365
transform -1 0 78288 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_153
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_154
timestamp 1698431365
transform -1 0 45696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_155
timestamp 1698431365
transform -1 0 56112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_156
timestamp 1698431365
transform -1 0 51408 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_157
timestamp 1698431365
transform -1 0 49728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_158
timestamp 1698431365
transform -1 0 49056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_159
timestamp 1698431365
transform -1 0 58352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_160
timestamp 1698431365
transform -1 0 53760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_161
timestamp 1698431365
transform -1 0 54208 0 -1 7840
box -86 -86 534 870
<< labels >>
flabel metal2 s 73024 0 73136 800 0 FreeSans 448 90 0 0 irq[0]
port 0 nsew signal tristate
flabel metal2 s 73248 0 73360 800 0 FreeSans 448 90 0 0 irq[1]
port 1 nsew signal tristate
flabel metal2 s 73472 0 73584 800 0 FreeSans 448 90 0 0 irq[2]
port 2 nsew signal tristate
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 3 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 4 nsew signal input
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 5 nsew signal input
flabel metal2 s 38080 0 38192 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 6 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 7 nsew signal input
flabel metal2 s 39424 0 39536 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 8 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 9 nsew signal input
flabel metal2 s 40768 0 40880 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 10 nsew signal input
flabel metal2 s 41440 0 41552 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 11 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 12 nsew signal input
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 13 nsew signal input
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 14 nsew signal input
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 15 nsew signal input
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 16 nsew signal input
flabel metal2 s 44800 0 44912 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 17 nsew signal input
flabel metal2 s 45472 0 45584 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 18 nsew signal input
flabel metal2 s 46144 0 46256 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 19 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 20 nsew signal input
flabel metal2 s 47488 0 47600 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 21 nsew signal input
flabel metal2 s 48160 0 48272 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 22 nsew signal input
flabel metal2 s 48832 0 48944 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 23 nsew signal input
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 24 nsew signal input
flabel metal2 s 31360 0 31472 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 25 nsew signal input
flabel metal2 s 50176 0 50288 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 26 nsew signal input
flabel metal2 s 50848 0 50960 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 27 nsew signal input
flabel metal2 s 51520 0 51632 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 28 nsew signal input
flabel metal2 s 52192 0 52304 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 29 nsew signal input
flabel metal2 s 52864 0 52976 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 30 nsew signal input
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 31 nsew signal input
flabel metal2 s 54208 0 54320 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 32 nsew signal input
flabel metal2 s 54880 0 54992 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 33 nsew signal input
flabel metal2 s 55552 0 55664 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 34 nsew signal input
flabel metal2 s 56224 0 56336 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 35 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 36 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 37 nsew signal input
flabel metal2 s 57568 0 57680 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 38 nsew signal input
flabel metal2 s 58240 0 58352 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 39 nsew signal input
flabel metal2 s 58912 0 59024 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 40 nsew signal input
flabel metal2 s 59584 0 59696 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 41 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 42 nsew signal input
flabel metal2 s 60928 0 61040 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 43 nsew signal input
flabel metal2 s 61600 0 61712 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 44 nsew signal input
flabel metal2 s 62272 0 62384 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 45 nsew signal input
flabel metal2 s 62944 0 63056 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 46 nsew signal input
flabel metal2 s 32704 0 32816 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 47 nsew signal input
flabel metal2 s 63616 0 63728 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 48 nsew signal input
flabel metal2 s 64288 0 64400 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 49 nsew signal input
flabel metal2 s 64960 0 65072 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 50 nsew signal input
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 51 nsew signal input
flabel metal2 s 66304 0 66416 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 52 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 53 nsew signal input
flabel metal2 s 67648 0 67760 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 54 nsew signal input
flabel metal2 s 68320 0 68432 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 55 nsew signal input
flabel metal2 s 68992 0 69104 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 56 nsew signal input
flabel metal2 s 69664 0 69776 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 57 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 58 nsew signal input
flabel metal2 s 70336 0 70448 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 59 nsew signal input
flabel metal2 s 71008 0 71120 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 60 nsew signal input
flabel metal2 s 71680 0 71792 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 61 nsew signal input
flabel metal2 s 72352 0 72464 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 62 nsew signal input
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 63 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 64 nsew signal input
flabel metal2 s 35392 0 35504 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 65 nsew signal input
flabel metal2 s 36064 0 36176 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 66 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 la_data_out[0]
port 67 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 la_data_out[10]
port 68 nsew signal tristate
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 la_data_out[11]
port 69 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 la_data_out[12]
port 70 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 71 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 la_data_out[14]
port 72 nsew signal tristate
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 la_data_out[15]
port 73 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 la_data_out[16]
port 74 nsew signal tristate
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 75 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 76 nsew signal tristate
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 77 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 la_data_out[1]
port 78 nsew signal tristate
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 la_data_out[20]
port 79 nsew signal tristate
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 la_data_out[21]
port 80 nsew signal tristate
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 la_data_out[22]
port 81 nsew signal tristate
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 82 nsew signal tristate
flabel metal2 s 46368 0 46480 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 83 nsew signal tristate
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 84 nsew signal tristate
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 la_data_out[26]
port 85 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 la_data_out[27]
port 86 nsew signal tristate
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 la_data_out[28]
port 87 nsew signal tristate
flabel metal2 s 49728 0 49840 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 88 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 la_data_out[2]
port 89 nsew signal tristate
flabel metal2 s 50400 0 50512 800 0 FreeSans 448 90 0 0 la_data_out[30]
port 90 nsew signal tristate
flabel metal2 s 51072 0 51184 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 91 nsew signal tristate
flabel metal2 s 51744 0 51856 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 92 nsew signal tristate
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 93 nsew signal tristate
flabel metal2 s 53088 0 53200 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 94 nsew signal tristate
flabel metal2 s 53760 0 53872 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 95 nsew signal tristate
flabel metal2 s 54432 0 54544 800 0 FreeSans 448 90 0 0 la_data_out[36]
port 96 nsew signal tristate
flabel metal2 s 55104 0 55216 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 97 nsew signal tristate
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 la_data_out[38]
port 98 nsew signal tristate
flabel metal2 s 56448 0 56560 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 99 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 la_data_out[3]
port 100 nsew signal tristate
flabel metal2 s 57120 0 57232 800 0 FreeSans 448 90 0 0 la_data_out[40]
port 101 nsew signal tristate
flabel metal2 s 57792 0 57904 800 0 FreeSans 448 90 0 0 la_data_out[41]
port 102 nsew signal tristate
flabel metal2 s 58464 0 58576 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 103 nsew signal tristate
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 104 nsew signal tristate
flabel metal2 s 59808 0 59920 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 105 nsew signal tristate
flabel metal2 s 60480 0 60592 800 0 FreeSans 448 90 0 0 la_data_out[45]
port 106 nsew signal tristate
flabel metal2 s 61152 0 61264 800 0 FreeSans 448 90 0 0 la_data_out[46]
port 107 nsew signal tristate
flabel metal2 s 61824 0 61936 800 0 FreeSans 448 90 0 0 la_data_out[47]
port 108 nsew signal tristate
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 109 nsew signal tristate
flabel metal2 s 63168 0 63280 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 110 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 la_data_out[4]
port 111 nsew signal tristate
flabel metal2 s 63840 0 63952 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 112 nsew signal tristate
flabel metal2 s 64512 0 64624 800 0 FreeSans 448 90 0 0 la_data_out[51]
port 113 nsew signal tristate
flabel metal2 s 65184 0 65296 800 0 FreeSans 448 90 0 0 la_data_out[52]
port 114 nsew signal tristate
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_out[53]
port 115 nsew signal tristate
flabel metal2 s 66528 0 66640 800 0 FreeSans 448 90 0 0 la_data_out[54]
port 116 nsew signal tristate
flabel metal2 s 67200 0 67312 800 0 FreeSans 448 90 0 0 la_data_out[55]
port 117 nsew signal tristate
flabel metal2 s 67872 0 67984 800 0 FreeSans 448 90 0 0 la_data_out[56]
port 118 nsew signal tristate
flabel metal2 s 68544 0 68656 800 0 FreeSans 448 90 0 0 la_data_out[57]
port 119 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_out[58]
port 120 nsew signal tristate
flabel metal2 s 69888 0 70000 800 0 FreeSans 448 90 0 0 la_data_out[59]
port 121 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 la_data_out[5]
port 122 nsew signal tristate
flabel metal2 s 70560 0 70672 800 0 FreeSans 448 90 0 0 la_data_out[60]
port 123 nsew signal tristate
flabel metal2 s 71232 0 71344 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 124 nsew signal tristate
flabel metal2 s 71904 0 72016 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 125 nsew signal tristate
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_out[63]
port 126 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 la_data_out[6]
port 127 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 la_data_out[7]
port 128 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 la_data_out[8]
port 129 nsew signal tristate
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 la_data_out[9]
port 130 nsew signal tristate
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 131 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 la_oenb[10]
port 132 nsew signal input
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 la_oenb[11]
port 133 nsew signal input
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 la_oenb[12]
port 134 nsew signal input
flabel metal2 s 39200 0 39312 800 0 FreeSans 448 90 0 0 la_oenb[13]
port 135 nsew signal input
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 136 nsew signal input
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 137 nsew signal input
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 138 nsew signal input
flabel metal2 s 41888 0 42000 800 0 FreeSans 448 90 0 0 la_oenb[17]
port 139 nsew signal input
flabel metal2 s 42560 0 42672 800 0 FreeSans 448 90 0 0 la_oenb[18]
port 140 nsew signal input
flabel metal2 s 43232 0 43344 800 0 FreeSans 448 90 0 0 la_oenb[19]
port 141 nsew signal input
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 142 nsew signal input
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 la_oenb[20]
port 143 nsew signal input
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 la_oenb[21]
port 144 nsew signal input
flabel metal2 s 45248 0 45360 800 0 FreeSans 448 90 0 0 la_oenb[22]
port 145 nsew signal input
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 146 nsew signal input
flabel metal2 s 46592 0 46704 800 0 FreeSans 448 90 0 0 la_oenb[24]
port 147 nsew signal input
flabel metal2 s 47264 0 47376 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 148 nsew signal input
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 la_oenb[26]
port 149 nsew signal input
flabel metal2 s 48608 0 48720 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 150 nsew signal input
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 la_oenb[28]
port 151 nsew signal input
flabel metal2 s 49952 0 50064 800 0 FreeSans 448 90 0 0 la_oenb[29]
port 152 nsew signal input
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 153 nsew signal input
flabel metal2 s 50624 0 50736 800 0 FreeSans 448 90 0 0 la_oenb[30]
port 154 nsew signal input
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 la_oenb[31]
port 155 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 la_oenb[32]
port 156 nsew signal input
flabel metal2 s 52640 0 52752 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 157 nsew signal input
flabel metal2 s 53312 0 53424 800 0 FreeSans 448 90 0 0 la_oenb[34]
port 158 nsew signal input
flabel metal2 s 53984 0 54096 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 159 nsew signal input
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 160 nsew signal input
flabel metal2 s 55328 0 55440 800 0 FreeSans 448 90 0 0 la_oenb[37]
port 161 nsew signal input
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 162 nsew signal input
flabel metal2 s 56672 0 56784 800 0 FreeSans 448 90 0 0 la_oenb[39]
port 163 nsew signal input
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 164 nsew signal input
flabel metal2 s 57344 0 57456 800 0 FreeSans 448 90 0 0 la_oenb[40]
port 165 nsew signal input
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 la_oenb[41]
port 166 nsew signal input
flabel metal2 s 58688 0 58800 800 0 FreeSans 448 90 0 0 la_oenb[42]
port 167 nsew signal input
flabel metal2 s 59360 0 59472 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 168 nsew signal input
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 169 nsew signal input
flabel metal2 s 60704 0 60816 800 0 FreeSans 448 90 0 0 la_oenb[45]
port 170 nsew signal input
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 171 nsew signal input
flabel metal2 s 62048 0 62160 800 0 FreeSans 448 90 0 0 la_oenb[47]
port 172 nsew signal input
flabel metal2 s 62720 0 62832 800 0 FreeSans 448 90 0 0 la_oenb[48]
port 173 nsew signal input
flabel metal2 s 63392 0 63504 800 0 FreeSans 448 90 0 0 la_oenb[49]
port 174 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 la_oenb[4]
port 175 nsew signal input
flabel metal2 s 64064 0 64176 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 176 nsew signal input
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 la_oenb[51]
port 177 nsew signal input
flabel metal2 s 65408 0 65520 800 0 FreeSans 448 90 0 0 la_oenb[52]
port 178 nsew signal input
flabel metal2 s 66080 0 66192 800 0 FreeSans 448 90 0 0 la_oenb[53]
port 179 nsew signal input
flabel metal2 s 66752 0 66864 800 0 FreeSans 448 90 0 0 la_oenb[54]
port 180 nsew signal input
flabel metal2 s 67424 0 67536 800 0 FreeSans 448 90 0 0 la_oenb[55]
port 181 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 182 nsew signal input
flabel metal2 s 68768 0 68880 800 0 FreeSans 448 90 0 0 la_oenb[57]
port 183 nsew signal input
flabel metal2 s 69440 0 69552 800 0 FreeSans 448 90 0 0 la_oenb[58]
port 184 nsew signal input
flabel metal2 s 70112 0 70224 800 0 FreeSans 448 90 0 0 la_oenb[59]
port 185 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 186 nsew signal input
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 la_oenb[60]
port 187 nsew signal input
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 188 nsew signal input
flabel metal2 s 72128 0 72240 800 0 FreeSans 448 90 0 0 la_oenb[62]
port 189 nsew signal input
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 la_oenb[63]
port 190 nsew signal input
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 la_oenb[6]
port 191 nsew signal input
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 192 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 la_oenb[8]
port 193 nsew signal input
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 la_oenb[9]
port 194 nsew signal input
flabel metal4 s 10844 3076 11164 36908 0 FreeSans 1280 90 0 0 vdd
port 195 nsew power bidirectional
flabel metal4 s 30164 3076 30484 36908 0 FreeSans 1280 90 0 0 vdd
port 195 nsew power bidirectional
flabel metal4 s 49484 3076 49804 36908 0 FreeSans 1280 90 0 0 vdd
port 195 nsew power bidirectional
flabel metal4 s 68804 3076 69124 36908 0 FreeSans 1280 90 0 0 vdd
port 195 nsew power bidirectional
flabel metal4 s 20504 3076 20824 36908 0 FreeSans 1280 90 0 0 vss
port 196 nsew ground bidirectional
flabel metal4 s 39824 3076 40144 36908 0 FreeSans 1280 90 0 0 vss
port 196 nsew ground bidirectional
flabel metal4 s 59144 3076 59464 36908 0 FreeSans 1280 90 0 0 vss
port 196 nsew ground bidirectional
flabel metal4 s 78464 3076 78784 36908 0 FreeSans 1280 90 0 0 vss
port 196 nsew ground bidirectional
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 wb_clk_i
port 197 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 wb_rst_i
port 198 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 199 nsew signal tristate
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 200 nsew signal input
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 201 nsew signal input
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 202 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 203 nsew signal input
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 204 nsew signal input
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 205 nsew signal input
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 206 nsew signal input
flabel metal2 s 19264 0 19376 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 207 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 208 nsew signal input
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 209 nsew signal input
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 210 nsew signal input
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 211 nsew signal input
flabel metal2 s 21952 0 22064 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 212 nsew signal input
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 213 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 214 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 215 nsew signal input
flabel metal2 s 24640 0 24752 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 216 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 217 nsew signal input
flabel metal2 s 25984 0 26096 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 218 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 219 nsew signal input
flabel metal2 s 27328 0 27440 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 220 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 221 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 222 nsew signal input
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 223 nsew signal input
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 224 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 225 nsew signal input
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 226 nsew signal input
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 227 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 228 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 229 nsew signal input
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 230 nsew signal input
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 231 nsew signal input
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 232 nsew signal input
flabel metal2 s 7840 0 7952 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 233 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 234 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 235 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 236 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 237 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 238 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 239 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 240 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 241 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 242 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 243 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 244 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 245 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 246 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 247 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 248 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 249 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 250 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 251 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 252 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 253 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 254 nsew signal input
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 255 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 256 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 257 nsew signal input
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 258 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 259 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 260 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 261 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 262 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 263 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 264 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 265 nsew signal tristate
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 266 nsew signal tristate
flabel metal2 s 16352 0 16464 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 267 nsew signal tristate
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 268 nsew signal tristate
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 269 nsew signal tristate
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 270 nsew signal tristate
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 271 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 272 nsew signal tristate
flabel metal2 s 20384 0 20496 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 273 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 274 nsew signal tristate
flabel metal2 s 21728 0 21840 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 275 nsew signal tristate
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 276 nsew signal tristate
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 277 nsew signal tristate
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 278 nsew signal tristate
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 279 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 280 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 281 nsew signal tristate
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 282 nsew signal tristate
flabel metal2 s 26432 0 26544 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 283 nsew signal tristate
flabel metal2 s 27104 0 27216 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 284 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 285 nsew signal tristate
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 286 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 287 nsew signal tristate
flabel metal2 s 29120 0 29232 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 288 nsew signal tristate
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 289 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 290 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 291 nsew signal tristate
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 292 nsew signal tristate
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 293 nsew signal tristate
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 294 nsew signal tristate
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 295 nsew signal tristate
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 296 nsew signal tristate
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 297 nsew signal input
flabel metal2 s 9184 0 9296 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 298 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 299 nsew signal input
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 300 nsew signal input
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 301 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 wbs_we_i
port 302 nsew signal input
rlabel metal1 39984 36848 39984 36848 0 vdd
rlabel via1 40064 36064 40064 36064 0 vss
rlabel metal3 19040 5096 19040 5096 0 _000_
rlabel metal2 29400 11872 29400 11872 0 _001_
rlabel metal3 26600 7560 26600 7560 0 _002_
rlabel metal2 25592 7952 25592 7952 0 _003_
rlabel metal2 26488 9464 26488 9464 0 _004_
rlabel metal3 33152 12040 33152 12040 0 _005_
rlabel metal2 34664 12712 34664 12712 0 _006_
rlabel metal2 33432 13104 33432 13104 0 _007_
rlabel metal2 38696 11592 38696 11592 0 _008_
rlabel metal2 38136 12656 38136 12656 0 _009_
rlabel metal2 42056 9912 42056 9912 0 _010_
rlabel metal2 53032 8232 53032 8232 0 _011_
rlabel metal3 53088 9128 53088 9128 0 _012_
rlabel metal2 48832 8904 48832 8904 0 _013_
rlabel metal2 43288 11872 43288 11872 0 _014_
rlabel metal2 44184 9632 44184 9632 0 _015_
rlabel metal2 47936 9240 47936 9240 0 _016_
rlabel metal2 17864 5544 17864 5544 0 _017_
rlabel metal2 6664 6608 6664 6608 0 _018_
rlabel metal2 9184 5208 9184 5208 0 _019_
rlabel metal2 13048 6216 13048 6216 0 _020_
rlabel metal3 10136 8232 10136 8232 0 _021_
rlabel metal2 10304 9688 10304 9688 0 _022_
rlabel metal2 11256 12600 11256 12600 0 _023_
rlabel metal2 14392 12488 14392 12488 0 _024_
rlabel metal2 22008 6048 22008 6048 0 _025_
rlabel metal3 19992 12264 19992 12264 0 _026_
rlabel metal2 20328 8400 20328 8400 0 _027_
rlabel metal2 16072 8456 16072 8456 0 _028_
rlabel metal2 22120 10528 22120 10528 0 _029_
rlabel metal2 17528 9464 17528 9464 0 _030_
rlabel metal2 16744 7224 16744 7224 0 _031_
rlabel metal2 25592 11032 25592 11032 0 _032_
rlabel metal3 60144 5880 60144 5880 0 _033_
rlabel metal3 53200 7672 53200 7672 0 _034_
rlabel metal2 55328 5992 55328 5992 0 _035_
rlabel metal2 54824 7952 54824 7952 0 _036_
rlabel metal2 49784 7784 49784 7784 0 _037_
rlabel metal2 70168 10304 70168 10304 0 _038_
rlabel metal2 23576 8624 23576 8624 0 _039_
rlabel metal2 23688 10584 23688 10584 0 _040_
rlabel metal2 25704 3360 25704 3360 0 _041_
rlabel metal2 39760 10696 39760 10696 0 _042_
rlabel metal3 56672 7448 56672 7448 0 _043_
rlabel metal3 32200 15512 32200 15512 0 _044_
rlabel metal2 19880 9520 19880 9520 0 _045_
rlabel metal3 25480 12712 25480 12712 0 _046_
rlabel metal2 55272 5040 55272 5040 0 _047_
rlabel metal2 55496 3864 55496 3864 0 _048_
rlabel metal2 59752 4200 59752 4200 0 _049_
rlabel metal2 59976 4312 59976 4312 0 _050_
rlabel metal3 62888 6776 62888 6776 0 _051_
rlabel metal3 63056 8232 63056 8232 0 _052_
rlabel metal2 60032 6440 60032 6440 0 _053_
rlabel metal2 62776 4872 62776 4872 0 _054_
rlabel metal3 62048 5880 62048 5880 0 _055_
rlabel metal2 63784 7056 63784 7056 0 _056_
rlabel metal2 44296 7728 44296 7728 0 _057_
rlabel metal2 59752 5712 59752 5712 0 _058_
rlabel metal2 59696 6440 59696 6440 0 _059_
rlabel metal2 43848 7728 43848 7728 0 _060_
rlabel metal2 59416 3976 59416 3976 0 _061_
rlabel metal3 60032 2968 60032 2968 0 _062_
rlabel metal2 59528 4032 59528 4032 0 _063_
rlabel metal2 54824 4592 54824 4592 0 _064_
rlabel metal2 39032 7616 39032 7616 0 _065_
rlabel metal2 23744 12712 23744 12712 0 _066_
rlabel metal2 26152 4256 26152 4256 0 _067_
rlabel metal2 23128 6272 23128 6272 0 _068_
rlabel metal2 17640 4984 17640 4984 0 _069_
rlabel metal2 23352 4480 23352 4480 0 _070_
rlabel metal3 22904 5096 22904 5096 0 _071_
rlabel metal3 23800 5320 23800 5320 0 _072_
rlabel metal2 25032 7560 25032 7560 0 _073_
rlabel metal2 25704 8288 25704 8288 0 _074_
rlabel metal3 42448 16968 42448 16968 0 _075_
rlabel metal2 23184 12040 23184 12040 0 _076_
rlabel metal2 26936 4088 26936 4088 0 _077_
rlabel metal2 27384 3920 27384 3920 0 _078_
rlabel metal3 28560 3192 28560 3192 0 _079_
rlabel metal2 26320 3416 26320 3416 0 _080_
rlabel metal3 24640 6440 24640 6440 0 _081_
rlabel metal2 25592 4704 25592 4704 0 _082_
rlabel metal3 25088 3752 25088 3752 0 _083_
rlabel metal3 27496 3304 27496 3304 0 _084_
rlabel metal2 58408 7952 58408 7952 0 _085_
rlabel metal2 57960 7672 57960 7672 0 _086_
rlabel metal2 26824 7000 26824 7000 0 _087_
rlabel metal2 29064 5488 29064 5488 0 _088_
rlabel metal3 25144 4312 25144 4312 0 _089_
rlabel metal2 29400 5096 29400 5096 0 _090_
rlabel metal3 54152 3640 54152 3640 0 _091_
rlabel metal3 41048 13216 41048 13216 0 _092_
rlabel metal3 40824 6664 40824 6664 0 _093_
rlabel metal3 36512 7448 36512 7448 0 _094_
rlabel metal2 33544 7840 33544 7840 0 _095_
rlabel metal2 25256 5600 25256 5600 0 _096_
rlabel metal2 33432 6048 33432 6048 0 _097_
rlabel metal2 35560 8736 35560 8736 0 _098_
rlabel metal3 33376 14056 33376 14056 0 _099_
rlabel metal2 37128 12992 37128 12992 0 _100_
rlabel metal2 56840 3192 56840 3192 0 _101_
rlabel metal3 36792 10024 36792 10024 0 _102_
rlabel metal3 34888 13384 34888 13384 0 _103_
rlabel metal2 32536 5656 32536 5656 0 _104_
rlabel metal2 32424 3696 32424 3696 0 _105_
rlabel metal2 38248 6720 38248 6720 0 _106_
rlabel metal2 36176 10696 36176 10696 0 _107_
rlabel metal2 39648 4200 39648 4200 0 _108_
rlabel metal2 39592 5488 39592 5488 0 _109_
rlabel metal2 33880 6440 33880 6440 0 _110_
rlabel metal2 40264 8008 40264 8008 0 _111_
rlabel metal3 45640 5040 45640 5040 0 _112_
rlabel metal3 39704 6552 39704 6552 0 _113_
rlabel metal3 33040 16856 33040 16856 0 _114_
rlabel metal2 39928 9632 39928 9632 0 _115_
rlabel metal3 20888 1344 20888 1344 0 _116_
rlabel metal2 44968 3920 44968 3920 0 _117_
rlabel metal2 44744 3136 44744 3136 0 _118_
rlabel metal3 40432 7448 40432 7448 0 _119_
rlabel metal2 38304 7336 38304 7336 0 _120_
rlabel metal2 40936 9296 40936 9296 0 _121_
rlabel metal2 42280 6048 42280 6048 0 _122_
rlabel metal2 48664 5824 48664 5824 0 _123_
rlabel metal3 43288 4312 43288 4312 0 _124_
rlabel metal2 42952 6832 42952 6832 0 _125_
rlabel metal2 37464 8120 37464 8120 0 _126_
rlabel metal2 41048 9408 41048 9408 0 _127_
rlabel metal2 41384 8736 41384 8736 0 _128_
rlabel metal2 41720 9464 41720 9464 0 _129_
rlabel metal2 42728 6384 42728 6384 0 _130_
rlabel metal2 50568 9520 50568 9520 0 _131_
rlabel metal3 44408 11928 44408 11928 0 _132_
rlabel metal2 48216 5432 48216 5432 0 _133_
rlabel metal2 49000 5320 49000 5320 0 _134_
rlabel metal2 52360 4592 52360 4592 0 _135_
rlabel metal2 51800 7056 51800 7056 0 _136_
rlabel metal2 50680 7840 50680 7840 0 _137_
rlabel metal3 21392 17080 21392 17080 0 _138_
rlabel metal2 16072 3108 16072 3108 0 _139_
rlabel metal2 41104 5880 41104 5880 0 _140_
rlabel metal2 46760 9408 46760 9408 0 _141_
rlabel metal2 51464 7000 51464 7000 0 _142_
rlabel metal2 51464 5992 51464 5992 0 _143_
rlabel metal2 46368 12152 46368 12152 0 _144_
rlabel metal2 22904 8736 22904 8736 0 _145_
rlabel metal3 45584 3416 45584 3416 0 _146_
rlabel metal2 46984 3360 46984 3360 0 _147_
rlabel metal2 17976 11984 17976 11984 0 _148_
rlabel metal2 39928 5992 39928 5992 0 _149_
rlabel metal2 44072 9856 44072 9856 0 _150_
rlabel metal2 45080 8400 45080 8400 0 _151_
rlabel metal2 43736 9072 43736 9072 0 _152_
rlabel metal2 52696 3976 52696 3976 0 _153_
rlabel metal2 44296 4536 44296 4536 0 _154_
rlabel metal2 43176 7112 43176 7112 0 _155_
rlabel metal2 16968 11200 16968 11200 0 _156_
rlabel metal2 45192 5208 45192 5208 0 _157_
rlabel metal2 44632 4928 44632 4928 0 _158_
rlabel metal2 56056 2296 56056 2296 0 _159_
rlabel metal2 44072 5824 44072 5824 0 _160_
rlabel metal2 47544 9520 47544 9520 0 _161_
rlabel metal2 47208 7840 47208 7840 0 _162_
rlabel metal2 47880 7896 47880 7896 0 _163_
rlabel metal2 18200 7728 18200 7728 0 _164_
rlabel metal2 17304 6048 17304 6048 0 _165_
rlabel metal2 17304 4424 17304 4424 0 _166_
rlabel via2 15736 5992 15736 5992 0 _167_
rlabel metal2 9688 6272 9688 6272 0 _168_
rlabel metal2 7896 7672 7896 7672 0 _169_
rlabel metal3 13608 6664 13608 6664 0 _170_
rlabel metal2 13160 11704 13160 11704 0 _171_
rlabel metal2 10920 9016 10920 9016 0 _172_
rlabel metal2 10920 9688 10920 9688 0 _173_
rlabel metal2 11816 12152 11816 12152 0 _174_
rlabel metal2 14168 11760 14168 11760 0 _175_
rlabel metal3 16464 8232 16464 8232 0 _176_
rlabel metal3 21112 6664 21112 6664 0 _177_
rlabel metal2 19544 12264 19544 12264 0 _178_
rlabel metal2 19880 8288 19880 8288 0 _179_
rlabel metal2 17640 6160 17640 6160 0 _180_
rlabel metal2 22568 10248 22568 10248 0 _181_
rlabel metal2 17864 8736 17864 8736 0 _182_
rlabel metal2 21280 5096 21280 5096 0 _183_
rlabel metal3 24920 10696 24920 10696 0 _184_
rlabel metal2 40936 11200 40936 11200 0 clknet_0_counter.clk
rlabel metal2 22568 12544 22568 12544 0 clknet_2_0__leaf_counter.clk
rlabel metal2 15288 11088 15288 11088 0 clknet_2_1__leaf_counter.clk
rlabel metal2 41496 10192 41496 10192 0 clknet_2_2__leaf_counter.clk
rlabel metal2 30856 10528 30856 10528 0 clknet_2_3__leaf_counter.clk
rlabel metal2 34440 8344 34440 8344 0 counter.clk
rlabel metal2 62552 3920 62552 3920 0 la_data_in[46]
rlabel metal2 67256 4760 67256 4760 0 la_data_in[47]
rlabel metal3 65912 3696 65912 3696 0 la_data_in[48]
rlabel metal3 63504 6552 63504 6552 0 la_data_in[49]
rlabel metal2 63672 2058 63672 2058 0 la_data_in[50]
rlabel metal2 71288 7616 71288 7616 0 la_data_in[51]
rlabel metal2 70056 7504 70056 7504 0 la_data_in[52]
rlabel metal2 65688 1638 65688 1638 0 la_data_in[53]
rlabel metal3 66696 7560 66696 7560 0 la_data_in[54]
rlabel metal3 67872 6552 67872 6552 0 la_data_in[55]
rlabel metal2 77616 4984 77616 4984 0 la_data_in[56]
rlabel metal2 68376 1918 68376 1918 0 la_data_in[57]
rlabel metal2 74984 4256 74984 4256 0 la_data_in[58]
rlabel metal2 74760 6832 74760 6832 0 la_data_in[59]
rlabel metal2 70448 3192 70448 3192 0 la_data_in[60]
rlabel metal2 71064 2058 71064 2058 0 la_data_in[61]
rlabel metal2 71736 1526 71736 1526 0 la_data_in[62]
rlabel metal2 76328 5880 76328 5880 0 la_data_in[63]
rlabel metal2 30296 2058 30296 2058 0 la_data_out[0]
rlabel metal2 37016 854 37016 854 0 la_data_out[10]
rlabel metal2 37688 2086 37688 2086 0 la_data_out[11]
rlabel metal2 38360 2478 38360 2478 0 la_data_out[12]
rlabel metal2 39032 854 39032 854 0 la_data_out[13]
rlabel metal2 39816 4088 39816 4088 0 la_data_out[14]
rlabel metal2 40376 2058 40376 2058 0 la_data_out[15]
rlabel metal3 31472 4872 31472 4872 0 la_data_out[1]
rlabel metal2 31640 2058 31640 2058 0 la_data_out[2]
rlabel metal2 32312 1022 32312 1022 0 la_data_out[3]
rlabel metal2 32984 2982 32984 2982 0 la_data_out[4]
rlabel metal2 33656 2058 33656 2058 0 la_data_out[5]
rlabel metal2 34440 5656 34440 5656 0 la_data_out[6]
rlabel metal2 35000 2058 35000 2058 0 la_data_out[7]
rlabel metal3 35056 3640 35056 3640 0 la_data_out[8]
rlabel metal2 36344 1022 36344 1022 0 la_data_out[9]
rlabel metal3 68320 4984 68320 4984 0 la_oenb[46]
rlabel metal2 62888 3696 62888 3696 0 la_oenb[47]
rlabel metal2 68488 3080 68488 3080 0 la_oenb[48]
rlabel metal3 63504 4424 63504 4424 0 la_oenb[49]
rlabel metal2 65128 5600 65128 5600 0 la_oenb[50]
rlabel metal2 64792 2058 64792 2058 0 la_oenb[51]
rlabel metal2 76104 3976 76104 3976 0 la_oenb[52]
rlabel metal2 70336 3416 70336 3416 0 la_oenb[53]
rlabel metal2 70392 5824 70392 5824 0 la_oenb[54]
rlabel metal1 67760 2968 67760 2968 0 la_oenb[55]
rlabel metal2 73192 4648 73192 4648 0 la_oenb[56]
rlabel metal2 74312 4256 74312 4256 0 la_oenb[57]
rlabel metal2 75208 5824 75208 5824 0 la_oenb[58]
rlabel metal2 72408 6328 72408 6328 0 la_oenb[59]
rlabel metal2 73584 6552 73584 6552 0 la_oenb[60]
rlabel metal2 75152 4424 75152 4424 0 la_oenb[61]
rlabel metal2 78120 3472 78120 3472 0 la_oenb[62]
rlabel metal2 74424 6272 74424 6272 0 la_oenb[63]
rlabel metal2 48328 5544 48328 5544 0 net1
rlabel metal2 76888 10248 76888 10248 0 net10
rlabel metal2 50456 2058 50456 2058 0 net100
rlabel metal2 51128 1246 51128 1246 0 net101
rlabel metal2 51688 3864 51688 3864 0 net102
rlabel metal2 52472 2758 52472 2758 0 net103
rlabel metal3 54320 4984 54320 4984 0 net104
rlabel metal3 54880 8008 54880 8008 0 net105
rlabel metal3 55440 6888 55440 6888 0 net106
rlabel metal2 55104 3640 55104 3640 0 net107
rlabel metal2 55832 1246 55832 1246 0 net108
rlabel metal3 56840 3752 56840 3752 0 net109
rlabel metal2 71736 9464 71736 9464 0 net11
rlabel metal2 57176 2142 57176 2142 0 net110
rlabel metal2 57848 2254 57848 2254 0 net111
rlabel metal2 58520 3318 58520 3318 0 net112
rlabel metal2 59192 1750 59192 1750 0 net113
rlabel metal2 59864 1974 59864 1974 0 net114
rlabel metal1 61096 8792 61096 8792 0 net115
rlabel metal2 61208 2058 61208 2058 0 net116
rlabel metal2 61880 2030 61880 2030 0 net117
rlabel metal2 62552 1862 62552 1862 0 net118
rlabel metal2 63224 2702 63224 2702 0 net119
rlabel metal2 77560 10304 77560 10304 0 net12
rlabel metal2 63896 1862 63896 1862 0 net120
rlabel metal2 64568 2254 64568 2254 0 net121
rlabel metal2 71512 7168 71512 7168 0 net122
rlabel metal3 66864 4984 66864 4984 0 net123
rlabel metal2 66584 2590 66584 2590 0 net124
rlabel metal2 67256 2422 67256 2422 0 net125
rlabel metal2 67928 2814 67928 2814 0 net126
rlabel metal2 68768 4536 68768 4536 0 net127
rlabel metal2 69272 1918 69272 1918 0 net128
rlabel metal2 69944 1918 69944 1918 0 net129
rlabel metal3 67368 3304 67368 3304 0 net13
rlabel metal2 70616 2870 70616 2870 0 net130
rlabel metal2 71288 2058 71288 2058 0 net131
rlabel metal2 78120 4312 78120 4312 0 net132
rlabel metal2 74368 9576 74368 9576 0 net133
rlabel metal2 19768 2058 19768 2058 0 net134
rlabel metal2 20496 6440 20496 6440 0 net135
rlabel metal2 21112 2758 21112 2758 0 net136
rlabel metal2 21616 5656 21616 5656 0 net137
rlabel metal2 22456 2702 22456 2702 0 net138
rlabel metal2 23128 2058 23128 2058 0 net139
rlabel metal2 70728 10528 70728 10528 0 net14
rlabel metal3 23352 4872 23352 4872 0 net140
rlabel metal2 24472 3766 24472 3766 0 net141
rlabel metal3 24472 3640 24472 3640 0 net142
rlabel metal3 25368 4760 25368 4760 0 net143
rlabel metal2 26488 854 26488 854 0 net144
rlabel metal3 16968 560 16968 560 0 net145
rlabel metal2 27832 1022 27832 1022 0 net146
rlabel metal2 28504 3486 28504 3486 0 net147
rlabel metal2 29176 1862 29176 1862 0 net148
rlabel metal2 24696 3360 24696 3360 0 net149
rlabel metal2 78008 3696 78008 3696 0 net15
rlabel metal3 75964 6440 75964 6440 0 net150
rlabel metal2 76104 9576 76104 9576 0 net151
rlabel metal2 73528 1974 73528 1974 0 net152
rlabel metal2 41048 2086 41048 2086 0 net153
rlabel metal2 41720 2058 41720 2058 0 net154
rlabel metal2 55720 1512 55720 1512 0 net155
rlabel metal2 49672 8904 49672 8904 0 net156
rlabel metal2 49448 8960 49448 8960 0 net157
rlabel metal2 43120 11816 43120 11816 0 net158
rlabel metal2 45080 1638 45080 1638 0 net159
rlabel metal2 75656 4592 75656 4592 0 net16
rlabel metal2 45752 1526 45752 1526 0 net160
rlabel metal3 50008 10920 50008 10920 0 net161
rlabel metal2 78232 6384 78232 6384 0 net162
rlabel metal2 59080 2268 59080 2268 0 net163
rlabel metal2 44408 11312 44408 11312 0 net164
rlabel metal3 45304 8904 45304 8904 0 net165
rlabel metal2 70952 9520 70952 9520 0 net166
rlabel metal3 50792 1680 50792 1680 0 net167
rlabel metal2 43512 10640 43512 10640 0 net168
rlabel metal2 44072 12656 44072 12656 0 net169
rlabel metal3 74088 9128 74088 9128 0 net17
rlabel metal2 77112 9688 77112 9688 0 net170
rlabel metal2 57568 4200 57568 4200 0 net171
rlabel metal2 42504 9128 42504 9128 0 net172
rlabel metal2 41104 11256 41104 11256 0 net173
rlabel metal2 76216 6664 76216 6664 0 net174
rlabel metal2 52808 4816 52808 4816 0 net175
rlabel metal2 52136 5432 52136 5432 0 net176
rlabel metal2 52360 7952 52360 7952 0 net177
rlabel metal2 75600 8904 75600 8904 0 net178
rlabel metal3 59080 6832 59080 6832 0 net179
rlabel metal2 77560 8624 77560 8624 0 net18
rlabel metal2 50232 6160 50232 6160 0 net180
rlabel metal3 53312 8904 53312 8904 0 net181
rlabel metal2 78120 6608 78120 6608 0 net182
rlabel metal3 49000 6608 49000 6608 0 net183
rlabel metal2 48664 8456 48664 8456 0 net184
rlabel metal2 48440 10864 48440 10864 0 net185
rlabel metal2 74088 7448 74088 7448 0 net186
rlabel metal2 63168 4872 63168 4872 0 net187
rlabel metal2 49224 7280 49224 7280 0 net188
rlabel metal2 49336 10136 49336 10136 0 net189
rlabel metal2 69160 3192 69160 3192 0 net19
rlabel metal2 67816 8848 67816 8848 0 net190
rlabel metal2 42840 6160 42840 6160 0 net191
rlabel metal2 41944 9296 41944 9296 0 net192
rlabel metal2 38920 13328 38920 13328 0 net193
rlabel metal2 63896 8736 63896 8736 0 net194
rlabel metal2 28168 5208 28168 5208 0 net195
rlabel metal2 26040 6104 26040 6104 0 net196
rlabel metal2 27720 8568 27720 8568 0 net197
rlabel metal2 65688 8904 65688 8904 0 net198
rlabel metal3 37968 17080 37968 17080 0 net199
rlabel metal2 63560 9688 63560 9688 0 net2
rlabel metal2 55832 6216 55832 6216 0 net20
rlabel metal2 27384 5432 27384 5432 0 net200
rlabel metal3 26152 8344 26152 8344 0 net201
rlabel metal3 70392 8848 70392 8848 0 net202
rlabel metal2 50344 3864 50344 3864 0 net203
rlabel metal2 38920 10976 38920 10976 0 net204
rlabel metal2 35672 11088 35672 11088 0 net205
rlabel metal2 67144 8176 67144 8176 0 net206
rlabel metal2 40544 12376 40544 12376 0 net207
rlabel metal2 39144 10416 39144 10416 0 net208
rlabel metal2 35672 13328 35672 13328 0 net209
rlabel metal3 64064 6440 64064 6440 0 net21
rlabel metal2 65800 3864 65800 3864 0 net210
rlabel metal2 47992 5600 47992 5600 0 net211
rlabel metal2 30968 8064 30968 8064 0 net212
rlabel metal2 30184 10976 30184 10976 0 net213
rlabel metal2 64904 8736 64904 8736 0 net214
rlabel metal3 29624 15848 29624 15848 0 net215
rlabel metal2 28168 5544 28168 5544 0 net216
rlabel metal3 28784 9912 28784 9912 0 net217
rlabel metal2 66920 8288 66920 8288 0 net218
rlabel metal2 31976 15624 31976 15624 0 net219
rlabel metal2 63672 8288 63672 8288 0 net22
rlabel metal2 32480 15624 32480 15624 0 net220
rlabel metal2 34832 9912 34832 9912 0 net221
rlabel metal2 68264 8624 68264 8624 0 net222
rlabel metal2 39144 7672 39144 7672 0 net223
rlabel metal2 34776 11984 34776 11984 0 net224
rlabel metal2 32200 10640 32200 10640 0 net225
rlabel metal2 77672 7588 77672 7588 0 net226
rlabel metal2 76216 8512 76216 8512 0 net227
rlabel metal2 40824 12544 40824 12544 0 net228
rlabel metal2 76384 9016 76384 9016 0 net229
rlabel metal2 55384 4144 55384 4144 0 net23
rlabel metal2 70616 7392 70616 7392 0 net230
rlabel metal2 43400 8848 43400 8848 0 net231
rlabel metal2 72184 5600 72184 5600 0 net232
rlabel metal2 74536 7280 74536 7280 0 net233
rlabel metal2 47544 12432 47544 12432 0 net234
rlabel metal2 71288 5544 71288 5544 0 net235
rlabel metal2 77336 5824 77336 5824 0 net236
rlabel metal2 77112 5152 77112 5152 0 net237
rlabel metal2 75656 7168 75656 7168 0 net238
rlabel metal2 47208 8904 47208 8904 0 net239
rlabel metal3 56224 2744 56224 2744 0 net24
rlabel metal2 66696 4368 66696 4368 0 net240
rlabel metal2 72632 5544 72632 5544 0 net241
rlabel metal2 65352 5376 65352 5376 0 net242
rlabel metal2 77840 7000 77840 7000 0 net243
rlabel metal2 67368 6496 67368 6496 0 net244
rlabel metal2 66360 5152 66360 5152 0 net245
rlabel metal2 69552 3528 69552 3528 0 net246
rlabel metal2 69496 4312 69496 4312 0 net247
rlabel metal2 73752 3416 73752 3416 0 net248
rlabel metal2 73192 3080 73192 3080 0 net25
rlabel metal2 70840 6748 70840 6748 0 net26
rlabel metal2 66920 7616 66920 7616 0 net27
rlabel metal2 67704 6832 67704 6832 0 net28
rlabel metal2 70504 5880 70504 5880 0 net29
rlabel metal2 65296 9240 65296 9240 0 net3
rlabel metal2 60200 9408 60200 9408 0 net30
rlabel metal2 77672 9688 77672 9688 0 net31
rlabel metal3 72968 8848 72968 8848 0 net32
rlabel metal2 77560 6216 77560 6216 0 net33
rlabel metal2 77112 7784 77112 7784 0 net34
rlabel metal2 77896 3808 77896 3808 0 net35
rlabel metal2 75880 9520 75880 9520 0 net36
rlabel metal3 36008 17416 36008 17416 0 net37
rlabel metal2 64568 8960 64568 8960 0 net38
rlabel metal2 22008 5432 22008 5432 0 net39
rlabel metal2 53592 10416 53592 10416 0 net4
rlabel metal2 5880 2184 5880 2184 0 net40
rlabel metal2 18648 3052 18648 3052 0 net41
rlabel metal2 19488 6104 19488 6104 0 net42
rlabel metal2 9688 3136 9688 3136 0 net43
rlabel metal2 13832 2352 13832 2352 0 net44
rlabel metal3 18984 784 18984 784 0 net45
rlabel metal3 9016 4536 9016 4536 0 net46
rlabel metal2 23240 6552 23240 6552 0 net47
rlabel metal2 23128 5432 23128 5432 0 net48
rlabel metal3 21000 12320 21000 12320 0 net49
rlabel metal2 66696 8344 66696 8344 0 net5
rlabel metal2 10696 8232 10696 8232 0 net50
rlabel metal2 3192 2856 3192 2856 0 net51
rlabel metal2 25032 5656 25032 5656 0 net52
rlabel metal2 14784 9688 14784 9688 0 net53
rlabel metal3 23744 3528 23744 3528 0 net54
rlabel metal2 2576 4536 2576 4536 0 net55
rlabel metal2 2520 3584 2520 3584 0 net56
rlabel metal3 29624 15288 29624 15288 0 net57
rlabel metal3 7896 5208 7896 5208 0 net58
rlabel metal2 28056 10304 28056 10304 0 net59
rlabel metal3 63364 9128 63364 9128 0 net6
rlabel metal2 38472 14280 38472 14280 0 net60
rlabel metal2 42504 12376 42504 12376 0 net61
rlabel metal2 47096 9856 47096 9856 0 net62
rlabel metal2 41832 12096 41832 12096 0 net63
rlabel metal2 43064 5432 43064 5432 0 net64
rlabel metal2 24248 12264 24248 12264 0 net65
rlabel metal2 31192 5600 31192 5600 0 net66
rlabel metal2 24696 7952 24696 7952 0 net67
rlabel metal2 15064 8736 15064 8736 0 net68
rlabel metal2 32648 9408 32648 9408 0 net69
rlabel metal2 58184 8400 58184 8400 0 net7
rlabel metal3 21000 8848 21000 8848 0 net70
rlabel metal3 35280 9800 35280 9800 0 net71
rlabel metal3 19320 10752 19320 10752 0 net72
rlabel metal2 35168 7448 35168 7448 0 net73
rlabel metal2 21504 11144 21504 11144 0 net74
rlabel metal2 16688 18536 16688 18536 0 net75
rlabel metal2 16072 5936 16072 5936 0 net76
rlabel metal2 19208 7168 19208 7168 0 net77
rlabel metal3 17416 5824 17416 5824 0 net78
rlabel metal2 24248 9576 24248 9576 0 net79
rlabel metal2 69272 9632 69272 9632 0 net8
rlabel metal2 17920 8232 17920 8232 0 net80
rlabel metal3 19152 5208 19152 5208 0 net81
rlabel metal3 22624 11480 22624 11480 0 net82
rlabel metal2 10584 5824 10584 5824 0 net83
rlabel metal2 7112 5432 7112 5432 0 net84
rlabel metal2 13720 5936 13720 5936 0 net85
rlabel metal2 12040 7504 12040 7504 0 net86
rlabel metal2 12488 9688 12488 9688 0 net87
rlabel metal2 12936 12040 12936 12040 0 net88
rlabel metal2 16520 9744 16520 9744 0 net89
rlabel metal3 62776 11928 62776 11928 0 net9
rlabel metal2 19880 5320 19880 5320 0 net90
rlabel metal2 18200 11088 18200 11088 0 net91
rlabel metal3 26096 4872 26096 4872 0 net92
rlabel metal2 13384 10080 13384 10080 0 net93
rlabel metal2 26712 11984 26712 11984 0 net94
rlabel metal2 47096 2366 47096 2366 0 net95
rlabel metal2 47768 1974 47768 1974 0 net96
rlabel metal2 48440 2058 48440 2058 0 net97
rlabel metal2 49168 12264 49168 12264 0 net98
rlabel metal2 49784 2198 49784 2198 0 net99
rlabel metal3 38136 15176 38136 15176 0 wb_clk_i
rlabel metal2 4648 4984 4648 4984 0 wb_rst_i
rlabel metal2 6776 1806 6776 1806 0 wbs_ack_o
rlabel metal2 2968 4368 2968 4368 0 wbs_cyc_i
rlabel metal2 4760 5992 4760 5992 0 wbs_dat_i[0]
rlabel metal2 3304 4032 3304 4032 0 wbs_dat_i[10]
rlabel metal2 18536 7000 18536 7000 0 wbs_dat_i[11]
rlabel metal2 19320 6104 19320 6104 0 wbs_dat_i[12]
rlabel metal2 17528 1302 17528 1302 0 wbs_dat_i[13]
rlabel metal2 18200 2142 18200 2142 0 wbs_dat_i[14]
rlabel metal2 18816 4312 18816 4312 0 wbs_dat_i[15]
rlabel metal2 8792 2058 8792 2058 0 wbs_dat_i[1]
rlabel metal2 9688 1750 9688 1750 0 wbs_dat_i[2]
rlabel metal2 10584 2058 10584 2058 0 wbs_dat_i[3]
rlabel metal2 9632 7448 9632 7448 0 wbs_dat_i[4]
rlabel metal2 11984 3304 11984 3304 0 wbs_dat_i[5]
rlabel metal2 2856 2968 2856 2968 0 wbs_dat_i[6]
rlabel metal2 13496 1918 13496 1918 0 wbs_dat_i[7]
rlabel metal2 14168 1470 14168 1470 0 wbs_dat_i[8]
rlabel metal2 14840 1470 14840 1470 0 wbs_dat_i[9]
rlabel metal2 8120 2058 8120 2058 0 wbs_dat_o[0]
rlabel metal2 15736 2478 15736 2478 0 wbs_dat_o[10]
rlabel metal2 16408 2198 16408 2198 0 wbs_dat_o[11]
rlabel metal2 17080 1246 17080 1246 0 wbs_dat_o[12]
rlabel metal2 17752 1246 17752 1246 0 wbs_dat_o[13]
rlabel metal2 18424 2086 18424 2086 0 wbs_dat_o[14]
rlabel metal2 19320 4088 19320 4088 0 wbs_dat_o[15]
rlabel metal2 9016 2058 9016 2058 0 wbs_dat_o[1]
rlabel metal3 7392 4088 7392 4088 0 wbs_dat_o[2]
rlabel metal2 11032 3752 11032 3752 0 wbs_dat_o[3]
rlabel metal2 11536 6552 11536 6552 0 wbs_dat_o[4]
rlabel metal2 12152 4872 12152 4872 0 wbs_dat_o[5]
rlabel metal2 13048 2058 13048 2058 0 wbs_dat_o[6]
rlabel metal2 13944 4088 13944 4088 0 wbs_dat_o[7]
rlabel metal3 11088 3416 11088 3416 0 wbs_dat_o[8]
rlabel metal2 15176 4592 15176 4592 0 wbs_dat_o[9]
rlabel metal2 2072 4592 2072 4592 0 wbs_sel_i[0]
rlabel metal2 2016 4200 2016 4200 0 wbs_sel_i[1]
rlabel metal2 4536 3472 4536 3472 0 wbs_stb_i
rlabel metal2 5768 5824 5768 5824 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
